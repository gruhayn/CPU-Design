
`include "ramVariables.h"

module ram
	#(
		parameter dataLength=`dataLength,
		parameter addressLegth=`addressLegth
	)
		(
			input [dataLength-1:0] SRAM_data_in ,
			output [dataLength-1:0] SRAM_data_out ,
			input SRAM_wr_n,
			input SRAM_cs_n ,
			input SRAM_oe_n ,
			input [addressLegth-1:0] SRAM_ADD_in ,
			
			output [addressLegth-1:0] SRAM_ADDR_out ,
			inout [dataLength-1:0] SRAM_DQ,
			output SRAM_WE_N,
			output SRAM_OE_N,
			output SRAM_UB_N,
			output SRAM_LB_N,
			output SRAM_CE_N
		);

reg [dataLength-1:0] sram_mem [2**addressLegth-1:0];

assign SRAM_LB_N=0;
assign SRAM_UB_N=0;
assign SRAM_CE_N = SRAM_cs_n;
assign SRAM_WE_N = SRAM_wr_n;
assign SRAM_OE_N = SRAM_oe_n;
assign SRAM_ADDR_out = SRAM_ADD_in;
//assign SRAM_data_out = ( (!SRAM_cs_n & !SRAM_oe_n & SRAM_wr_n) ) ? sram_mem[SRAM_ADD_in] : {16{1'bz}};
assign SRAM_data_out = sram_mem[SRAM_ADD_in];

always @(*) begin
	if (SRAM_cs_n==0 && SRAM_wr_n==0) begin
		sram_mem[SRAM_ADD_in] = SRAM_data_in ;
	end
end

initial begin

	sram_mem[0] = 16'b1001111111111100;
	sram_mem[1] = 16'b1010001111111100;
	sram_mem[2] = 16'b1011110110001101;
	sram_mem[3] = 16'b1010010000000000;
	sram_mem[4] = 16'b1010100000000000;
	sram_mem[5] = 16'b1011110111101000;
	sram_mem[6] = 16'b1001110000000000;
	sram_mem[7] = 16'b1010000000000000;
	sram_mem[8] = 16'b1011110110001001;
	sram_mem[9] = 16'b1010010000010000;
	sram_mem[10] = 16'b1010100000000000;
	sram_mem[11] = 16'b1010110111101010;
	sram_mem[12] = 16'b0001110101000000;
	sram_mem[13] = 16'b1010010011000000;
	sram_mem[14] = 16'b1010100000000000;
	sram_mem[15] = 16'b1001000100101010;
	sram_mem[16] = 16'b0101010111100000;
	sram_mem[17] = 16'b1011110110001011;
	sram_mem[18] = 16'b1011110101000100;
	sram_mem[19] = 16'b0000100100100100;
	sram_mem[20] = 16'b0010000010000000;
	sram_mem[21] = 16'b1010010010110000;
	sram_mem[22] = 16'b1010100000000000;
	sram_mem[23] = 16'b1001000101100100;
	sram_mem[24] = 16'b0101010111100000;
	sram_mem[25] = 16'b1011110100000100;
	sram_mem[26] = 16'b0000000101100100;
	sram_mem[27] = 16'b1011110010000101;
	sram_mem[28] = 16'b0001100010100000;
	sram_mem[29] = 16'b1010110010000110;
	sram_mem[30] = 16'b1010110010100111;
	sram_mem[31] = 16'b1010010010100000;
	sram_mem[32] = 16'b1010100000000000;
	sram_mem[33] = 16'b1001000011000111;
	sram_mem[34] = 16'b0110010111100000;
	sram_mem[35] = 16'b1011110011000000;
	sram_mem[36] = 16'b1011110011100110;
	sram_mem[37] = 16'b1011110000000111;
	sram_mem[38] = 16'b1011100011000100;
	sram_mem[39] = 16'b1011100011100101;
	sram_mem[40] = 16'b0001100101100000;
	sram_mem[41] = 16'b1010010001001000;
	sram_mem[42] = 16'b1010100000000000;
	sram_mem[43] = 16'b1000110111100000;
	sram_mem[44] = 16'b0001100100100000;
	sram_mem[45] = 16'b1010010000110100;
	sram_mem[46] = 16'b1010100000000000;
	sram_mem[47] = 16'b1000110111100000;
	sram_mem[48] = 16'b1011110110001001;
	sram_mem[49] = 16'b1010010011100000;
	sram_mem[50] = 16'b1010100000000000;
	sram_mem[51] = 16'b1001000100101010;
	sram_mem[52] = 16'b0100110111100000;
	sram_mem[53] = 16'b1010110100000100;
	sram_mem[54] = 16'b0001100100000000;
	sram_mem[55] = 16'b0001100100100000;
	sram_mem[56] = 16'b1101110000000000;
	sram_mem[65536] = 16'b0000000000000010;
	sram_mem[65537] = 16'b1111111111110111;
	sram_mem[65538] = 16'b0000000000000001;
	sram_mem[65539] = 16'b0000000000000011;
	sram_mem[65540] = 16'b0000000000000100;
	sram_mem[65541] = 16'b0000000000000000;
	sram_mem[65542] = 16'b0000000000000000;
	sram_mem[65543] = 16'b0000000000000000;
	sram_mem[65544] = 16'b0000000000000000;
	sram_mem[65545] = 16'b0000000000000000;
	sram_mem[65546] = 16'b0000000000000000;
	sram_mem[65547] = 16'b0000000000000000;
	sram_mem[65548] = 16'b0000000000000000;
	sram_mem[65549] = 16'b0000000000000000;
	sram_mem[65550] = 16'b0000000000000000;
	sram_mem[65551] = 16'b0000000000000000;
	sram_mem[65552] = 16'b0000000000000000;
	sram_mem[65553] = 16'b0000000000000000;
	sram_mem[65554] = 16'b0000000000000000;
	sram_mem[65555] = 16'b0000000000000000;
	sram_mem[65556] = 16'b0000000000000000;
	sram_mem[65557] = 16'b0000000000000000;
	sram_mem[65558] = 16'b0000000000000000;
	sram_mem[65559] = 16'b0000000000000000;
	sram_mem[65560] = 16'b0000000000000000;
	sram_mem[65561] = 16'b0000000000000000;
	sram_mem[65562] = 16'b0000000000000000;
	sram_mem[65563] = 16'b0000000000000000;
	sram_mem[65564] = 16'b0000000000000000;
	sram_mem[65565] = 16'b0000000000000000;
	sram_mem[65566] = 16'b0000000000000000;
	sram_mem[65567] = 16'b0000000000000000;
	sram_mem[65568] = 16'b0000000000000000;
	sram_mem[65569] = 16'b0000000000000000;
	sram_mem[65570] = 16'b0000000000000000;
	sram_mem[65571] = 16'b0000000000000000;
	sram_mem[65572] = 16'b0000000000000000;
	sram_mem[65573] = 16'b0000000000000000;
	sram_mem[65574] = 16'b0000000000000000;
	sram_mem[65575] = 16'b0000000000000000;
	sram_mem[65576] = 16'b0000000000000000;
	sram_mem[65577] = 16'b0000000000000000;
	sram_mem[65578] = 16'b0000000000000000;
	sram_mem[65579] = 16'b0000000000000000;
	sram_mem[65580] = 16'b0000000000000000;
	sram_mem[65581] = 16'b0000000000000000;
	sram_mem[65582] = 16'b0000000000000000;
	sram_mem[65583] = 16'b0000000000000000;
	sram_mem[65584] = 16'b0000000000000000;
	sram_mem[65585] = 16'b0000000000000000;
	sram_mem[65586] = 16'b0000000000000000;
	sram_mem[65587] = 16'b0000000000000000;
	sram_mem[65588] = 16'b0000000000000000;
	sram_mem[65589] = 16'b0000000000000000;
	sram_mem[65590] = 16'b0000000000000000;
	sram_mem[65591] = 16'b0000000000000000;
	sram_mem[65592] = 16'b0000000000000000;
	sram_mem[65593] = 16'b0000000000000000;
	sram_mem[65594] = 16'b0000000000000000;
	sram_mem[65595] = 16'b0000000000000000;
	sram_mem[65596] = 16'b0000000000000000;
	sram_mem[65597] = 16'b0000000000000000;
	sram_mem[65598] = 16'b0000000000000000;
	sram_mem[65599] = 16'b0000000000000000;
	sram_mem[65600] = 16'b0000000000000000;
	sram_mem[65601] = 16'b0000000000000000;
	sram_mem[65602] = 16'b0000000000000000;
	sram_mem[65603] = 16'b0000000000000000;
	sram_mem[65604] = 16'b0000000000000000;
	sram_mem[65605] = 16'b0000000000000000;
	sram_mem[65606] = 16'b0000000000000000;
	sram_mem[65607] = 16'b0000000000000000;
	sram_mem[65608] = 16'b0000000000000000;
	sram_mem[65609] = 16'b0000000000000000;
	sram_mem[65610] = 16'b0000000000000000;
	sram_mem[65611] = 16'b0000000000000000;
	sram_mem[65612] = 16'b0000000000000000;
	sram_mem[65613] = 16'b0000000000000000;
	sram_mem[65614] = 16'b0000000000000000;
	sram_mem[65615] = 16'b0000000000000000;
	sram_mem[65616] = 16'b0000000000000000;
	sram_mem[65617] = 16'b0000000000000000;
	sram_mem[65618] = 16'b0000000000000000;
	sram_mem[65619] = 16'b0000000000000000;
	sram_mem[65620] = 16'b0000000000000000;
	sram_mem[65621] = 16'b0000000000000000;
	sram_mem[65622] = 16'b0000000000000000;
	sram_mem[65623] = 16'b0000000000000000;
	sram_mem[65624] = 16'b0000000000000000;
	sram_mem[65625] = 16'b0000000000000000;
	sram_mem[65626] = 16'b0000000000000000;
	sram_mem[65627] = 16'b0000000000000000;
	sram_mem[65628] = 16'b0000000000000000;
	sram_mem[65629] = 16'b0000000000000000;
	sram_mem[65630] = 16'b0000000000000000;
	sram_mem[65631] = 16'b0000000000000000;
	sram_mem[65632] = 16'b0000000000000000;
	sram_mem[65633] = 16'b0000000000000000;
	sram_mem[65634] = 16'b0000000000000000;
	sram_mem[65635] = 16'b0000000000000000;
	sram_mem[65636] = 16'b0000000000000000;
	sram_mem[65637] = 16'b0000000000000000;
	sram_mem[65638] = 16'b0000000000000000;
	sram_mem[65639] = 16'b0000000000000000;
	sram_mem[65640] = 16'b0000000000000000;
	sram_mem[65641] = 16'b0000000000000000;
	sram_mem[65642] = 16'b0000000000000000;
	sram_mem[65643] = 16'b0000000000000000;
	sram_mem[65644] = 16'b0000000000000000;
	sram_mem[65645] = 16'b0000000000000000;
	sram_mem[65646] = 16'b0000000000000000;
	sram_mem[65647] = 16'b0000000000000000;
	sram_mem[65648] = 16'b0000000000000000;
	sram_mem[65649] = 16'b0000000000000000;
	sram_mem[65650] = 16'b0000000000000000;
	sram_mem[65651] = 16'b0000000000000000;
	sram_mem[65652] = 16'b0000000000000000;
	sram_mem[65653] = 16'b0000000000000000;
	sram_mem[65654] = 16'b0000000000000000;
	sram_mem[65655] = 16'b0000000000000000;
	sram_mem[65656] = 16'b0000000000000000;
	sram_mem[65657] = 16'b0000000000000000;
	sram_mem[65658] = 16'b0000000000000000;
	sram_mem[65659] = 16'b0000000000000000;
	sram_mem[65660] = 16'b0000000000000000;
	sram_mem[65661] = 16'b0000000000000000;
	sram_mem[65662] = 16'b0000000000000000;
	sram_mem[65663] = 16'b0000000000000000;
	sram_mem[65664] = 16'b0000000000000000;
	sram_mem[65665] = 16'b0000000000000000;
	sram_mem[65666] = 16'b0000000000000000;
	sram_mem[65667] = 16'b0000000000000000;
	sram_mem[65668] = 16'b0000000000000000;
	sram_mem[65669] = 16'b0000000000000000;
	sram_mem[65670] = 16'b0000000000000000;
	sram_mem[65671] = 16'b0000000000000000;
	sram_mem[65672] = 16'b0000000000000000;
	sram_mem[65673] = 16'b0000000000000000;
	sram_mem[65674] = 16'b0000000000000000;
	sram_mem[65675] = 16'b0000000000000000;
	sram_mem[65676] = 16'b0000000000000000;
	sram_mem[65677] = 16'b0000000000000000;
	sram_mem[65678] = 16'b0000000000000000;
	sram_mem[65679] = 16'b0000000000000000;
	sram_mem[65680] = 16'b0000000000000000;
	sram_mem[65681] = 16'b0000000000000000;
	sram_mem[65682] = 16'b0000000000000000;
	sram_mem[65683] = 16'b0000000000000000;
	sram_mem[65684] = 16'b0000000000000000;
	sram_mem[65685] = 16'b0000000000000000;
	sram_mem[65686] = 16'b0000000000000000;
	sram_mem[65687] = 16'b0000000000000000;
	sram_mem[65688] = 16'b0000000000000000;
	sram_mem[65689] = 16'b0000000000000000;
	sram_mem[65690] = 16'b0000000000000000;
	sram_mem[65691] = 16'b0000000000000000;
	sram_mem[65692] = 16'b0000000000000000;
	sram_mem[65693] = 16'b0000000000000000;
	sram_mem[65694] = 16'b0000000000000000;
	sram_mem[65695] = 16'b0000000000000000;
	sram_mem[65696] = 16'b0000000000000000;
	sram_mem[65697] = 16'b0000000000000000;
	sram_mem[65698] = 16'b0000000000000000;
	sram_mem[65699] = 16'b0000000000000000;
	sram_mem[65700] = 16'b0000000000000000;
	sram_mem[65701] = 16'b0000000000000000;
	sram_mem[65702] = 16'b0000000000000000;
	sram_mem[65703] = 16'b0000000000000000;
	sram_mem[65704] = 16'b0000000000000000;
	sram_mem[65705] = 16'b0000000000000000;
	sram_mem[65706] = 16'b0000000000000000;
	sram_mem[65707] = 16'b0000000000000000;
	sram_mem[65708] = 16'b0000000000000000;
	sram_mem[65709] = 16'b0000000000000000;
	sram_mem[65710] = 16'b0000000000000000;
	sram_mem[65711] = 16'b0000000000000000;
	sram_mem[65712] = 16'b0000000000000000;
	sram_mem[65713] = 16'b0000000000000000;
	sram_mem[65714] = 16'b0000000000000000;
	sram_mem[65715] = 16'b0000000000000000;
	sram_mem[65716] = 16'b0000000000000000;
	sram_mem[65717] = 16'b0000000000000000;
	sram_mem[65718] = 16'b0000000000000000;
	sram_mem[65719] = 16'b0000000000000000;
	sram_mem[65720] = 16'b0000000000000000;
	sram_mem[65721] = 16'b0000000000000000;
	sram_mem[65722] = 16'b0000000000000000;
	sram_mem[65723] = 16'b0000000000000000;
	sram_mem[65724] = 16'b0000000000000000;
	sram_mem[65725] = 16'b0000000000000000;
	sram_mem[65726] = 16'b0000000000000000;
	sram_mem[65727] = 16'b0000000000000000;
	sram_mem[65728] = 16'b0000000000000000;
	sram_mem[65729] = 16'b0000000000000000;
	sram_mem[65730] = 16'b0000000000000000;
	sram_mem[65731] = 16'b0000000000000000;
	sram_mem[65732] = 16'b0000000000000000;
	sram_mem[65733] = 16'b0000000000000000;
	sram_mem[65734] = 16'b0000000000000000;
	sram_mem[65735] = 16'b0000000000000000;
	sram_mem[65736] = 16'b0000000000000000;
	sram_mem[65737] = 16'b0000000000000000;
	sram_mem[65738] = 16'b0000000000000000;
	sram_mem[65739] = 16'b0000000000000000;
	sram_mem[65740] = 16'b0000000000000000;
	sram_mem[65741] = 16'b0000000000000000;
	sram_mem[65742] = 16'b0000000000000000;
	sram_mem[65743] = 16'b0000000000000000;
	sram_mem[65744] = 16'b0000000000000000;
	sram_mem[65745] = 16'b0000000000000000;
	sram_mem[65746] = 16'b0000000000000000;
	sram_mem[65747] = 16'b0000000000000000;
	sram_mem[65748] = 16'b0000000000000000;
	sram_mem[65749] = 16'b0000000000000000;
	sram_mem[65750] = 16'b0000000000000000;
	sram_mem[65751] = 16'b0000000000000000;
	sram_mem[65752] = 16'b0000000000000000;
	sram_mem[65753] = 16'b0000000000000000;
	sram_mem[65754] = 16'b0000000000000000;
	sram_mem[65755] = 16'b0000000000000000;
	sram_mem[65756] = 16'b0000000000000000;
	sram_mem[65757] = 16'b0000000000000000;
	sram_mem[65758] = 16'b0000000000000000;
	sram_mem[65759] = 16'b0000000000000000;
	sram_mem[65760] = 16'b0000000000000000;
	sram_mem[65761] = 16'b0000000000000000;
	sram_mem[65762] = 16'b0000000000000000;
	sram_mem[65763] = 16'b0000000000000000;
	sram_mem[65764] = 16'b0000000000000000;
	sram_mem[65765] = 16'b0000000000000000;
	sram_mem[65766] = 16'b0000000000000000;
	sram_mem[65767] = 16'b0000000000000000;
	sram_mem[65768] = 16'b0000000000000000;
	sram_mem[65769] = 16'b0000000000000000;
	sram_mem[65770] = 16'b0000000000000000;
	sram_mem[65771] = 16'b0000000000000000;
	sram_mem[65772] = 16'b0000000000000000;
	sram_mem[65773] = 16'b0000000000000000;
	sram_mem[65774] = 16'b0000000000000000;
	sram_mem[65775] = 16'b0000000000000000;
	sram_mem[65776] = 16'b0000000000000000;
	sram_mem[65777] = 16'b0000000000000000;
	sram_mem[65778] = 16'b0000000000000000;
	sram_mem[65779] = 16'b0000000000000000;
	sram_mem[65780] = 16'b0000000000000000;
	sram_mem[65781] = 16'b0000000000000000;
	sram_mem[65782] = 16'b0000000000000000;
	sram_mem[65783] = 16'b0000000000000000;
	sram_mem[65784] = 16'b0000000000000000;
	sram_mem[65785] = 16'b0000000000000000;
	sram_mem[65786] = 16'b0000000000000000;
	sram_mem[65787] = 16'b0000000000000000;
	sram_mem[65788] = 16'b0000000000000000;
	sram_mem[65789] = 16'b0000000000000000;
	sram_mem[65790] = 16'b0000000000000000;
	sram_mem[65791] = 16'b0000000000000000;
	sram_mem[65792] = 16'b0000000000000000;
	sram_mem[65793] = 16'b0000000000000000;
	sram_mem[65794] = 16'b0000000000000000;
	sram_mem[65795] = 16'b0000000000000000;
	sram_mem[65796] = 16'b0000000000000000;
	sram_mem[65797] = 16'b0000000000000000;
	sram_mem[65798] = 16'b0000000000000000;
	sram_mem[65799] = 16'b0000000000000000;
	sram_mem[65800] = 16'b0000000000000000;
	sram_mem[65801] = 16'b0000000000000000;
	sram_mem[65802] = 16'b0000000000000000;
	sram_mem[65803] = 16'b0000000000000000;
	sram_mem[65804] = 16'b0000000000000000;
	sram_mem[65805] = 16'b0000000000000000;
	sram_mem[65806] = 16'b0000000000000000;
	sram_mem[65807] = 16'b0000000000000000;
	sram_mem[65808] = 16'b0000000000000000;
	sram_mem[65809] = 16'b0000000000000000;
	sram_mem[65810] = 16'b0000000000000000;
	sram_mem[65811] = 16'b0000000000000000;
	sram_mem[65812] = 16'b0000000000000000;
	sram_mem[65813] = 16'b0000000000000000;
	sram_mem[65814] = 16'b0000000000000000;
	sram_mem[65815] = 16'b0000000000000000;
	sram_mem[65816] = 16'b0000000000000000;
	sram_mem[65817] = 16'b0000000000000000;
	sram_mem[65818] = 16'b0000000000000000;
	sram_mem[65819] = 16'b0000000000000000;
	sram_mem[65820] = 16'b0000000000000000;
	sram_mem[65821] = 16'b0000000000000000;
	sram_mem[65822] = 16'b0000000000000000;
	sram_mem[65823] = 16'b0000000000000000;
	sram_mem[65824] = 16'b0000000000000000;
	sram_mem[65825] = 16'b0000000000000000;
	sram_mem[65826] = 16'b0000000000000000;
	sram_mem[65827] = 16'b0000000000000000;
	sram_mem[65828] = 16'b0000000000000000;
	sram_mem[65829] = 16'b0000000000000000;
	sram_mem[65830] = 16'b0000000000000000;
	sram_mem[65831] = 16'b0000000000000000;
	sram_mem[65832] = 16'b0000000000000000;
	sram_mem[65833] = 16'b0000000000000000;
	sram_mem[65834] = 16'b0000000000000000;
	sram_mem[65835] = 16'b0000000000000000;
	sram_mem[65836] = 16'b0000000000000000;
	sram_mem[65837] = 16'b0000000000000000;
	sram_mem[65838] = 16'b0000000000000000;
	sram_mem[65839] = 16'b0000000000000000;
	sram_mem[65840] = 16'b0000000000000000;
	sram_mem[65841] = 16'b0000000000000000;
	sram_mem[65842] = 16'b0000000000000000;
	sram_mem[65843] = 16'b0000000000000000;
	sram_mem[65844] = 16'b0000000000000000;
	sram_mem[65845] = 16'b0000000000000000;
	sram_mem[65846] = 16'b0000000000000000;
	sram_mem[65847] = 16'b0000000000000000;
	sram_mem[65848] = 16'b0000000000000000;
	sram_mem[65849] = 16'b0000000000000000;
	sram_mem[65850] = 16'b0000000000000000;
	sram_mem[65851] = 16'b0000000000000000;
	sram_mem[65852] = 16'b0000000000000000;
	sram_mem[65853] = 16'b0000000000000000;
	sram_mem[65854] = 16'b0000000000000000;
	sram_mem[65855] = 16'b0000000000000000;
	sram_mem[65856] = 16'b0000000000000000;
	sram_mem[65857] = 16'b0000000000000000;
	sram_mem[65858] = 16'b0000000000000000;
	sram_mem[65859] = 16'b0000000000000000;
	sram_mem[65860] = 16'b0000000000000000;
	sram_mem[65861] = 16'b0000000000000000;
	sram_mem[65862] = 16'b0000000000000000;
	sram_mem[65863] = 16'b0000000000000000;
	sram_mem[65864] = 16'b0000000000000000;
	sram_mem[65865] = 16'b0000000000000000;
	sram_mem[65866] = 16'b0000000000000000;
	sram_mem[65867] = 16'b0000000000000000;
	sram_mem[65868] = 16'b0000000000000000;
	sram_mem[65869] = 16'b0000000000000000;
	sram_mem[65870] = 16'b0000000000000000;
	sram_mem[65871] = 16'b0000000000000000;
	sram_mem[65872] = 16'b0000000000000000;
	sram_mem[65873] = 16'b0000000000000000;
	sram_mem[65874] = 16'b0000000000000000;
	sram_mem[65875] = 16'b0000000000000000;
	sram_mem[65876] = 16'b0000000000000000;
	sram_mem[65877] = 16'b0000000000000000;
	sram_mem[65878] = 16'b0000000000000000;
	sram_mem[65879] = 16'b0000000000000000;
	sram_mem[65880] = 16'b0000000000000000;
	sram_mem[65881] = 16'b0000000000000000;
	sram_mem[65882] = 16'b0000000000000000;
	sram_mem[65883] = 16'b0000000000000000;
	sram_mem[65884] = 16'b0000000000000000;
	sram_mem[65885] = 16'b0000000000000000;
	sram_mem[65886] = 16'b0000000000000000;
	sram_mem[65887] = 16'b0000000000000000;
	sram_mem[65888] = 16'b0000000000000000;
	sram_mem[65889] = 16'b0000000000000000;
	sram_mem[65890] = 16'b0000000000000000;
	sram_mem[65891] = 16'b0000000000000000;
	sram_mem[65892] = 16'b0000000000000000;
	sram_mem[65893] = 16'b0000000000000000;
	sram_mem[65894] = 16'b0000000000000000;
	sram_mem[65895] = 16'b0000000000000000;
	sram_mem[65896] = 16'b0000000000000000;
	sram_mem[65897] = 16'b0000000000000000;
	sram_mem[65898] = 16'b0000000000000000;
	sram_mem[65899] = 16'b0000000000000000;
	sram_mem[65900] = 16'b0000000000000000;
	sram_mem[65901] = 16'b0000000000000000;
	sram_mem[65902] = 16'b0000000000000000;
	sram_mem[65903] = 16'b0000000000000000;
	sram_mem[65904] = 16'b0000000000000000;
	sram_mem[65905] = 16'b0000000000000000;
	sram_mem[65906] = 16'b0000000000000000;
	sram_mem[65907] = 16'b0000000000000000;
	sram_mem[65908] = 16'b0000000000000000;
	sram_mem[65909] = 16'b0000000000000000;
	sram_mem[65910] = 16'b0000000000000000;
	sram_mem[65911] = 16'b0000000000000000;
	sram_mem[65912] = 16'b0000000000000000;
	sram_mem[65913] = 16'b0000000000000000;
	sram_mem[65914] = 16'b0000000000000000;
	sram_mem[65915] = 16'b0000000000000000;
	sram_mem[65916] = 16'b0000000000000000;
	sram_mem[65917] = 16'b0000000000000000;
	sram_mem[65918] = 16'b0000000000000000;
	sram_mem[65919] = 16'b0000000000000000;
	sram_mem[65920] = 16'b0000000000000000;
	sram_mem[65921] = 16'b0000000000000000;
	sram_mem[65922] = 16'b0000000000000000;
	sram_mem[65923] = 16'b0000000000000000;
	sram_mem[65924] = 16'b0000000000000000;
	sram_mem[65925] = 16'b0000000000000000;
	sram_mem[65926] = 16'b0000000000000000;
	sram_mem[65927] = 16'b0000000000000000;
	sram_mem[65928] = 16'b0000000000000000;
	sram_mem[65929] = 16'b0000000000000000;
	sram_mem[65930] = 16'b0000000000000000;
	sram_mem[65931] = 16'b0000000000000000;
	sram_mem[65932] = 16'b0000000000000000;
	sram_mem[65933] = 16'b0000000000000000;
	sram_mem[65934] = 16'b0000000000000000;
	sram_mem[65935] = 16'b0000000000000000;
	sram_mem[65936] = 16'b0000000000000000;
	sram_mem[65937] = 16'b0000000000000000;
	sram_mem[65938] = 16'b0000000000000000;
	sram_mem[65939] = 16'b0000000000000000;
	sram_mem[65940] = 16'b0000000000000000;
	sram_mem[65941] = 16'b0000000000000000;
	sram_mem[65942] = 16'b0000000000000000;
	sram_mem[65943] = 16'b0000000000000000;
	sram_mem[65944] = 16'b0000000000000000;
	sram_mem[65945] = 16'b0000000000000000;
	sram_mem[65946] = 16'b0000000000000000;
	sram_mem[65947] = 16'b0000000000000000;
	sram_mem[65948] = 16'b0000000000000000;
	sram_mem[65949] = 16'b0000000000000000;
	sram_mem[65950] = 16'b0000000000000000;
	sram_mem[65951] = 16'b0000000000000000;
	sram_mem[65952] = 16'b0000000000000000;
	sram_mem[65953] = 16'b0000000000000000;
	sram_mem[65954] = 16'b0000000000000000;
	sram_mem[65955] = 16'b0000000000000000;
	sram_mem[65956] = 16'b0000000000000000;
	sram_mem[65957] = 16'b0000000000000000;
	sram_mem[65958] = 16'b0000000000000000;
	sram_mem[65959] = 16'b0000000000000000;
	sram_mem[65960] = 16'b0000000000000000;
	sram_mem[65961] = 16'b0000000000000000;
	sram_mem[65962] = 16'b0000000000000000;
	sram_mem[65963] = 16'b0000000000000000;
	sram_mem[65964] = 16'b0000000000000000;
	sram_mem[65965] = 16'b0000000000000000;
	sram_mem[65966] = 16'b0000000000000000;
	sram_mem[65967] = 16'b0000000000000000;
	sram_mem[65968] = 16'b0000000000000000;
	sram_mem[65969] = 16'b0000000000000000;
	sram_mem[65970] = 16'b0000000000000000;
	sram_mem[65971] = 16'b0000000000000000;
	sram_mem[65972] = 16'b0000000000000000;
	sram_mem[65973] = 16'b0000000000000000;
	sram_mem[65974] = 16'b0000000000000000;
	sram_mem[65975] = 16'b0000000000000000;
	sram_mem[65976] = 16'b0000000000000000;
	sram_mem[65977] = 16'b0000000000000000;
	sram_mem[65978] = 16'b0000000000000000;
	sram_mem[65979] = 16'b0000000000000000;
	sram_mem[65980] = 16'b0000000000000000;
	sram_mem[65981] = 16'b0000000000000000;
	sram_mem[65982] = 16'b0000000000000000;
	sram_mem[65983] = 16'b0000000000000000;
	sram_mem[65984] = 16'b0000000000000000;
	sram_mem[65985] = 16'b0000000000000000;
	sram_mem[65986] = 16'b0000000000000000;
	sram_mem[65987] = 16'b0000000000000000;
	sram_mem[65988] = 16'b0000000000000000;
	sram_mem[65989] = 16'b0000000000000000;
	sram_mem[65990] = 16'b0000000000000000;
	sram_mem[65991] = 16'b0000000000000000;
	sram_mem[65992] = 16'b0000000000000000;
	sram_mem[65993] = 16'b0000000000000000;
	sram_mem[65994] = 16'b0000000000000000;
	sram_mem[65995] = 16'b0000000000000000;
	sram_mem[65996] = 16'b0000000000000000;
	sram_mem[65997] = 16'b0000000000000000;
	sram_mem[65998] = 16'b0000000000000000;
	sram_mem[65999] = 16'b0000000000000000;
	sram_mem[66000] = 16'b0000000000000000;
	sram_mem[66001] = 16'b0000000000000000;
	sram_mem[66002] = 16'b0000000000000000;
	sram_mem[66003] = 16'b0000000000000000;
	sram_mem[66004] = 16'b0000000000000000;
	sram_mem[66005] = 16'b0000000000000000;
	sram_mem[66006] = 16'b0000000000000000;
	sram_mem[66007] = 16'b0000000000000000;
	sram_mem[66008] = 16'b0000000000000000;
	sram_mem[66009] = 16'b0000000000000000;
	sram_mem[66010] = 16'b0000000000000000;
	sram_mem[66011] = 16'b0000000000000000;
	sram_mem[66012] = 16'b0000000000000000;
	sram_mem[66013] = 16'b0000000000000000;
	sram_mem[66014] = 16'b0000000000000000;
	sram_mem[66015] = 16'b0000000000000000;
	sram_mem[66016] = 16'b0000000000000000;
	sram_mem[66017] = 16'b0000000000000000;
	sram_mem[66018] = 16'b0000000000000000;
	sram_mem[66019] = 16'b0000000000000000;
	sram_mem[66020] = 16'b0000000000000000;
	sram_mem[66021] = 16'b0000000000000000;
	sram_mem[66022] = 16'b0000000000000000;
	sram_mem[66023] = 16'b0000000000000000;
	sram_mem[66024] = 16'b0000000000000000;
	sram_mem[66025] = 16'b0000000000000000;
	sram_mem[66026] = 16'b0000000000000000;
	sram_mem[66027] = 16'b0000000000000000;
	sram_mem[66028] = 16'b0000000000000000;
	sram_mem[66029] = 16'b0000000000000000;
	sram_mem[66030] = 16'b0000000000000000;
	sram_mem[66031] = 16'b0000000000000000;
	sram_mem[66032] = 16'b0000000000000000;
	sram_mem[66033] = 16'b0000000000000000;
	sram_mem[66034] = 16'b0000000000000000;
	sram_mem[66035] = 16'b0000000000000000;
	sram_mem[66036] = 16'b0000000000000000;
	sram_mem[66037] = 16'b0000000000000000;
	sram_mem[66038] = 16'b0000000000000000;
	sram_mem[66039] = 16'b0000000000000000;
	sram_mem[66040] = 16'b0000000000000000;
	sram_mem[66041] = 16'b0000000000000000;
	sram_mem[66042] = 16'b0000000000000000;
	sram_mem[66043] = 16'b0000000000000000;
	sram_mem[66044] = 16'b0000000000000000;
	sram_mem[66045] = 16'b0000000000000000;
	sram_mem[66046] = 16'b0000000000000000;
	sram_mem[66047] = 16'b0000000000000000;
	sram_mem[66048] = 16'b0000000000000000;
	sram_mem[66049] = 16'b0000000000000000;
	sram_mem[66050] = 16'b0000000000000000;
	sram_mem[66051] = 16'b0000000000000000;
	sram_mem[66052] = 16'b0000000000000000;
	sram_mem[66053] = 16'b0000000000000000;
	sram_mem[66054] = 16'b0000000000000000;
	sram_mem[66055] = 16'b0000000000000000;
	sram_mem[66056] = 16'b0000000000000000;
	sram_mem[66057] = 16'b0000000000000000;
	sram_mem[66058] = 16'b0000000000000000;
	sram_mem[66059] = 16'b0000000000000000;
	sram_mem[66060] = 16'b0000000000000000;
	sram_mem[66061] = 16'b0000000000000000;
	sram_mem[66062] = 16'b0000000000000000;
	sram_mem[66063] = 16'b0000000000000000;
	sram_mem[66064] = 16'b0000000000000000;
	sram_mem[66065] = 16'b0000000000000000;
	sram_mem[66066] = 16'b0000000000000000;
	sram_mem[66067] = 16'b0000000000000000;
	sram_mem[66068] = 16'b0000000000000000;
	sram_mem[66069] = 16'b0000000000000000;
	sram_mem[66070] = 16'b0000000000000000;
	sram_mem[66071] = 16'b0000000000000000;
	sram_mem[66072] = 16'b0000000000000000;
	sram_mem[66073] = 16'b0000000000000000;
	sram_mem[66074] = 16'b0000000000000000;
	sram_mem[66075] = 16'b0000000000000000;
	sram_mem[66076] = 16'b0000000000000000;
	sram_mem[66077] = 16'b0000000000000000;
	sram_mem[66078] = 16'b0000000000000000;
	sram_mem[66079] = 16'b0000000000000000;
	sram_mem[66080] = 16'b0000000000000000;
	sram_mem[66081] = 16'b0000000000000000;
	sram_mem[66082] = 16'b0000000000000000;
	sram_mem[66083] = 16'b0000000000000000;
	sram_mem[66084] = 16'b0000000000000000;
	sram_mem[66085] = 16'b0000000000000000;
	sram_mem[66086] = 16'b0000000000000000;
	sram_mem[66087] = 16'b0000000000000000;
	sram_mem[66088] = 16'b0000000000000000;
	sram_mem[66089] = 16'b0000000000000000;
	sram_mem[66090] = 16'b0000000000000000;
	sram_mem[66091] = 16'b0000000000000000;
	sram_mem[66092] = 16'b0000000000000000;
	sram_mem[66093] = 16'b0000000000000000;
	sram_mem[66094] = 16'b0000000000000000;
	sram_mem[66095] = 16'b0000000000000000;
	sram_mem[66096] = 16'b0000000000000000;
	sram_mem[66097] = 16'b0000000000000000;
	sram_mem[66098] = 16'b0000000000000000;
	sram_mem[66099] = 16'b0000000000000000;
	sram_mem[66100] = 16'b0000000000000000;
	sram_mem[66101] = 16'b0000000000000000;
	sram_mem[66102] = 16'b0000000000000000;
	sram_mem[66103] = 16'b0000000000000000;
	sram_mem[66104] = 16'b0000000000000000;
	sram_mem[66105] = 16'b0000000000000000;
	sram_mem[66106] = 16'b0000000000000000;
	sram_mem[66107] = 16'b0000000000000000;
	sram_mem[66108] = 16'b0000000000000000;
	sram_mem[66109] = 16'b0000000000000000;
	sram_mem[66110] = 16'b0000000000000000;
	sram_mem[66111] = 16'b0000000000000000;
	sram_mem[66112] = 16'b0000000000000000;
	sram_mem[66113] = 16'b0000000000000000;
	sram_mem[66114] = 16'b0000000000000000;
	sram_mem[66115] = 16'b0000000000000000;
	sram_mem[66116] = 16'b0000000000000000;
	sram_mem[66117] = 16'b0000000000000000;
	sram_mem[66118] = 16'b0000000000000000;
	sram_mem[66119] = 16'b0000000000000000;
	sram_mem[66120] = 16'b0000000000000000;
	sram_mem[66121] = 16'b0000000000000000;
	sram_mem[66122] = 16'b0000000000000000;
	sram_mem[66123] = 16'b0000000000000000;
	sram_mem[66124] = 16'b0000000000000000;
	sram_mem[66125] = 16'b0000000000000000;
	sram_mem[66126] = 16'b0000000000000000;
	sram_mem[66127] = 16'b0000000000000000;
	sram_mem[66128] = 16'b0000000000000000;
	sram_mem[66129] = 16'b0000000000000000;
	sram_mem[66130] = 16'b0000000000000000;
	sram_mem[66131] = 16'b0000000000000000;
	sram_mem[66132] = 16'b0000000000000000;
	sram_mem[66133] = 16'b0000000000000000;
	sram_mem[66134] = 16'b0000000000000000;
	sram_mem[66135] = 16'b0000000000000000;
	sram_mem[66136] = 16'b0000000000000000;
	sram_mem[66137] = 16'b0000000000000000;
	sram_mem[66138] = 16'b0000000000000000;
	sram_mem[66139] = 16'b0000000000000000;
	sram_mem[66140] = 16'b0000000000000000;
	sram_mem[66141] = 16'b0000000000000000;
	sram_mem[66142] = 16'b0000000000000000;
	sram_mem[66143] = 16'b0000000000000000;
	sram_mem[66144] = 16'b0000000000000000;
	sram_mem[66145] = 16'b0000000000000000;
	sram_mem[66146] = 16'b0000000000000000;
	sram_mem[66147] = 16'b0000000000000000;
	sram_mem[66148] = 16'b0000000000000000;
	sram_mem[66149] = 16'b0000000000000000;
	sram_mem[66150] = 16'b0000000000000000;
	sram_mem[66151] = 16'b0000000000000000;
	sram_mem[66152] = 16'b0000000000000000;
	sram_mem[66153] = 16'b0000000000000000;
	sram_mem[66154] = 16'b0000000000000000;
	sram_mem[66155] = 16'b0000000000000000;
	sram_mem[66156] = 16'b0000000000000000;
	sram_mem[66157] = 16'b0000000000000000;
	sram_mem[66158] = 16'b0000000000000000;
	sram_mem[66159] = 16'b0000000000000000;
	sram_mem[66160] = 16'b0000000000000000;
	sram_mem[66161] = 16'b0000000000000000;
	sram_mem[66162] = 16'b0000000000000000;
	sram_mem[66163] = 16'b0000000000000000;
	sram_mem[66164] = 16'b0000000000000000;
	sram_mem[66165] = 16'b0000000000000000;
	sram_mem[66166] = 16'b0000000000000000;
	sram_mem[66167] = 16'b0000000000000000;
	sram_mem[66168] = 16'b0000000000000000;
	sram_mem[66169] = 16'b0000000000000000;
	sram_mem[66170] = 16'b0000000000000000;
	sram_mem[66171] = 16'b0000000000000000;
	sram_mem[66172] = 16'b0000000000000000;
	sram_mem[66173] = 16'b0000000000000000;
	sram_mem[66174] = 16'b0000000000000000;
	sram_mem[66175] = 16'b0000000000000000;
	sram_mem[66176] = 16'b0000000000000000;
	sram_mem[66177] = 16'b0000000000000000;
	sram_mem[66178] = 16'b0000000000000000;
	sram_mem[66179] = 16'b0000000000000000;
	sram_mem[66180] = 16'b0000000000000000;
	sram_mem[66181] = 16'b0000000000000000;
	sram_mem[66182] = 16'b0000000000000000;
	sram_mem[66183] = 16'b0000000000000000;
	sram_mem[66184] = 16'b0000000000000000;
	sram_mem[66185] = 16'b0000000000000000;
	sram_mem[66186] = 16'b0000000000000000;
	sram_mem[66187] = 16'b0000000000000000;
	sram_mem[66188] = 16'b0000000000000000;
	sram_mem[66189] = 16'b0000000000000000;
	sram_mem[66190] = 16'b0000000000000000;
	sram_mem[66191] = 16'b0000000000000000;
	sram_mem[66192] = 16'b0000000000000000;
	sram_mem[66193] = 16'b0000000000000000;
	sram_mem[66194] = 16'b0000000000000000;
	sram_mem[66195] = 16'b0000000000000000;
	sram_mem[66196] = 16'b0000000000000000;
	sram_mem[66197] = 16'b0000000000000000;
	sram_mem[66198] = 16'b0000000000000000;
	sram_mem[66199] = 16'b0000000000000000;
	sram_mem[66200] = 16'b0000000000000000;
	sram_mem[66201] = 16'b0000000000000000;
	sram_mem[66202] = 16'b0000000000000000;
	sram_mem[66203] = 16'b0000000000000000;
	sram_mem[66204] = 16'b0000000000000000;
	sram_mem[66205] = 16'b0000000000000000;
	sram_mem[66206] = 16'b0000000000000000;
	sram_mem[66207] = 16'b0000000000000000;
	sram_mem[66208] = 16'b0000000000000000;
	sram_mem[66209] = 16'b0000000000000000;
	sram_mem[66210] = 16'b0000000000000000;
	sram_mem[66211] = 16'b0000000000000000;
	sram_mem[66212] = 16'b0000000000000000;
	sram_mem[66213] = 16'b0000000000000000;
	sram_mem[66214] = 16'b0000000000000000;
	sram_mem[66215] = 16'b0000000000000000;
	sram_mem[66216] = 16'b0000000000000000;
	sram_mem[66217] = 16'b0000000000000000;
	sram_mem[66218] = 16'b0000000000000000;
	sram_mem[66219] = 16'b0000000000000000;
	sram_mem[66220] = 16'b0000000000000000;
	sram_mem[66221] = 16'b0000000000000000;
	sram_mem[66222] = 16'b0000000000000000;
	sram_mem[66223] = 16'b0000000000000000;
	sram_mem[66224] = 16'b0000000000000000;
	sram_mem[66225] = 16'b0000000000000000;
	sram_mem[66226] = 16'b0000000000000000;
	sram_mem[66227] = 16'b0000000000000000;
	sram_mem[66228] = 16'b0000000000000000;
	sram_mem[66229] = 16'b0000000000000000;
	sram_mem[66230] = 16'b0000000000000000;
	sram_mem[66231] = 16'b0000000000000000;
	sram_mem[66232] = 16'b0000000000000000;
	sram_mem[66233] = 16'b0000000000000000;
	sram_mem[66234] = 16'b0000000000000000;
	sram_mem[66235] = 16'b0000000000000000;
	sram_mem[66236] = 16'b0000000000000000;
	sram_mem[66237] = 16'b0000000000000000;
	sram_mem[66238] = 16'b0000000000000000;
	sram_mem[66239] = 16'b0000000000000000;
	sram_mem[66240] = 16'b0000000000000000;
	sram_mem[66241] = 16'b0000000000000000;
	sram_mem[66242] = 16'b0000000000000000;
	sram_mem[66243] = 16'b0000000000000000;
	sram_mem[66244] = 16'b0000000000000000;
	sram_mem[66245] = 16'b0000000000000000;
	sram_mem[66246] = 16'b0000000000000000;
	sram_mem[66247] = 16'b0000000000000000;
	sram_mem[66248] = 16'b0000000000000000;
	sram_mem[66249] = 16'b0000000000000000;
	sram_mem[66250] = 16'b0000000000000000;
	sram_mem[66251] = 16'b0000000000000000;
	sram_mem[66252] = 16'b0000000000000000;
	sram_mem[66253] = 16'b0000000000000000;
	sram_mem[66254] = 16'b0000000000000000;
	sram_mem[66255] = 16'b0000000000000000;
	sram_mem[66256] = 16'b0000000000000000;
	sram_mem[66257] = 16'b0000000000000000;
	sram_mem[66258] = 16'b0000000000000000;
	sram_mem[66259] = 16'b0000000000000000;
	sram_mem[66260] = 16'b0000000000000000;
	sram_mem[66261] = 16'b0000000000000000;
	sram_mem[66262] = 16'b0000000000000000;
	sram_mem[66263] = 16'b0000000000000000;
	sram_mem[66264] = 16'b0000000000000000;
	sram_mem[66265] = 16'b0000000000000000;
	sram_mem[66266] = 16'b0000000000000000;
	sram_mem[66267] = 16'b0000000000000000;
	sram_mem[66268] = 16'b0000000000000000;
	sram_mem[66269] = 16'b0000000000000000;
	sram_mem[66270] = 16'b0000000000000000;
	sram_mem[66271] = 16'b0000000000000000;
	sram_mem[66272] = 16'b0000000000000000;
	sram_mem[66273] = 16'b0000000000000000;
	sram_mem[66274] = 16'b0000000000000000;
	sram_mem[66275] = 16'b0000000000000000;
	sram_mem[66276] = 16'b0000000000000000;
	sram_mem[66277] = 16'b0000000000000000;
	sram_mem[66278] = 16'b0000000000000000;
	sram_mem[66279] = 16'b0000000000000000;
	sram_mem[66280] = 16'b0000000000000000;
	sram_mem[66281] = 16'b0000000000000000;
	sram_mem[66282] = 16'b0000000000000000;
	sram_mem[66283] = 16'b0000000000000000;
	sram_mem[66284] = 16'b0000000000000000;
	sram_mem[66285] = 16'b0000000000000000;
	sram_mem[66286] = 16'b0000000000000000;
	sram_mem[66287] = 16'b0000000000000000;
	sram_mem[66288] = 16'b0000000000000000;
	sram_mem[66289] = 16'b0000000000000000;
	sram_mem[66290] = 16'b0000000000000000;
	sram_mem[66291] = 16'b0000000000000000;
	sram_mem[66292] = 16'b0000000000000000;
	sram_mem[66293] = 16'b0000000000000000;
	sram_mem[66294] = 16'b0000000000000000;
	sram_mem[66295] = 16'b0000000000000000;
	sram_mem[66296] = 16'b0000000000000000;
	sram_mem[66297] = 16'b0000000000000000;
	sram_mem[66298] = 16'b0000000000000000;
	sram_mem[66299] = 16'b0000000000000000;
	sram_mem[66300] = 16'b0000000000000000;
	sram_mem[66301] = 16'b0000000000000000;
	sram_mem[66302] = 16'b0000000000000000;
	sram_mem[66303] = 16'b0000000000000000;
	sram_mem[66304] = 16'b0000000000000000;
	sram_mem[66305] = 16'b0000000000000000;
	sram_mem[66306] = 16'b0000000000000000;
	sram_mem[66307] = 16'b0000000000000000;
	sram_mem[66308] = 16'b0000000000000000;
	sram_mem[66309] = 16'b0000000000000000;
	sram_mem[66310] = 16'b0000000000000000;
	sram_mem[66311] = 16'b0000000000000000;
	sram_mem[66312] = 16'b0000000000000000;
	sram_mem[66313] = 16'b0000000000000000;
	sram_mem[66314] = 16'b0000000000000000;
	sram_mem[66315] = 16'b0000000000000000;
	sram_mem[66316] = 16'b0000000000000000;
	sram_mem[66317] = 16'b0000000000000000;
	sram_mem[66318] = 16'b0000000000000000;
	sram_mem[66319] = 16'b0000000000000000;
	sram_mem[66320] = 16'b0000000000000000;
	sram_mem[66321] = 16'b0000000000000000;
	sram_mem[66322] = 16'b0000000000000000;
	sram_mem[66323] = 16'b0000000000000000;
	sram_mem[66324] = 16'b0000000000000000;
	sram_mem[66325] = 16'b0000000000000000;
	sram_mem[66326] = 16'b0000000000000000;
	sram_mem[66327] = 16'b0000000000000000;
	sram_mem[66328] = 16'b0000000000000000;
	sram_mem[66329] = 16'b0000000000000000;
	sram_mem[66330] = 16'b0000000000000000;
	sram_mem[66331] = 16'b0000000000000000;
	sram_mem[66332] = 16'b0000000000000000;
	sram_mem[66333] = 16'b0000000000000000;
	sram_mem[66334] = 16'b0000000000000000;
	sram_mem[66335] = 16'b0000000000000000;
	sram_mem[66336] = 16'b0000000000000000;
	sram_mem[66337] = 16'b0000000000000000;
	sram_mem[66338] = 16'b0000000000000000;
	sram_mem[66339] = 16'b0000000000000000;
	sram_mem[66340] = 16'b0000000000000000;
	sram_mem[66341] = 16'b0000000000000000;
	sram_mem[66342] = 16'b0000000000000000;
	sram_mem[66343] = 16'b0000000000000000;
	sram_mem[66344] = 16'b0000000000000000;
	sram_mem[66345] = 16'b0000000000000000;
	sram_mem[66346] = 16'b0000000000000000;
	sram_mem[66347] = 16'b0000000000000000;
	sram_mem[66348] = 16'b0000000000000000;
	sram_mem[66349] = 16'b0000000000000000;
	sram_mem[66350] = 16'b0000000000000000;
	sram_mem[66351] = 16'b0000000000000000;
	sram_mem[66352] = 16'b0000000000000000;
	sram_mem[66353] = 16'b0000000000000000;
	sram_mem[66354] = 16'b0000000000000000;
	sram_mem[66355] = 16'b0000000000000000;
	sram_mem[66356] = 16'b0000000000000000;
	sram_mem[66357] = 16'b0000000000000000;
	sram_mem[66358] = 16'b0000000000000000;
	sram_mem[66359] = 16'b0000000000000000;
	sram_mem[66360] = 16'b0000000000000000;
	sram_mem[66361] = 16'b0000000000000000;
	sram_mem[66362] = 16'b0000000000000000;
	sram_mem[66363] = 16'b0000000000000000;
	sram_mem[66364] = 16'b0000000000000000;
	sram_mem[66365] = 16'b0000000000000000;
	sram_mem[66366] = 16'b0000000000000000;
	sram_mem[66367] = 16'b0000000000000000;
	sram_mem[66368] = 16'b0000000000000000;
	sram_mem[66369] = 16'b0000000000000000;
	sram_mem[66370] = 16'b0000000000000000;
	sram_mem[66371] = 16'b0000000000000000;
	sram_mem[66372] = 16'b0000000000000000;
	sram_mem[66373] = 16'b0000000000000000;
	sram_mem[66374] = 16'b0000000000000000;
	sram_mem[66375] = 16'b0000000000000000;
	sram_mem[66376] = 16'b0000000000000000;
	sram_mem[66377] = 16'b0000000000000000;
	sram_mem[66378] = 16'b0000000000000000;
	sram_mem[66379] = 16'b0000000000000000;
	sram_mem[66380] = 16'b0000000000000000;
	sram_mem[66381] = 16'b0000000000000000;
	sram_mem[66382] = 16'b0000000000000000;
	sram_mem[66383] = 16'b0000000000000000;
	sram_mem[66384] = 16'b0000000000000000;
	sram_mem[66385] = 16'b0000000000000000;
	sram_mem[66386] = 16'b0000000000000000;
	sram_mem[66387] = 16'b0000000000000000;
	sram_mem[66388] = 16'b0000000000000000;
	sram_mem[66389] = 16'b0000000000000000;
	sram_mem[66390] = 16'b0000000000000000;
	sram_mem[66391] = 16'b0000000000000000;
	sram_mem[66392] = 16'b0000000000000000;
	sram_mem[66393] = 16'b0000000000000000;
	sram_mem[66394] = 16'b0000000000000000;
	sram_mem[66395] = 16'b0000000000000000;
	sram_mem[66396] = 16'b0000000000000000;
	sram_mem[66397] = 16'b0000000000000000;
	sram_mem[66398] = 16'b0000000000000000;
	sram_mem[66399] = 16'b0000000000000000;
	sram_mem[66400] = 16'b0000000000000000;
	sram_mem[66401] = 16'b0000000000000000;
	sram_mem[66402] = 16'b0000000000000000;
	sram_mem[66403] = 16'b0000000000000000;
	sram_mem[66404] = 16'b0000000000000000;
	sram_mem[66405] = 16'b0000000000000000;
	sram_mem[66406] = 16'b0000000000000000;
	sram_mem[66407] = 16'b0000000000000000;
	sram_mem[66408] = 16'b0000000000000000;
	sram_mem[66409] = 16'b0000000000000000;
	sram_mem[66410] = 16'b0000000000000000;
	sram_mem[66411] = 16'b0000000000000000;
	sram_mem[66412] = 16'b0000000000000000;
	sram_mem[66413] = 16'b0000000000000000;
	sram_mem[66414] = 16'b0000000000000000;
	sram_mem[66415] = 16'b0000000000000000;
	sram_mem[66416] = 16'b0000000000000000;
	sram_mem[66417] = 16'b0000000000000000;
	sram_mem[66418] = 16'b0000000000000000;
	sram_mem[66419] = 16'b0000000000000000;
	sram_mem[66420] = 16'b0000000000000000;
	sram_mem[66421] = 16'b0000000000000000;
	sram_mem[66422] = 16'b0000000000000000;
	sram_mem[66423] = 16'b0000000000000000;
	sram_mem[66424] = 16'b0000000000000000;
	sram_mem[66425] = 16'b0000000000000000;
	sram_mem[66426] = 16'b0000000000000000;
	sram_mem[66427] = 16'b0000000000000000;
	sram_mem[66428] = 16'b0000000000000000;
	sram_mem[66429] = 16'b0000000000000000;
	sram_mem[66430] = 16'b0000000000000000;
	sram_mem[66431] = 16'b0000000000000000;
	sram_mem[66432] = 16'b0000000000000000;
	sram_mem[66433] = 16'b0000000000000000;
	sram_mem[66434] = 16'b0000000000000000;
	sram_mem[66435] = 16'b0000000000000000;
	sram_mem[66436] = 16'b0000000000000000;
	sram_mem[66437] = 16'b0000000000000000;
	sram_mem[66438] = 16'b0000000000000000;
	sram_mem[66439] = 16'b0000000000000000;
	sram_mem[66440] = 16'b0000000000000000;
	sram_mem[66441] = 16'b0000000000000000;
	sram_mem[66442] = 16'b0000000000000000;
	sram_mem[66443] = 16'b0000000000000000;
	sram_mem[66444] = 16'b0000000000000000;
	sram_mem[66445] = 16'b0000000000000000;
	sram_mem[66446] = 16'b0000000000000000;
	sram_mem[66447] = 16'b0000000000000000;
	sram_mem[66448] = 16'b0000000000000000;
	sram_mem[66449] = 16'b0000000000000000;
	sram_mem[66450] = 16'b0000000000000000;
	sram_mem[66451] = 16'b0000000000000000;
	sram_mem[66452] = 16'b0000000000000000;
	sram_mem[66453] = 16'b0000000000000000;
	sram_mem[66454] = 16'b0000000000000000;
	sram_mem[66455] = 16'b0000000000000000;
	sram_mem[66456] = 16'b0000000000000000;
	sram_mem[66457] = 16'b0000000000000000;
	sram_mem[66458] = 16'b0000000000000000;
	sram_mem[66459] = 16'b0000000000000000;
	sram_mem[66460] = 16'b0000000000000000;
	sram_mem[66461] = 16'b0000000000000000;
	sram_mem[66462] = 16'b0000000000000000;
	sram_mem[66463] = 16'b0000000000000000;
	sram_mem[66464] = 16'b0000000000000000;
	sram_mem[66465] = 16'b0000000000000000;
	sram_mem[66466] = 16'b0000000000000000;
	sram_mem[66467] = 16'b0000000000000000;
	sram_mem[66468] = 16'b0000000000000000;
	sram_mem[66469] = 16'b0000000000000000;
	sram_mem[66470] = 16'b0000000000000000;
	sram_mem[66471] = 16'b0000000000000000;
	sram_mem[66472] = 16'b0000000000000000;
	sram_mem[66473] = 16'b0000000000000000;
	sram_mem[66474] = 16'b0000000000000000;
	sram_mem[66475] = 16'b0000000000000000;
	sram_mem[66476] = 16'b0000000000000000;
	sram_mem[66477] = 16'b0000000000000000;
	sram_mem[66478] = 16'b0000000000000000;
	sram_mem[66479] = 16'b0000000000000000;
	sram_mem[66480] = 16'b0000000000000000;
	sram_mem[66481] = 16'b0000000000000000;
	sram_mem[66482] = 16'b0000000000000000;
	sram_mem[66483] = 16'b0000000000000000;
	sram_mem[66484] = 16'b0000000000000000;
	sram_mem[66485] = 16'b0000000000000000;
	sram_mem[66486] = 16'b0000000000000000;
	sram_mem[66487] = 16'b0000000000000000;
	sram_mem[66488] = 16'b0000000000000000;
	sram_mem[66489] = 16'b0000000000000000;
	sram_mem[66490] = 16'b0000000000000000;
	sram_mem[66491] = 16'b0000000000000000;
	sram_mem[66492] = 16'b0000000000000000;
	sram_mem[66493] = 16'b0000000000000000;
	sram_mem[66494] = 16'b0000000000000000;
	sram_mem[66495] = 16'b0000000000000000;
	sram_mem[66496] = 16'b0000000000000000;
	sram_mem[66497] = 16'b0000000000000000;
	sram_mem[66498] = 16'b0000000000000000;
	sram_mem[66499] = 16'b0000000000000000;
	sram_mem[66500] = 16'b0000000000000000;
	sram_mem[66501] = 16'b0000000000000000;
	sram_mem[66502] = 16'b0000000000000000;
	sram_mem[66503] = 16'b0000000000000000;
	sram_mem[66504] = 16'b0000000000000000;
	sram_mem[66505] = 16'b0000000000000000;
	sram_mem[66506] = 16'b0000000000000000;
	sram_mem[66507] = 16'b0000000000000000;
	sram_mem[66508] = 16'b0000000000000000;
	sram_mem[66509] = 16'b0000000000000000;
	sram_mem[66510] = 16'b0000000000000000;
	sram_mem[66511] = 16'b0000000000000000;
	sram_mem[66512] = 16'b0000000000000000;
	sram_mem[66513] = 16'b0000000000000000;
	sram_mem[66514] = 16'b0000000000000000;
	sram_mem[66515] = 16'b0000000000000000;
	sram_mem[66516] = 16'b0000000000000000;
	sram_mem[66517] = 16'b0000000000000000;
	sram_mem[66518] = 16'b0000000000000000;
	sram_mem[66519] = 16'b0000000000000000;
	sram_mem[66520] = 16'b0000000000000000;
	sram_mem[66521] = 16'b0000000000000000;
	sram_mem[66522] = 16'b0000000000000000;
	sram_mem[66523] = 16'b0000000000000000;
	sram_mem[66524] = 16'b0000000000000000;
	sram_mem[66525] = 16'b0000000000000000;
	sram_mem[66526] = 16'b0000000000000000;
	sram_mem[66527] = 16'b0000000000000000;
	sram_mem[66528] = 16'b0000000000000000;
	sram_mem[66529] = 16'b0000000000000000;
	sram_mem[66530] = 16'b0000000000000000;
	sram_mem[66531] = 16'b0000000000000000;
	sram_mem[66532] = 16'b0000000000000000;
	sram_mem[66533] = 16'b0000000000000000;
	sram_mem[66534] = 16'b0000000000000000;
	sram_mem[66535] = 16'b0000000000000000;
	sram_mem[66536] = 16'b0000000000000000;
	sram_mem[66537] = 16'b0000000000000000;
	sram_mem[66538] = 16'b0000000000000000;
	sram_mem[66539] = 16'b0000000000000000;
	sram_mem[66540] = 16'b0000000000000000;
	sram_mem[66541] = 16'b0000000000000000;
	sram_mem[66542] = 16'b0000000000000000;
	sram_mem[66543] = 16'b0000000000000000;
	sram_mem[66544] = 16'b0000000000000000;
	sram_mem[66545] = 16'b0000000000000000;
	sram_mem[66546] = 16'b0000000000000000;
	sram_mem[66547] = 16'b0000000000000000;
	sram_mem[66548] = 16'b0000000000000000;
	sram_mem[66549] = 16'b0000000000000000;
	sram_mem[66550] = 16'b0000000000000000;
	sram_mem[66551] = 16'b0000000000000000;
	sram_mem[66552] = 16'b0000000000000000;
	sram_mem[66553] = 16'b0000000000000000;
	sram_mem[66554] = 16'b0000000000000000;
	sram_mem[66555] = 16'b0000000000000000;
	sram_mem[66556] = 16'b0000000000000000;
	sram_mem[66557] = 16'b0000000000000000;
	sram_mem[66558] = 16'b0000000000000000;
	sram_mem[66559] = 16'b0000000000000000;
	sram_mem[66560] = 16'b0000000000000000;
	sram_mem[66561] = 16'b0000000000000000;
	sram_mem[66562] = 16'b0000000000000000;
	sram_mem[66563] = 16'b0000000000000000;
	sram_mem[66564] = 16'b0000000000000000;
	sram_mem[66565] = 16'b0000000000000000;
	sram_mem[66566] = 16'b0000000000000000;
	sram_mem[66567] = 16'b0000000000000000;
	sram_mem[66568] = 16'b0000000000000000;
	sram_mem[66569] = 16'b0000000000000000;
	sram_mem[66570] = 16'b0000000000000000;
	sram_mem[66571] = 16'b0000000000000000;
	sram_mem[66572] = 16'b0000000000000000;
	sram_mem[66573] = 16'b0000000000000000;
	sram_mem[66574] = 16'b0000000000000000;
	sram_mem[66575] = 16'b0000000000000000;
	sram_mem[66576] = 16'b0000000000000000;
	sram_mem[66577] = 16'b0000000000000000;
	sram_mem[66578] = 16'b0000000000000000;
	sram_mem[66579] = 16'b0000000000000000;
	sram_mem[66580] = 16'b0000000000000000;
	sram_mem[66581] = 16'b0000000000000000;
	sram_mem[66582] = 16'b0000000000000000;
	sram_mem[66583] = 16'b0000000000000000;
	sram_mem[66584] = 16'b0000000000000000;
	sram_mem[66585] = 16'b0000000000000000;
	sram_mem[66586] = 16'b0000000000000000;
	sram_mem[66587] = 16'b0000000000000000;
	sram_mem[66588] = 16'b0000000000000000;
	sram_mem[66589] = 16'b0000000000000000;
	sram_mem[66590] = 16'b0000000000000000;
	sram_mem[66591] = 16'b0000000000000000;
	sram_mem[66592] = 16'b0000000000000000;
	sram_mem[66593] = 16'b0000000000000000;
	sram_mem[66594] = 16'b0000000000000000;
	sram_mem[66595] = 16'b0000000000000000;
	sram_mem[66596] = 16'b0000000000000000;
	sram_mem[66597] = 16'b0000000000000000;
	sram_mem[66598] = 16'b0000000000000000;
	sram_mem[66599] = 16'b0000000000000000;
	sram_mem[66600] = 16'b0000000000000000;
	sram_mem[66601] = 16'b0000000000000000;
	sram_mem[66602] = 16'b0000000000000000;
	sram_mem[66603] = 16'b0000000000000000;
	sram_mem[66604] = 16'b0000000000000000;
	sram_mem[66605] = 16'b0000000000000000;
	sram_mem[66606] = 16'b0000000000000000;
	sram_mem[66607] = 16'b0000000000000000;
	sram_mem[66608] = 16'b0000000000000000;
	sram_mem[66609] = 16'b0000000000000000;
	sram_mem[66610] = 16'b0000000000000000;
	sram_mem[66611] = 16'b0000000000000000;
	sram_mem[66612] = 16'b0000000000000000;
	sram_mem[66613] = 16'b0000000000000000;
	sram_mem[66614] = 16'b0000000000000000;
	sram_mem[66615] = 16'b0000000000000000;
	sram_mem[66616] = 16'b0000000000000000;
	sram_mem[66617] = 16'b0000000000000000;
	sram_mem[66618] = 16'b0000000000000000;
	sram_mem[66619] = 16'b0000000000000000;
	sram_mem[66620] = 16'b0000000000000000;
	sram_mem[66621] = 16'b0000000000000000;
	sram_mem[66622] = 16'b0000000000000000;
	sram_mem[66623] = 16'b0000000000000000;
	sram_mem[66624] = 16'b0000000000000000;
	sram_mem[66625] = 16'b0000000000000000;
	sram_mem[66626] = 16'b0000000000000000;
	sram_mem[66627] = 16'b0000000000000000;
	sram_mem[66628] = 16'b0000000000000000;
	sram_mem[66629] = 16'b0000000000000000;
	sram_mem[66630] = 16'b0000000000000000;
	sram_mem[66631] = 16'b0000000000000000;
	sram_mem[66632] = 16'b0000000000000000;
	sram_mem[66633] = 16'b0000000000000000;
	sram_mem[66634] = 16'b0000000000000000;
	sram_mem[66635] = 16'b0000000000000000;
	sram_mem[66636] = 16'b0000000000000000;
	sram_mem[66637] = 16'b0000000000000000;
	sram_mem[66638] = 16'b0000000000000000;
	sram_mem[66639] = 16'b0000000000000000;
	sram_mem[66640] = 16'b0000000000000000;
	sram_mem[66641] = 16'b0000000000000000;
	sram_mem[66642] = 16'b0000000000000000;
	sram_mem[66643] = 16'b0000000000000000;
	sram_mem[66644] = 16'b0000000000000000;
	sram_mem[66645] = 16'b0000000000000000;
	sram_mem[66646] = 16'b0000000000000000;
	sram_mem[66647] = 16'b0000000000000000;
	sram_mem[66648] = 16'b0000000000000000;
	sram_mem[66649] = 16'b0000000000000000;
	sram_mem[66650] = 16'b0000000000000000;
	sram_mem[66651] = 16'b0000000000000000;
	sram_mem[66652] = 16'b0000000000000000;
	sram_mem[66653] = 16'b0000000000000000;
	sram_mem[66654] = 16'b0000000000000000;
	sram_mem[66655] = 16'b0000000000000000;
	sram_mem[66656] = 16'b0000000000000000;
	sram_mem[66657] = 16'b0000000000000000;
	sram_mem[66658] = 16'b0000000000000000;
	sram_mem[66659] = 16'b0000000000000000;
	sram_mem[66660] = 16'b0000000000000000;
	sram_mem[66661] = 16'b0000000000000000;
	sram_mem[66662] = 16'b0000000000000000;
	sram_mem[66663] = 16'b0000000000000000;
	sram_mem[66664] = 16'b0000000000000000;
	sram_mem[66665] = 16'b0000000000000000;
	sram_mem[66666] = 16'b0000000000000000;
	sram_mem[66667] = 16'b0000000000000000;
	sram_mem[66668] = 16'b0000000000000000;
	sram_mem[66669] = 16'b0000000000000000;
	sram_mem[66670] = 16'b0000000000000000;
	sram_mem[66671] = 16'b0000000000000000;
	sram_mem[66672] = 16'b0000000000000000;
	sram_mem[66673] = 16'b0000000000000000;
	sram_mem[66674] = 16'b0000000000000000;
	sram_mem[66675] = 16'b0000000000000000;
	sram_mem[66676] = 16'b0000000000000000;
	sram_mem[66677] = 16'b0000000000000000;
	sram_mem[66678] = 16'b0000000000000000;
	sram_mem[66679] = 16'b0000000000000000;
	sram_mem[66680] = 16'b0000000000000000;
	sram_mem[66681] = 16'b0000000000000000;
	sram_mem[66682] = 16'b0000000000000000;
	sram_mem[66683] = 16'b0000000000000000;
	sram_mem[66684] = 16'b0000000000000000;
	sram_mem[66685] = 16'b0000000000000000;
	sram_mem[66686] = 16'b0000000000000000;
	sram_mem[66687] = 16'b0000000000000000;
	sram_mem[66688] = 16'b0000000000000000;
	sram_mem[66689] = 16'b0000000000000000;
	sram_mem[66690] = 16'b0000000000000000;
	sram_mem[66691] = 16'b0000000000000000;
	sram_mem[66692] = 16'b0000000000000000;
	sram_mem[66693] = 16'b0000000000000000;
	sram_mem[66694] = 16'b0000000000000000;
	sram_mem[66695] = 16'b0000000000000000;
	sram_mem[66696] = 16'b0000000000000000;
	sram_mem[66697] = 16'b0000000000000000;
	sram_mem[66698] = 16'b0000000000000000;
	sram_mem[66699] = 16'b0000000000000000;
	sram_mem[66700] = 16'b0000000000000000;
	sram_mem[66701] = 16'b0000000000000000;
	sram_mem[66702] = 16'b0000000000000000;
	sram_mem[66703] = 16'b0000000000000000;
	sram_mem[66704] = 16'b0000000000000000;
	sram_mem[66705] = 16'b0000000000000000;
	sram_mem[66706] = 16'b0000000000000000;
	sram_mem[66707] = 16'b0000000000000000;
	sram_mem[66708] = 16'b0000000000000000;
	sram_mem[66709] = 16'b0000000000000000;
	sram_mem[66710] = 16'b0000000000000000;
	sram_mem[66711] = 16'b0000000000000000;
	sram_mem[66712] = 16'b0000000000000000;
	sram_mem[66713] = 16'b0000000000000000;
	sram_mem[66714] = 16'b0000000000000000;
	sram_mem[66715] = 16'b0000000000000000;
	sram_mem[66716] = 16'b0000000000000000;
	sram_mem[66717] = 16'b0000000000000000;
	sram_mem[66718] = 16'b0000000000000000;
	sram_mem[66719] = 16'b0000000000000000;
	sram_mem[66720] = 16'b0000000000000000;
	sram_mem[66721] = 16'b0000000000000000;
	sram_mem[66722] = 16'b0000000000000000;
	sram_mem[66723] = 16'b0000000000000000;
	sram_mem[66724] = 16'b0000000000000000;
	sram_mem[66725] = 16'b0000000000000000;
	sram_mem[66726] = 16'b0000000000000000;
	sram_mem[66727] = 16'b0000000000000000;
	sram_mem[66728] = 16'b0000000000000000;
	sram_mem[66729] = 16'b0000000000000000;
	sram_mem[66730] = 16'b0000000000000000;
	sram_mem[66731] = 16'b0000000000000000;
	sram_mem[66732] = 16'b0000000000000000;
	sram_mem[66733] = 16'b0000000000000000;
	sram_mem[66734] = 16'b0000000000000000;
	sram_mem[66735] = 16'b0000000000000000;
	sram_mem[66736] = 16'b0000000000000000;
	sram_mem[66737] = 16'b0000000000000000;
	sram_mem[66738] = 16'b0000000000000000;
	sram_mem[66739] = 16'b0000000000000000;
	sram_mem[66740] = 16'b0000000000000000;
	sram_mem[66741] = 16'b0000000000000000;
	sram_mem[66742] = 16'b0000000000000000;
	sram_mem[66743] = 16'b0000000000000000;
	sram_mem[66744] = 16'b0000000000000000;
	sram_mem[66745] = 16'b0000000000000000;
	sram_mem[66746] = 16'b0000000000000000;
	sram_mem[66747] = 16'b0000000000000000;
	sram_mem[66748] = 16'b0000000000000000;
	sram_mem[66749] = 16'b0000000000000000;
	sram_mem[66750] = 16'b0000000000000000;
	sram_mem[66751] = 16'b0000000000000000;
	sram_mem[66752] = 16'b0000000000000000;
	sram_mem[66753] = 16'b0000000000000000;
	sram_mem[66754] = 16'b0000000000000000;
	sram_mem[66755] = 16'b0000000000000000;
	sram_mem[66756] = 16'b0000000000000000;
	sram_mem[66757] = 16'b0000000000000000;
	sram_mem[66758] = 16'b0000000000000000;
	sram_mem[66759] = 16'b0000000000000000;
	sram_mem[66760] = 16'b0000000000000000;
	sram_mem[66761] = 16'b0000000000000000;
	sram_mem[66762] = 16'b0000000000000000;
	sram_mem[66763] = 16'b0000000000000000;
	sram_mem[66764] = 16'b0000000000000000;
	sram_mem[66765] = 16'b0000000000000000;
	sram_mem[66766] = 16'b0000000000000000;
	sram_mem[66767] = 16'b0000000000000000;
	sram_mem[66768] = 16'b0000000000000000;
	sram_mem[66769] = 16'b0000000000000000;
	sram_mem[66770] = 16'b0000000000000000;
	sram_mem[66771] = 16'b0000000000000000;
	sram_mem[66772] = 16'b0000000000000000;
	sram_mem[66773] = 16'b0000000000000000;
	sram_mem[66774] = 16'b0000000000000000;
	sram_mem[66775] = 16'b0000000000000000;
	sram_mem[66776] = 16'b0000000000000000;
	sram_mem[66777] = 16'b0000000000000000;
	sram_mem[66778] = 16'b0000000000000000;
	sram_mem[66779] = 16'b0000000000000000;
	sram_mem[66780] = 16'b0000000000000000;
	sram_mem[66781] = 16'b0000000000000000;
	sram_mem[66782] = 16'b0000000000000000;
	sram_mem[66783] = 16'b0000000000000000;
	sram_mem[66784] = 16'b0000000000000000;
	sram_mem[66785] = 16'b0000000000000000;
	sram_mem[66786] = 16'b0000000000000000;
	sram_mem[66787] = 16'b0000000000000000;
	sram_mem[66788] = 16'b0000000000000000;
	sram_mem[66789] = 16'b0000000000000000;
	sram_mem[66790] = 16'b0000000000000000;
	sram_mem[66791] = 16'b0000000000000000;
	sram_mem[66792] = 16'b0000000000000000;
	sram_mem[66793] = 16'b0000000000000000;
	sram_mem[66794] = 16'b0000000000000000;
	sram_mem[66795] = 16'b0000000000000000;
	sram_mem[66796] = 16'b0000000000000000;
	sram_mem[66797] = 16'b0000000000000000;
	sram_mem[66798] = 16'b0000000000000000;
	sram_mem[66799] = 16'b0000000000000000;
	sram_mem[66800] = 16'b0000000000000000;
	sram_mem[66801] = 16'b0000000000000000;
	sram_mem[66802] = 16'b0000000000000000;
	sram_mem[66803] = 16'b0000000000000000;
	sram_mem[66804] = 16'b0000000000000000;
	sram_mem[66805] = 16'b0000000000000000;
	sram_mem[66806] = 16'b0000000000000000;
	sram_mem[66807] = 16'b0000000000000000;
	sram_mem[66808] = 16'b0000000000000000;
	sram_mem[66809] = 16'b0000000000000000;
	sram_mem[66810] = 16'b0000000000000000;
	sram_mem[66811] = 16'b0000000000000000;
	sram_mem[66812] = 16'b0000000000000000;
	sram_mem[66813] = 16'b0000000000000000;
	sram_mem[66814] = 16'b0000000000000000;
	sram_mem[66815] = 16'b0000000000000000;
	sram_mem[66816] = 16'b0000000000000000;
	sram_mem[66817] = 16'b0000000000000000;
	sram_mem[66818] = 16'b0000000000000000;
	sram_mem[66819] = 16'b0000000000000000;
	sram_mem[66820] = 16'b0000000000000000;
	sram_mem[66821] = 16'b0000000000000000;
	sram_mem[66822] = 16'b0000000000000000;
	sram_mem[66823] = 16'b0000000000000000;
	sram_mem[66824] = 16'b0000000000000000;
	sram_mem[66825] = 16'b0000000000000000;
	sram_mem[66826] = 16'b0000000000000000;
	sram_mem[66827] = 16'b0000000000000000;
	sram_mem[66828] = 16'b0000000000000000;
	sram_mem[66829] = 16'b0000000000000000;
	sram_mem[66830] = 16'b0000000000000000;
	sram_mem[66831] = 16'b0000000000000000;
	sram_mem[66832] = 16'b0000000000000000;
	sram_mem[66833] = 16'b0000000000000000;
	sram_mem[66834] = 16'b0000000000000000;
	sram_mem[66835] = 16'b0000000000000000;
	sram_mem[66836] = 16'b0000000000000000;
	sram_mem[66837] = 16'b0000000000000000;
	sram_mem[66838] = 16'b0000000000000000;
	sram_mem[66839] = 16'b0000000000000000;
	sram_mem[66840] = 16'b0000000000000000;
	sram_mem[66841] = 16'b0000000000000000;
	sram_mem[66842] = 16'b0000000000000000;
	sram_mem[66843] = 16'b0000000000000000;
	sram_mem[66844] = 16'b0000000000000000;
	sram_mem[66845] = 16'b0000000000000000;
	sram_mem[66846] = 16'b0000000000000000;
	sram_mem[66847] = 16'b0000000000000000;
	sram_mem[66848] = 16'b0000000000000000;
	sram_mem[66849] = 16'b0000000000000000;
	sram_mem[66850] = 16'b0000000000000000;
	sram_mem[66851] = 16'b0000000000000000;
	sram_mem[66852] = 16'b0000000000000000;
	sram_mem[66853] = 16'b0000000000000000;
	sram_mem[66854] = 16'b0000000000000000;
	sram_mem[66855] = 16'b0000000000000000;
	sram_mem[66856] = 16'b0000000000000000;
	sram_mem[66857] = 16'b0000000000000000;
	sram_mem[66858] = 16'b0000000000000000;
	sram_mem[66859] = 16'b0000000000000000;
	sram_mem[66860] = 16'b0000000000000000;
	sram_mem[66861] = 16'b0000000000000000;
	sram_mem[66862] = 16'b0000000000000000;
	sram_mem[66863] = 16'b0000000000000000;
	sram_mem[66864] = 16'b0000000000000000;
	sram_mem[66865] = 16'b0000000000000000;
	sram_mem[66866] = 16'b0000000000000000;
	sram_mem[66867] = 16'b0000000000000000;
	sram_mem[66868] = 16'b0000000000000000;
	sram_mem[66869] = 16'b0000000000000000;
	sram_mem[66870] = 16'b0000000000000000;
	sram_mem[66871] = 16'b0000000000000000;
	sram_mem[66872] = 16'b0000000000000000;
	sram_mem[66873] = 16'b0000000000000000;
	sram_mem[66874] = 16'b0000000000000000;
	sram_mem[66875] = 16'b0000000000000000;
	sram_mem[66876] = 16'b0000000000000000;
	sram_mem[66877] = 16'b0000000000000000;
	sram_mem[66878] = 16'b0000000000000000;
	sram_mem[66879] = 16'b0000000000000000;
	sram_mem[66880] = 16'b0000000000000000;
	sram_mem[66881] = 16'b0000000000000000;
	sram_mem[66882] = 16'b0000000000000000;
	sram_mem[66883] = 16'b0000000000000000;
	sram_mem[66884] = 16'b0000000000000000;
	sram_mem[66885] = 16'b0000000000000000;
	sram_mem[66886] = 16'b0000000000000000;
	sram_mem[66887] = 16'b0000000000000000;
	sram_mem[66888] = 16'b0000000000000000;
	sram_mem[66889] = 16'b0000000000000000;
	sram_mem[66890] = 16'b0000000000000000;
	sram_mem[66891] = 16'b0000000000000000;
	sram_mem[66892] = 16'b0000000000000000;
	sram_mem[66893] = 16'b0000000000000000;
	sram_mem[66894] = 16'b0000000000000000;
	sram_mem[66895] = 16'b0000000000000000;
	sram_mem[66896] = 16'b0000000000000000;
	sram_mem[66897] = 16'b0000000000000000;
	sram_mem[66898] = 16'b0000000000000000;
	sram_mem[66899] = 16'b0000000000000000;
	sram_mem[66900] = 16'b0000000000000000;
	sram_mem[66901] = 16'b0000000000000000;
	sram_mem[66902] = 16'b0000000000000000;
	sram_mem[66903] = 16'b0000000000000000;
	sram_mem[66904] = 16'b0000000000000000;
	sram_mem[66905] = 16'b0000000000000000;
	sram_mem[66906] = 16'b0000000000000000;
	sram_mem[66907] = 16'b0000000000000000;
	sram_mem[66908] = 16'b0000000000000000;
	sram_mem[66909] = 16'b0000000000000000;
	sram_mem[66910] = 16'b0000000000000000;
	sram_mem[66911] = 16'b0000000000000000;
	sram_mem[66912] = 16'b0000000000000000;
	sram_mem[66913] = 16'b0000000000000000;
	sram_mem[66914] = 16'b0000000000000000;
	sram_mem[66915] = 16'b0000000000000000;
	sram_mem[66916] = 16'b0000000000000000;
	sram_mem[66917] = 16'b0000000000000000;
	sram_mem[66918] = 16'b0000000000000000;
	sram_mem[66919] = 16'b0000000000000000;
	sram_mem[66920] = 16'b0000000000000000;
	sram_mem[66921] = 16'b0000000000000000;
	sram_mem[66922] = 16'b0000000000000000;
	sram_mem[66923] = 16'b0000000000000000;
	sram_mem[66924] = 16'b0000000000000000;
	sram_mem[66925] = 16'b0000000000000000;
	sram_mem[66926] = 16'b0000000000000000;
	sram_mem[66927] = 16'b0000000000000000;
	sram_mem[66928] = 16'b0000000000000000;
	sram_mem[66929] = 16'b0000000000000000;
	sram_mem[66930] = 16'b0000000000000000;
	sram_mem[66931] = 16'b0000000000000000;
	sram_mem[66932] = 16'b0000000000000000;
	sram_mem[66933] = 16'b0000000000000000;
	sram_mem[66934] = 16'b0000000000000000;
	sram_mem[66935] = 16'b0000000000000000;
	sram_mem[66936] = 16'b0000000000000000;
	sram_mem[66937] = 16'b0000000000000000;
	sram_mem[66938] = 16'b0000000000000000;
	sram_mem[66939] = 16'b0000000000000000;
	sram_mem[66940] = 16'b0000000000000000;
	sram_mem[66941] = 16'b0000000000000000;
	sram_mem[66942] = 16'b0000000000000000;
	sram_mem[66943] = 16'b0000000000000000;
	sram_mem[66944] = 16'b0000000000000000;
	sram_mem[66945] = 16'b0000000000000000;
	sram_mem[66946] = 16'b0000000000000000;
	sram_mem[66947] = 16'b0000000000000000;
	sram_mem[66948] = 16'b0000000000000000;
	sram_mem[66949] = 16'b0000000000000000;
	sram_mem[66950] = 16'b0000000000000000;
	sram_mem[66951] = 16'b0000000000000000;
	sram_mem[66952] = 16'b0000000000000000;
	sram_mem[66953] = 16'b0000000000000000;
	sram_mem[66954] = 16'b0000000000000000;
	sram_mem[66955] = 16'b0000000000000000;
	sram_mem[66956] = 16'b0000000000000000;
	sram_mem[66957] = 16'b0000000000000000;
	sram_mem[66958] = 16'b0000000000000000;
	sram_mem[66959] = 16'b0000000000000000;
	sram_mem[66960] = 16'b0000000000000000;
	sram_mem[66961] = 16'b0000000000000000;
	sram_mem[66962] = 16'b0000000000000000;
	sram_mem[66963] = 16'b0000000000000000;
	sram_mem[66964] = 16'b0000000000000000;
	sram_mem[66965] = 16'b0000000000000000;
	sram_mem[66966] = 16'b0000000000000000;
	sram_mem[66967] = 16'b0000000000000000;
	sram_mem[66968] = 16'b0000000000000000;
	sram_mem[66969] = 16'b0000000000000000;
	sram_mem[66970] = 16'b0000000000000000;
	sram_mem[66971] = 16'b0000000000000000;
	sram_mem[66972] = 16'b0000000000000000;
	sram_mem[66973] = 16'b0000000000000000;
	sram_mem[66974] = 16'b0000000000000000;
	sram_mem[66975] = 16'b0000000000000000;
	sram_mem[66976] = 16'b0000000000000000;
	sram_mem[66977] = 16'b0000000000000000;
	sram_mem[66978] = 16'b0000000000000000;
	sram_mem[66979] = 16'b0000000000000000;
	sram_mem[66980] = 16'b0000000000000000;
	sram_mem[66981] = 16'b0000000000000000;
	sram_mem[66982] = 16'b0000000000000000;
	sram_mem[66983] = 16'b0000000000000000;
	sram_mem[66984] = 16'b0000000000000000;
	sram_mem[66985] = 16'b0000000000000000;
	sram_mem[66986] = 16'b0000000000000000;
	sram_mem[66987] = 16'b0000000000000000;
	sram_mem[66988] = 16'b0000000000000000;
	sram_mem[66989] = 16'b0000000000000000;
	sram_mem[66990] = 16'b0000000000000000;
	sram_mem[66991] = 16'b0000000000000000;
	sram_mem[66992] = 16'b0000000000000000;
	sram_mem[66993] = 16'b0000000000000000;
	sram_mem[66994] = 16'b0000000000000000;
	sram_mem[66995] = 16'b0000000000000000;
	sram_mem[66996] = 16'b0000000000000000;
	sram_mem[66997] = 16'b0000000000000000;
	sram_mem[66998] = 16'b0000000000000000;
	sram_mem[66999] = 16'b0000000000000000;
	sram_mem[67000] = 16'b0000000000000000;
	sram_mem[67001] = 16'b0000000000000000;
	sram_mem[67002] = 16'b0000000000000000;
	sram_mem[67003] = 16'b0000000000000000;
	sram_mem[67004] = 16'b0000000000000000;
	sram_mem[67005] = 16'b0000000000000000;
	sram_mem[67006] = 16'b0000000000000000;
	sram_mem[67007] = 16'b0000000000000000;
	sram_mem[67008] = 16'b0000000000000000;
	sram_mem[67009] = 16'b0000000000000000;
	sram_mem[67010] = 16'b0000000000000000;
	sram_mem[67011] = 16'b0000000000000000;
	sram_mem[67012] = 16'b0000000000000000;
	sram_mem[67013] = 16'b0000000000000000;
	sram_mem[67014] = 16'b0000000000000000;
	sram_mem[67015] = 16'b0000000000000000;
	sram_mem[67016] = 16'b0000000000000000;
	sram_mem[67017] = 16'b0000000000000000;
	sram_mem[67018] = 16'b0000000000000000;
	sram_mem[67019] = 16'b0000000000000000;
	sram_mem[67020] = 16'b0000000000000000;
	sram_mem[67021] = 16'b0000000000000000;
	sram_mem[67022] = 16'b0000000000000000;
	sram_mem[67023] = 16'b0000000000000000;
	sram_mem[67024] = 16'b0000000000000000;
	sram_mem[67025] = 16'b0000000000000000;
	sram_mem[67026] = 16'b0000000000000000;
	sram_mem[67027] = 16'b0000000000000000;
	sram_mem[67028] = 16'b0000000000000000;
	sram_mem[67029] = 16'b0000000000000000;
	sram_mem[67030] = 16'b0000000000000000;
	sram_mem[67031] = 16'b0000000000000000;
	sram_mem[67032] = 16'b0000000000000000;
	sram_mem[67033] = 16'b0000000000000000;
	sram_mem[67034] = 16'b0000000000000000;
	sram_mem[67035] = 16'b0000000000000000;
	sram_mem[67036] = 16'b0000000000000000;
	sram_mem[67037] = 16'b0000000000000000;
	sram_mem[67038] = 16'b0000000000000000;
	sram_mem[67039] = 16'b0000000000000000;
	sram_mem[67040] = 16'b0000000000000000;
	sram_mem[67041] = 16'b0000000000000000;
	sram_mem[67042] = 16'b0000000000000000;
	sram_mem[67043] = 16'b0000000000000000;
	sram_mem[67044] = 16'b0000000000000000;
	sram_mem[67045] = 16'b0000000000000000;
	sram_mem[67046] = 16'b0000000000000000;
	sram_mem[67047] = 16'b0000000000000000;
	sram_mem[67048] = 16'b0000000000000000;
	sram_mem[67049] = 16'b0000000000000000;
	sram_mem[67050] = 16'b0000000000000000;
	sram_mem[67051] = 16'b0000000000000000;
	sram_mem[67052] = 16'b0000000000000000;
	sram_mem[67053] = 16'b0000000000000000;
	sram_mem[67054] = 16'b0000000000000000;
	sram_mem[67055] = 16'b0000000000000000;
	sram_mem[67056] = 16'b0000000000000000;
	sram_mem[67057] = 16'b0000000000000000;
	sram_mem[67058] = 16'b0000000000000000;
	sram_mem[67059] = 16'b0000000000000000;
	sram_mem[67060] = 16'b0000000000000000;
	sram_mem[67061] = 16'b0000000000000000;
	sram_mem[67062] = 16'b0000000000000000;
	sram_mem[67063] = 16'b0000000000000000;
	sram_mem[67064] = 16'b0000000000000000;
	sram_mem[67065] = 16'b0000000000000000;
	sram_mem[67066] = 16'b0000000000000000;
	sram_mem[67067] = 16'b0000000000000000;
	sram_mem[67068] = 16'b0000000000000000;
	sram_mem[67069] = 16'b0000000000000000;
	sram_mem[67070] = 16'b0000000000000000;
	sram_mem[67071] = 16'b0000000000000000;
	sram_mem[67072] = 16'b0000000000000000;
	sram_mem[67073] = 16'b0000000000000000;
	sram_mem[67074] = 16'b0000000000000000;
	sram_mem[67075] = 16'b0000000000000000;
	sram_mem[67076] = 16'b0000000000000000;
	sram_mem[67077] = 16'b0000000000000000;
	sram_mem[67078] = 16'b0000000000000000;
	sram_mem[67079] = 16'b0000000000000000;
	sram_mem[67080] = 16'b0000000000000000;
	sram_mem[67081] = 16'b0000000000000000;
	sram_mem[67082] = 16'b0000000000000000;
	sram_mem[67083] = 16'b0000000000000000;
	sram_mem[67084] = 16'b0000000000000000;
	sram_mem[67085] = 16'b0000000000000000;
	sram_mem[67086] = 16'b0000000000000000;
	sram_mem[67087] = 16'b0000000000000000;
	sram_mem[67088] = 16'b0000000000000000;
	sram_mem[67089] = 16'b0000000000000000;
	sram_mem[67090] = 16'b0000000000000000;
	sram_mem[67091] = 16'b0000000000000000;
	sram_mem[67092] = 16'b0000000000000000;
	sram_mem[67093] = 16'b0000000000000000;
	sram_mem[67094] = 16'b0000000000000000;
	sram_mem[67095] = 16'b0000000000000000;
	sram_mem[67096] = 16'b0000000000000000;
	sram_mem[67097] = 16'b0000000000000000;
	sram_mem[67098] = 16'b0000000000000000;
	sram_mem[67099] = 16'b0000000000000000;
	sram_mem[67100] = 16'b0000000000000000;
	sram_mem[67101] = 16'b0000000000000000;
	sram_mem[67102] = 16'b0000000000000000;
	sram_mem[67103] = 16'b0000000000000000;
	sram_mem[67104] = 16'b0000000000000000;
	sram_mem[67105] = 16'b0000000000000000;
	sram_mem[67106] = 16'b0000000000000000;
	sram_mem[67107] = 16'b0000000000000000;
	sram_mem[67108] = 16'b0000000000000000;
	sram_mem[67109] = 16'b0000000000000000;
	sram_mem[67110] = 16'b0000000000000000;
	sram_mem[67111] = 16'b0000000000000000;
	sram_mem[67112] = 16'b0000000000000000;
	sram_mem[67113] = 16'b0000000000000000;
	sram_mem[67114] = 16'b0000000000000000;
	sram_mem[67115] = 16'b0000000000000000;
	sram_mem[67116] = 16'b0000000000000000;
	sram_mem[67117] = 16'b0000000000000000;
	sram_mem[67118] = 16'b0000000000000000;
	sram_mem[67119] = 16'b0000000000000000;
	sram_mem[67120] = 16'b0000000000000000;
	sram_mem[67121] = 16'b0000000000000000;
	sram_mem[67122] = 16'b0000000000000000;
	sram_mem[67123] = 16'b0000000000000000;
	sram_mem[67124] = 16'b0000000000000000;
	sram_mem[67125] = 16'b0000000000000000;
	sram_mem[67126] = 16'b0000000000000000;
	sram_mem[67127] = 16'b0000000000000000;
	sram_mem[67128] = 16'b0000000000000000;
	sram_mem[67129] = 16'b0000000000000000;
	sram_mem[67130] = 16'b0000000000000000;
	sram_mem[67131] = 16'b0000000000000000;
	sram_mem[67132] = 16'b0000000000000000;
	sram_mem[67133] = 16'b0000000000000000;
	sram_mem[67134] = 16'b0000000000000000;
	sram_mem[67135] = 16'b0000000000000000;
	sram_mem[67136] = 16'b0000000000000000;
	sram_mem[67137] = 16'b0000000000000000;
	sram_mem[67138] = 16'b0000000000000000;
	sram_mem[67139] = 16'b0000000000000000;
	sram_mem[67140] = 16'b0000000000000000;
	sram_mem[67141] = 16'b0000000000000000;
	sram_mem[67142] = 16'b0000000000000000;
	sram_mem[67143] = 16'b0000000000000000;
	sram_mem[67144] = 16'b0000000000000000;
	sram_mem[67145] = 16'b0000000000000000;
	sram_mem[67146] = 16'b0000000000000000;
	sram_mem[67147] = 16'b0000000000000000;
	sram_mem[67148] = 16'b0000000000000000;
	sram_mem[67149] = 16'b0000000000000000;
	sram_mem[67150] = 16'b0000000000000000;
	sram_mem[67151] = 16'b0000000000000000;
	sram_mem[67152] = 16'b0000000000000000;
	sram_mem[67153] = 16'b0000000000000000;
	sram_mem[67154] = 16'b0000000000000000;
	sram_mem[67155] = 16'b0000000000000000;
	sram_mem[67156] = 16'b0000000000000000;
	sram_mem[67157] = 16'b0000000000000000;
	sram_mem[67158] = 16'b0000000000000000;
	sram_mem[67159] = 16'b0000000000000000;
	sram_mem[67160] = 16'b0000000000000000;
	sram_mem[67161] = 16'b0000000000000000;
	sram_mem[67162] = 16'b0000000000000000;
	sram_mem[67163] = 16'b0000000000000000;
	sram_mem[67164] = 16'b0000000000000000;
	sram_mem[67165] = 16'b0000000000000000;
	sram_mem[67166] = 16'b0000000000000000;
	sram_mem[67167] = 16'b0000000000000000;
	sram_mem[67168] = 16'b0000000000000000;
	sram_mem[67169] = 16'b0000000000000000;
	sram_mem[67170] = 16'b0000000000000000;
	sram_mem[67171] = 16'b0000000000000000;
	sram_mem[67172] = 16'b0000000000000000;
	sram_mem[67173] = 16'b0000000000000000;
	sram_mem[67174] = 16'b0000000000000000;
	sram_mem[67175] = 16'b0000000000000000;
	sram_mem[67176] = 16'b0000000000000000;
	sram_mem[67177] = 16'b0000000000000000;
	sram_mem[67178] = 16'b0000000000000000;
	sram_mem[67179] = 16'b0000000000000000;
	sram_mem[67180] = 16'b0000000000000000;
	sram_mem[67181] = 16'b0000000000000000;
	sram_mem[67182] = 16'b0000000000000000;
	sram_mem[67183] = 16'b0000000000000000;
	sram_mem[67184] = 16'b0000000000000000;
	sram_mem[67185] = 16'b0000000000000000;
	sram_mem[67186] = 16'b0000000000000000;
	sram_mem[67187] = 16'b0000000000000000;
	sram_mem[67188] = 16'b0000000000000000;
	sram_mem[67189] = 16'b0000000000000000;
	sram_mem[67190] = 16'b0000000000000000;
	sram_mem[67191] = 16'b0000000000000000;
	sram_mem[67192] = 16'b0000000000000000;
	sram_mem[67193] = 16'b0000000000000000;
	sram_mem[67194] = 16'b0000000000000000;
	sram_mem[67195] = 16'b0000000000000000;
	sram_mem[67196] = 16'b0000000000000000;
	sram_mem[67197] = 16'b0000000000000000;
	sram_mem[67198] = 16'b0000000000000000;
	sram_mem[67199] = 16'b0000000000000000;
	sram_mem[67200] = 16'b0000000000000000;
	sram_mem[67201] = 16'b0000000000000000;
	sram_mem[67202] = 16'b0000000000000000;
	sram_mem[67203] = 16'b0000000000000000;
	sram_mem[67204] = 16'b0000000000000000;
	sram_mem[67205] = 16'b0000000000000000;
	sram_mem[67206] = 16'b0000000000000000;
	sram_mem[67207] = 16'b0000000000000000;
	sram_mem[67208] = 16'b0000000000000000;
	sram_mem[67209] = 16'b0000000000000000;
	sram_mem[67210] = 16'b0000000000000000;
	sram_mem[67211] = 16'b0000000000000000;
	sram_mem[67212] = 16'b0000000000000000;
	sram_mem[67213] = 16'b0000000000000000;
	sram_mem[67214] = 16'b0000000000000000;
	sram_mem[67215] = 16'b0000000000000000;
	sram_mem[67216] = 16'b0000000000000000;
	sram_mem[67217] = 16'b0000000000000000;
	sram_mem[67218] = 16'b0000000000000000;
	sram_mem[67219] = 16'b0000000000000000;
	sram_mem[67220] = 16'b0000000000000000;
	sram_mem[67221] = 16'b0000000000000000;
	sram_mem[67222] = 16'b0000000000000000;
	sram_mem[67223] = 16'b0000000000000000;
	sram_mem[67224] = 16'b0000000000000000;
	sram_mem[67225] = 16'b0000000000000000;
	sram_mem[67226] = 16'b0000000000000000;
	sram_mem[67227] = 16'b0000000000000000;
	sram_mem[67228] = 16'b0000000000000000;
	sram_mem[67229] = 16'b0000000000000000;
	sram_mem[67230] = 16'b0000000000000000;
	sram_mem[67231] = 16'b0000000000000000;
	sram_mem[67232] = 16'b0000000000000000;
	sram_mem[67233] = 16'b0000000000000000;
	sram_mem[67234] = 16'b0000000000000000;
	sram_mem[67235] = 16'b0000000000000000;
	sram_mem[67236] = 16'b0000000000000000;
	sram_mem[67237] = 16'b0000000000000000;
	sram_mem[67238] = 16'b0000000000000000;
	sram_mem[67239] = 16'b0000000000000000;
	sram_mem[67240] = 16'b0000000000000000;
	sram_mem[67241] = 16'b0000000000000000;
	sram_mem[67242] = 16'b0000000000000000;
	sram_mem[67243] = 16'b0000000000000000;
	sram_mem[67244] = 16'b0000000000000000;
	sram_mem[67245] = 16'b0000000000000000;
	sram_mem[67246] = 16'b0000000000000000;
	sram_mem[67247] = 16'b0000000000000000;
	sram_mem[67248] = 16'b0000000000000000;
	sram_mem[67249] = 16'b0000000000000000;
	sram_mem[67250] = 16'b0000000000000000;
	sram_mem[67251] = 16'b0000000000000000;
	sram_mem[67252] = 16'b0000000000000000;
	sram_mem[67253] = 16'b0000000000000000;
	sram_mem[67254] = 16'b0000000000000000;
	sram_mem[67255] = 16'b0000000000000000;
	sram_mem[67256] = 16'b0000000000000000;
	sram_mem[67257] = 16'b0000000000000000;
	sram_mem[67258] = 16'b0000000000000000;
	sram_mem[67259] = 16'b0000000000000000;
	sram_mem[67260] = 16'b0000000000000000;
	sram_mem[67261] = 16'b0000000000000000;
	sram_mem[67262] = 16'b0000000000000000;
	sram_mem[67263] = 16'b0000000000000000;
	sram_mem[67264] = 16'b0000000000000000;
	sram_mem[67265] = 16'b0000000000000000;
	sram_mem[67266] = 16'b0000000000000000;
	sram_mem[67267] = 16'b0000000000000000;
	sram_mem[67268] = 16'b0000000000000000;
	sram_mem[67269] = 16'b0000000000000000;
	sram_mem[67270] = 16'b0000000000000000;
	sram_mem[67271] = 16'b0000000000000000;
	sram_mem[67272] = 16'b0000000000000000;
	sram_mem[67273] = 16'b0000000000000000;
	sram_mem[67274] = 16'b0000000000000000;
	sram_mem[67275] = 16'b0000000000000000;
	sram_mem[67276] = 16'b0000000000000000;
	sram_mem[67277] = 16'b0000000000000000;
	sram_mem[67278] = 16'b0000000000000000;
	sram_mem[67279] = 16'b0000000000000000;
	sram_mem[67280] = 16'b0000000000000000;
	sram_mem[67281] = 16'b0000000000000000;
	sram_mem[67282] = 16'b0000000000000000;
	sram_mem[67283] = 16'b0000000000000000;
	sram_mem[67284] = 16'b0000000000000000;
	sram_mem[67285] = 16'b0000000000000000;
	sram_mem[67286] = 16'b0000000000000000;
	sram_mem[67287] = 16'b0000000000000000;
	sram_mem[67288] = 16'b0000000000000000;
	sram_mem[67289] = 16'b0000000000000000;
	sram_mem[67290] = 16'b0000000000000000;
	sram_mem[67291] = 16'b0000000000000000;
	sram_mem[67292] = 16'b0000000000000000;
	sram_mem[67293] = 16'b0000000000000000;
	sram_mem[67294] = 16'b0000000000000000;
	sram_mem[67295] = 16'b0000000000000000;
	sram_mem[67296] = 16'b0000000000000000;
	sram_mem[67297] = 16'b0000000000000000;
	sram_mem[67298] = 16'b0000000000000000;
	sram_mem[67299] = 16'b0000000000000000;
	sram_mem[67300] = 16'b0000000000000000;
	sram_mem[67301] = 16'b0000000000000000;
	sram_mem[67302] = 16'b0000000000000000;
	sram_mem[67303] = 16'b0000000000000000;
	sram_mem[67304] = 16'b0000000000000000;
	sram_mem[67305] = 16'b0000000000000000;
	sram_mem[67306] = 16'b0000000000000000;
	sram_mem[67307] = 16'b0000000000000000;
	sram_mem[67308] = 16'b0000000000000000;
	sram_mem[67309] = 16'b0000000000000000;
	sram_mem[67310] = 16'b0000000000000000;
	sram_mem[67311] = 16'b0000000000000000;
	sram_mem[67312] = 16'b0000000000000000;
	sram_mem[67313] = 16'b0000000000000000;
	sram_mem[67314] = 16'b0000000000000000;
	sram_mem[67315] = 16'b0000000000000000;
	sram_mem[67316] = 16'b0000000000000000;
	sram_mem[67317] = 16'b0000000000000000;
	sram_mem[67318] = 16'b0000000000000000;
	sram_mem[67319] = 16'b0000000000000000;
	sram_mem[67320] = 16'b0000000000000000;
	sram_mem[67321] = 16'b0000000000000000;
	sram_mem[67322] = 16'b0000000000000000;
	sram_mem[67323] = 16'b0000000000000000;
	sram_mem[67324] = 16'b0000000000000000;
	sram_mem[67325] = 16'b0000000000000000;
	sram_mem[67326] = 16'b0000000000000000;
	sram_mem[67327] = 16'b0000000000000000;
	sram_mem[67328] = 16'b0000000000000000;
	sram_mem[67329] = 16'b0000000000000000;
	sram_mem[67330] = 16'b0000000000000000;
	sram_mem[67331] = 16'b0000000000000000;
	sram_mem[67332] = 16'b0000000000000000;
	sram_mem[67333] = 16'b0000000000000000;
	sram_mem[67334] = 16'b0000000000000000;
	sram_mem[67335] = 16'b0000000000000000;
	sram_mem[67336] = 16'b0000000000000000;
	sram_mem[67337] = 16'b0000000000000000;
	sram_mem[67338] = 16'b0000000000000000;
	sram_mem[67339] = 16'b0000000000000000;
	sram_mem[67340] = 16'b0000000000000000;
	sram_mem[67341] = 16'b0000000000000000;
	sram_mem[67342] = 16'b0000000000000000;
	sram_mem[67343] = 16'b0000000000000000;
	sram_mem[67344] = 16'b0000000000000000;
	sram_mem[67345] = 16'b0000000000000000;
	sram_mem[67346] = 16'b0000000000000000;
	sram_mem[67347] = 16'b0000000000000000;
	sram_mem[67348] = 16'b0000000000000000;
	sram_mem[67349] = 16'b0000000000000000;
	sram_mem[67350] = 16'b0000000000000000;
	sram_mem[67351] = 16'b0000000000000000;
	sram_mem[67352] = 16'b0000000000000000;
	sram_mem[67353] = 16'b0000000000000000;
	sram_mem[67354] = 16'b0000000000000000;
	sram_mem[67355] = 16'b0000000000000000;
	sram_mem[67356] = 16'b0000000000000000;
	sram_mem[67357] = 16'b0000000000000000;
	sram_mem[67358] = 16'b0000000000000000;
	sram_mem[67359] = 16'b0000000000000000;
	sram_mem[67360] = 16'b0000000000000000;
	sram_mem[67361] = 16'b0000000000000000;
	sram_mem[67362] = 16'b0000000000000000;
	sram_mem[67363] = 16'b0000000000000000;
	sram_mem[67364] = 16'b0000000000000000;
	sram_mem[67365] = 16'b0000000000000000;
	sram_mem[67366] = 16'b0000000000000000;
	sram_mem[67367] = 16'b0000000000000000;
	sram_mem[67368] = 16'b0000000000000000;
	sram_mem[67369] = 16'b0000000000000000;
	sram_mem[67370] = 16'b0000000000000000;
	sram_mem[67371] = 16'b0000000000000000;
	sram_mem[67372] = 16'b0000000000000000;
	sram_mem[67373] = 16'b0000000000000000;
	sram_mem[67374] = 16'b0000000000000000;
	sram_mem[67375] = 16'b0000000000000000;
	sram_mem[67376] = 16'b0000000000000000;
	sram_mem[67377] = 16'b0000000000000000;
	sram_mem[67378] = 16'b0000000000000000;
	sram_mem[67379] = 16'b0000000000000000;
	sram_mem[67380] = 16'b0000000000000000;
	sram_mem[67381] = 16'b0000000000000000;
	sram_mem[67382] = 16'b0000000000000000;
	sram_mem[67383] = 16'b0000000000000000;
	sram_mem[67384] = 16'b0000000000000000;
	sram_mem[67385] = 16'b0000000000000000;
	sram_mem[67386] = 16'b0000000000000000;
	sram_mem[67387] = 16'b0000000000000000;
	sram_mem[67388] = 16'b0000000000000000;
	sram_mem[67389] = 16'b0000000000000000;
	sram_mem[67390] = 16'b0000000000000000;
	sram_mem[67391] = 16'b0000000000000000;
	sram_mem[67392] = 16'b0000000000000000;
	sram_mem[67393] = 16'b0000000000000000;
	sram_mem[67394] = 16'b0000000000000000;
	sram_mem[67395] = 16'b0000000000000000;
	sram_mem[67396] = 16'b0000000000000000;
	sram_mem[67397] = 16'b0000000000000000;
	sram_mem[67398] = 16'b0000000000000000;
	sram_mem[67399] = 16'b0000000000000000;
	sram_mem[67400] = 16'b0000000000000000;
	sram_mem[67401] = 16'b0000000000000000;
	sram_mem[67402] = 16'b0000000000000000;
	sram_mem[67403] = 16'b0000000000000000;
	sram_mem[67404] = 16'b0000000000000000;
	sram_mem[67405] = 16'b0000000000000000;
	sram_mem[67406] = 16'b0000000000000000;
	sram_mem[67407] = 16'b0000000000000000;
	sram_mem[67408] = 16'b0000000000000000;
	sram_mem[67409] = 16'b0000000000000000;
	sram_mem[67410] = 16'b0000000000000000;
	sram_mem[67411] = 16'b0000000000000000;
	sram_mem[67412] = 16'b0000000000000000;
	sram_mem[67413] = 16'b0000000000000000;
	sram_mem[67414] = 16'b0000000000000000;
	sram_mem[67415] = 16'b0000000000000000;
	sram_mem[67416] = 16'b0000000000000000;
	sram_mem[67417] = 16'b0000000000000000;
	sram_mem[67418] = 16'b0000000000000000;
	sram_mem[67419] = 16'b0000000000000000;
	sram_mem[67420] = 16'b0000000000000000;
	sram_mem[67421] = 16'b0000000000000000;
	sram_mem[67422] = 16'b0000000000000000;
	sram_mem[67423] = 16'b0000000000000000;
	sram_mem[67424] = 16'b0000000000000000;
	sram_mem[67425] = 16'b0000000000000000;
	sram_mem[67426] = 16'b0000000000000000;
	sram_mem[67427] = 16'b0000000000000000;
	sram_mem[67428] = 16'b0000000000000000;
	sram_mem[67429] = 16'b0000000000000000;
	sram_mem[67430] = 16'b0000000000000000;
	sram_mem[67431] = 16'b0000000000000000;
	sram_mem[67432] = 16'b0000000000000000;
	sram_mem[67433] = 16'b0000000000000000;
	sram_mem[67434] = 16'b0000000000000000;
	sram_mem[67435] = 16'b0000000000000000;
	sram_mem[67436] = 16'b0000000000000000;
	sram_mem[67437] = 16'b0000000000000000;
	sram_mem[67438] = 16'b0000000000000000;
	sram_mem[67439] = 16'b0000000000000000;
	sram_mem[67440] = 16'b0000000000000000;
	sram_mem[67441] = 16'b0000000000000000;
	sram_mem[67442] = 16'b0000000000000000;
	sram_mem[67443] = 16'b0000000000000000;
	sram_mem[67444] = 16'b0000000000000000;
	sram_mem[67445] = 16'b0000000000000000;
	sram_mem[67446] = 16'b0000000000000000;
	sram_mem[67447] = 16'b0000000000000000;
	sram_mem[67448] = 16'b0000000000000000;
	sram_mem[67449] = 16'b0000000000000000;
	sram_mem[67450] = 16'b0000000000000000;
	sram_mem[67451] = 16'b0000000000000000;
	sram_mem[67452] = 16'b0000000000000000;
	sram_mem[67453] = 16'b0000000000000000;
	sram_mem[67454] = 16'b0000000000000000;
	sram_mem[67455] = 16'b0000000000000000;
	sram_mem[67456] = 16'b0000000000000000;
	sram_mem[67457] = 16'b0000000000000000;
	sram_mem[67458] = 16'b0000000000000000;
	sram_mem[67459] = 16'b0000000000000000;
	sram_mem[67460] = 16'b0000000000000000;
	sram_mem[67461] = 16'b0000000000000000;
	sram_mem[67462] = 16'b0000000000000000;
	sram_mem[67463] = 16'b0000000000000000;
	sram_mem[67464] = 16'b0000000000000000;
	sram_mem[67465] = 16'b0000000000000000;
	sram_mem[67466] = 16'b0000000000000000;
	sram_mem[67467] = 16'b0000000000000000;
	sram_mem[67468] = 16'b0000000000000000;
	sram_mem[67469] = 16'b0000000000000000;
	sram_mem[67470] = 16'b0000000000000000;
	sram_mem[67471] = 16'b0000000000000000;
	sram_mem[67472] = 16'b0000000000000000;
	sram_mem[67473] = 16'b0000000000000000;
	sram_mem[67474] = 16'b0000000000000000;
	sram_mem[67475] = 16'b0000000000000000;
	sram_mem[67476] = 16'b0000000000000000;
	sram_mem[67477] = 16'b0000000000000000;
	sram_mem[67478] = 16'b0000000000000000;
	sram_mem[67479] = 16'b0000000000000000;
	sram_mem[67480] = 16'b0000000000000000;
	sram_mem[67481] = 16'b0000000000000000;
	sram_mem[67482] = 16'b0000000000000000;
	sram_mem[67483] = 16'b0000000000000000;
	sram_mem[67484] = 16'b0000000000000000;
	sram_mem[67485] = 16'b0000000000000000;
	sram_mem[67486] = 16'b0000000000000000;
	sram_mem[67487] = 16'b0000000000000000;
	sram_mem[67488] = 16'b0000000000000000;
	sram_mem[67489] = 16'b0000000000000000;
	sram_mem[67490] = 16'b0000000000000000;
	sram_mem[67491] = 16'b0000000000000000;
	sram_mem[67492] = 16'b0000000000000000;
	sram_mem[67493] = 16'b0000000000000000;
	sram_mem[67494] = 16'b0000000000000000;
	sram_mem[67495] = 16'b0000000000000000;
	sram_mem[67496] = 16'b0000000000000000;
	sram_mem[67497] = 16'b0000000000000000;
	sram_mem[67498] = 16'b0000000000000000;
	sram_mem[67499] = 16'b0000000000000000;
	sram_mem[67500] = 16'b0000000000000000;
	sram_mem[67501] = 16'b0000000000000000;
	sram_mem[67502] = 16'b0000000000000000;
	sram_mem[67503] = 16'b0000000000000000;
	sram_mem[67504] = 16'b0000000000000000;
	sram_mem[67505] = 16'b0000000000000000;
	sram_mem[67506] = 16'b0000000000000000;
	sram_mem[67507] = 16'b0000000000000000;
	sram_mem[67508] = 16'b0000000000000000;
	sram_mem[67509] = 16'b0000000000000000;
	sram_mem[67510] = 16'b0000000000000000;
	sram_mem[67511] = 16'b0000000000000000;
	sram_mem[67512] = 16'b0000000000000000;
	sram_mem[67513] = 16'b0000000000000000;
	sram_mem[67514] = 16'b0000000000000000;
	sram_mem[67515] = 16'b0000000000000000;
	sram_mem[67516] = 16'b0000000000000000;
	sram_mem[67517] = 16'b0000000000000000;
	sram_mem[67518] = 16'b0000000000000000;
	sram_mem[67519] = 16'b0000000000000000;
	sram_mem[67520] = 16'b0000000000000000;
	sram_mem[67521] = 16'b0000000000000000;
	sram_mem[67522] = 16'b0000000000000000;
	sram_mem[67523] = 16'b0000000000000000;
	sram_mem[67524] = 16'b0000000000000000;
	sram_mem[67525] = 16'b0000000000000000;
	sram_mem[67526] = 16'b0000000000000000;
	sram_mem[67527] = 16'b0000000000000000;
	sram_mem[67528] = 16'b0000000000000000;
	sram_mem[67529] = 16'b0000000000000000;
	sram_mem[67530] = 16'b0000000000000000;
	sram_mem[67531] = 16'b0000000000000000;
	sram_mem[67532] = 16'b0000000000000000;
	sram_mem[67533] = 16'b0000000000000000;
	sram_mem[67534] = 16'b0000000000000000;
	sram_mem[67535] = 16'b0000000000000000;
	sram_mem[67536] = 16'b0000000000000000;
	sram_mem[67537] = 16'b0000000000000000;
	sram_mem[67538] = 16'b0000000000000000;
	sram_mem[67539] = 16'b0000000000000000;
	sram_mem[67540] = 16'b0000000000000000;
	sram_mem[67541] = 16'b0000000000000000;
	sram_mem[67542] = 16'b0000000000000000;
	sram_mem[67543] = 16'b0000000000000000;
	sram_mem[67544] = 16'b0000000000000000;
	sram_mem[67545] = 16'b0000000000000000;
	sram_mem[67546] = 16'b0000000000000000;
	sram_mem[67547] = 16'b0000000000000000;
	sram_mem[67548] = 16'b0000000000000000;
	sram_mem[67549] = 16'b0000000000000000;
	sram_mem[67550] = 16'b0000000000000000;
	sram_mem[67551] = 16'b0000000000000000;
	sram_mem[67552] = 16'b0000000000000000;
	sram_mem[67553] = 16'b0000000000000000;
	sram_mem[67554] = 16'b0000000000000000;
	sram_mem[67555] = 16'b0000000000000000;
	sram_mem[67556] = 16'b0000000000000000;
	sram_mem[67557] = 16'b0000000000000000;
	sram_mem[67558] = 16'b0000000000000000;
	sram_mem[67559] = 16'b0000000000000000;
	sram_mem[67560] = 16'b0000000000000000;
	sram_mem[67561] = 16'b0000000000000000;
	sram_mem[67562] = 16'b0000000000000000;
	sram_mem[67563] = 16'b0000000000000000;
	sram_mem[67564] = 16'b0000000000000000;
	sram_mem[67565] = 16'b0000000000000000;
	sram_mem[67566] = 16'b0000000000000000;
	sram_mem[67567] = 16'b0000000000000000;
	sram_mem[67568] = 16'b0000000000000000;
	sram_mem[67569] = 16'b0000000000000000;
	sram_mem[67570] = 16'b0000000000000000;
	sram_mem[67571] = 16'b0000000000000000;
	sram_mem[67572] = 16'b0000000000000000;
	sram_mem[67573] = 16'b0000000000000000;
	sram_mem[67574] = 16'b0000000000000000;
	sram_mem[67575] = 16'b0000000000000000;
	sram_mem[67576] = 16'b0000000000000000;
	sram_mem[67577] = 16'b0000000000000000;
	sram_mem[67578] = 16'b0000000000000000;
	sram_mem[67579] = 16'b0000000000000000;
	sram_mem[67580] = 16'b0000000000000000;
	sram_mem[67581] = 16'b0000000000000000;
	sram_mem[67582] = 16'b0000000000000000;
	sram_mem[67583] = 16'b0000000000000000;
	sram_mem[67584] = 16'b0000000000000000;
	sram_mem[67585] = 16'b0000000000000000;
	sram_mem[67586] = 16'b0000000000000000;
	sram_mem[67587] = 16'b0000000000000000;
	sram_mem[67588] = 16'b0000000000000000;
	sram_mem[67589] = 16'b0000000000000000;
	sram_mem[67590] = 16'b0000000000000000;
	sram_mem[67591] = 16'b0000000000000000;
	sram_mem[67592] = 16'b0000000000000000;
	sram_mem[67593] = 16'b0000000000000000;
	sram_mem[67594] = 16'b0000000000000000;
	sram_mem[67595] = 16'b0000000000000000;
	sram_mem[67596] = 16'b0000000000000000;
	sram_mem[67597] = 16'b0000000000000000;
	sram_mem[67598] = 16'b0000000000000000;
	sram_mem[67599] = 16'b0000000000000000;
	sram_mem[67600] = 16'b0000000000000000;
	sram_mem[67601] = 16'b0000000000000000;
	sram_mem[67602] = 16'b0000000000000000;
	sram_mem[67603] = 16'b0000000000000000;
	sram_mem[67604] = 16'b0000000000000000;
	sram_mem[67605] = 16'b0000000000000000;
	sram_mem[67606] = 16'b0000000000000000;
	sram_mem[67607] = 16'b0000000000000000;
	sram_mem[67608] = 16'b0000000000000000;
	sram_mem[67609] = 16'b0000000000000000;
	sram_mem[67610] = 16'b0000000000000000;
	sram_mem[67611] = 16'b0000000000000000;
	sram_mem[67612] = 16'b0000000000000000;
	sram_mem[67613] = 16'b0000000000000000;
	sram_mem[67614] = 16'b0000000000000000;
	sram_mem[67615] = 16'b0000000000000000;
	sram_mem[67616] = 16'b0000000000000000;
	sram_mem[67617] = 16'b0000000000000000;
	sram_mem[67618] = 16'b0000000000000000;
	sram_mem[67619] = 16'b0000000000000000;
	sram_mem[67620] = 16'b0000000000000000;
	sram_mem[67621] = 16'b0000000000000000;
	sram_mem[67622] = 16'b0000000000000000;
	sram_mem[67623] = 16'b0000000000000000;
	sram_mem[67624] = 16'b0000000000000000;
	sram_mem[67625] = 16'b0000000000000000;
	sram_mem[67626] = 16'b0000000000000000;
	sram_mem[67627] = 16'b0000000000000000;
	sram_mem[67628] = 16'b0000000000000000;
	sram_mem[67629] = 16'b0000000000000000;
	sram_mem[67630] = 16'b0000000000000000;
	sram_mem[67631] = 16'b0000000000000000;
	sram_mem[67632] = 16'b0000000000000000;
	sram_mem[67633] = 16'b0000000000000000;
	sram_mem[67634] = 16'b0000000000000000;
	sram_mem[67635] = 16'b0000000000000000;
	sram_mem[67636] = 16'b0000000000000000;
	sram_mem[67637] = 16'b0000000000000000;
	sram_mem[67638] = 16'b0000000000000000;
	sram_mem[67639] = 16'b0000000000000000;
	sram_mem[67640] = 16'b0000000000000000;
	sram_mem[67641] = 16'b0000000000000000;
	sram_mem[67642] = 16'b0000000000000000;
	sram_mem[67643] = 16'b0000000000000000;
	sram_mem[67644] = 16'b0000000000000000;
	sram_mem[67645] = 16'b0000000000000000;
	sram_mem[67646] = 16'b0000000000000000;
	sram_mem[67647] = 16'b0000000000000000;
	sram_mem[67648] = 16'b0000000000000000;
	sram_mem[67649] = 16'b0000000000000000;
	sram_mem[67650] = 16'b0000000000000000;
	sram_mem[67651] = 16'b0000000000000000;
	sram_mem[67652] = 16'b0000000000000000;
	sram_mem[67653] = 16'b0000000000000000;
	sram_mem[67654] = 16'b0000000000000000;
	sram_mem[67655] = 16'b0000000000000000;
	sram_mem[67656] = 16'b0000000000000000;
	sram_mem[67657] = 16'b0000000000000000;
	sram_mem[67658] = 16'b0000000000000000;
	sram_mem[67659] = 16'b0000000000000000;
	sram_mem[67660] = 16'b0000000000000000;
	sram_mem[67661] = 16'b0000000000000000;
	sram_mem[67662] = 16'b0000000000000000;
	sram_mem[67663] = 16'b0000000000000000;
	sram_mem[67664] = 16'b0000000000000000;
	sram_mem[67665] = 16'b0000000000000000;
	sram_mem[67666] = 16'b0000000000000000;
	sram_mem[67667] = 16'b0000000000000000;
	sram_mem[67668] = 16'b0000000000000000;
	sram_mem[67669] = 16'b0000000000000000;
	sram_mem[67670] = 16'b0000000000000000;
	sram_mem[67671] = 16'b0000000000000000;
	sram_mem[67672] = 16'b0000000000000000;
	sram_mem[67673] = 16'b0000000000000000;
	sram_mem[67674] = 16'b0000000000000000;
	sram_mem[67675] = 16'b0000000000000000;
	sram_mem[67676] = 16'b0000000000000000;
	sram_mem[67677] = 16'b0000000000000000;
	sram_mem[67678] = 16'b0000000000000000;
	sram_mem[67679] = 16'b0000000000000000;
	sram_mem[67680] = 16'b0000000000000000;
	sram_mem[67681] = 16'b0000000000000000;
	sram_mem[67682] = 16'b0000000000000000;
	sram_mem[67683] = 16'b0000000000000000;
	sram_mem[67684] = 16'b0000000000000000;
	sram_mem[67685] = 16'b0000000000000000;
	sram_mem[67686] = 16'b0000000000000000;
	sram_mem[67687] = 16'b0000000000000000;
	sram_mem[67688] = 16'b0000000000000000;
	sram_mem[67689] = 16'b0000000000000000;
	sram_mem[67690] = 16'b0000000000000000;
	sram_mem[67691] = 16'b0000000000000000;
	sram_mem[67692] = 16'b0000000000000000;
	sram_mem[67693] = 16'b0000000000000000;
	sram_mem[67694] = 16'b0000000000000000;
	sram_mem[67695] = 16'b0000000000000000;
	sram_mem[67696] = 16'b0000000000000000;
	sram_mem[67697] = 16'b0000000000000000;
	sram_mem[67698] = 16'b0000000000000000;
	sram_mem[67699] = 16'b0000000000000000;
	sram_mem[67700] = 16'b0000000000000000;
	sram_mem[67701] = 16'b0000000000000000;
	sram_mem[67702] = 16'b0000000000000000;
	sram_mem[67703] = 16'b0000000000000000;
	sram_mem[67704] = 16'b0000000000000000;
	sram_mem[67705] = 16'b0000000000000000;
	sram_mem[67706] = 16'b0000000000000000;
	sram_mem[67707] = 16'b0000000000000000;
	sram_mem[67708] = 16'b0000000000000000;
	sram_mem[67709] = 16'b0000000000000000;
	sram_mem[67710] = 16'b0000000000000000;
	sram_mem[67711] = 16'b0000000000000000;
	sram_mem[67712] = 16'b0000000000000000;
	sram_mem[67713] = 16'b0000000000000000;
	sram_mem[67714] = 16'b0000000000000000;
	sram_mem[67715] = 16'b0000000000000000;
	sram_mem[67716] = 16'b0000000000000000;
	sram_mem[67717] = 16'b0000000000000000;
	sram_mem[67718] = 16'b0000000000000000;
	sram_mem[67719] = 16'b0000000000000000;
	sram_mem[67720] = 16'b0000000000000000;
	sram_mem[67721] = 16'b0000000000000000;
	sram_mem[67722] = 16'b0000000000000000;
	sram_mem[67723] = 16'b0000000000000000;
	sram_mem[67724] = 16'b0000000000000000;
	sram_mem[67725] = 16'b0000000000000000;
	sram_mem[67726] = 16'b0000000000000000;
	sram_mem[67727] = 16'b0000000000000000;
	sram_mem[67728] = 16'b0000000000000000;
	sram_mem[67729] = 16'b0000000000000000;
	sram_mem[67730] = 16'b0000000000000000;
	sram_mem[67731] = 16'b0000000000000000;
	sram_mem[67732] = 16'b0000000000000000;
	sram_mem[67733] = 16'b0000000000000000;
	sram_mem[67734] = 16'b0000000000000000;
	sram_mem[67735] = 16'b0000000000000000;
	sram_mem[67736] = 16'b0000000000000000;
	sram_mem[67737] = 16'b0000000000000000;
	sram_mem[67738] = 16'b0000000000000000;
	sram_mem[67739] = 16'b0000000000000000;
	sram_mem[67740] = 16'b0000000000000000;
	sram_mem[67741] = 16'b0000000000000000;
	sram_mem[67742] = 16'b0000000000000000;
	sram_mem[67743] = 16'b0000000000000000;
	sram_mem[67744] = 16'b0000000000000000;
	sram_mem[67745] = 16'b0000000000000000;
	sram_mem[67746] = 16'b0000000000000000;
	sram_mem[67747] = 16'b0000000000000000;
	sram_mem[67748] = 16'b0000000000000000;
	sram_mem[67749] = 16'b0000000000000000;
	sram_mem[67750] = 16'b0000000000000000;
	sram_mem[67751] = 16'b0000000000000000;
	sram_mem[67752] = 16'b0000000000000000;
	sram_mem[67753] = 16'b0000000000000000;
	sram_mem[67754] = 16'b0000000000000000;
	sram_mem[67755] = 16'b0000000000000000;
	sram_mem[67756] = 16'b0000000000000000;
	sram_mem[67757] = 16'b0000000000000000;
	sram_mem[67758] = 16'b0000000000000000;
	sram_mem[67759] = 16'b0000000000000000;
	sram_mem[67760] = 16'b0000000000000000;
	sram_mem[67761] = 16'b0000000000000000;
	sram_mem[67762] = 16'b0000000000000000;
	sram_mem[67763] = 16'b0000000000000000;
	sram_mem[67764] = 16'b0000000000000000;
	sram_mem[67765] = 16'b0000000000000000;
	sram_mem[67766] = 16'b0000000000000000;
	sram_mem[67767] = 16'b0000000000000000;
	sram_mem[67768] = 16'b0000000000000000;
	sram_mem[67769] = 16'b0000000000000000;
	sram_mem[67770] = 16'b0000000000000000;
	sram_mem[67771] = 16'b0000000000000000;
	sram_mem[67772] = 16'b0000000000000000;
	sram_mem[67773] = 16'b0000000000000000;
	sram_mem[67774] = 16'b0000000000000000;
	sram_mem[67775] = 16'b0000000000000000;
	sram_mem[67776] = 16'b0000000000000000;
	sram_mem[67777] = 16'b0000000000000000;
	sram_mem[67778] = 16'b0000000000000000;
	sram_mem[67779] = 16'b0000000000000000;
	sram_mem[67780] = 16'b0000000000000000;
	sram_mem[67781] = 16'b0000000000000000;
	sram_mem[67782] = 16'b0000000000000000;
	sram_mem[67783] = 16'b0000000000000000;
	sram_mem[67784] = 16'b0000000000000000;
	sram_mem[67785] = 16'b0000000000000000;
	sram_mem[67786] = 16'b0000000000000000;
	sram_mem[67787] = 16'b0000000000000000;
	sram_mem[67788] = 16'b0000000000000000;
	sram_mem[67789] = 16'b0000000000000000;
	sram_mem[67790] = 16'b0000000000000000;
	sram_mem[67791] = 16'b0000000000000000;
	sram_mem[67792] = 16'b0000000000000000;
	sram_mem[67793] = 16'b0000000000000000;
	sram_mem[67794] = 16'b0000000000000000;
	sram_mem[67795] = 16'b0000000000000000;
	sram_mem[67796] = 16'b0000000000000000;
	sram_mem[67797] = 16'b0000000000000000;
	sram_mem[67798] = 16'b0000000000000000;
	sram_mem[67799] = 16'b0000000000000000;
	sram_mem[67800] = 16'b0000000000000000;
	sram_mem[67801] = 16'b0000000000000000;
	sram_mem[67802] = 16'b0000000000000000;
	sram_mem[67803] = 16'b0000000000000000;
	sram_mem[67804] = 16'b0000000000000000;
	sram_mem[67805] = 16'b0000000000000000;
	sram_mem[67806] = 16'b0000000000000000;
	sram_mem[67807] = 16'b0000000000000000;
	sram_mem[67808] = 16'b0000000000000000;
	sram_mem[67809] = 16'b0000000000000000;
	sram_mem[67810] = 16'b0000000000000000;
	sram_mem[67811] = 16'b0000000000000000;
	sram_mem[67812] = 16'b0000000000000000;
	sram_mem[67813] = 16'b0000000000000000;
	sram_mem[67814] = 16'b0000000000000000;
	sram_mem[67815] = 16'b0000000000000000;
	sram_mem[67816] = 16'b0000000000000000;
	sram_mem[67817] = 16'b0000000000000000;
	sram_mem[67818] = 16'b0000000000000000;
	sram_mem[67819] = 16'b0000000000000000;
	sram_mem[67820] = 16'b0000000000000000;
	sram_mem[67821] = 16'b0000000000000000;
	sram_mem[67822] = 16'b0000000000000000;
	sram_mem[67823] = 16'b0000000000000000;
	sram_mem[67824] = 16'b0000000000000000;
	sram_mem[67825] = 16'b0000000000000000;
	sram_mem[67826] = 16'b0000000000000000;
	sram_mem[67827] = 16'b0000000000000000;
	sram_mem[67828] = 16'b0000000000000000;
	sram_mem[67829] = 16'b0000000000000000;
	sram_mem[67830] = 16'b0000000000000000;
	sram_mem[67831] = 16'b0000000000000000;
	sram_mem[67832] = 16'b0000000000000000;
	sram_mem[67833] = 16'b0000000000000000;
	sram_mem[67834] = 16'b0000000000000000;
	sram_mem[67835] = 16'b0000000000000000;
	sram_mem[67836] = 16'b0000000000000000;
	sram_mem[67837] = 16'b0000000000000000;
	sram_mem[67838] = 16'b0000000000000000;
	sram_mem[67839] = 16'b0000000000000000;
	sram_mem[67840] = 16'b0000000000000000;
	sram_mem[67841] = 16'b0000000000000000;
	sram_mem[67842] = 16'b0000000000000000;
	sram_mem[67843] = 16'b0000000000000000;
	sram_mem[67844] = 16'b0000000000000000;
	sram_mem[67845] = 16'b0000000000000000;
	sram_mem[67846] = 16'b0000000000000000;
	sram_mem[67847] = 16'b0000000000000000;
	sram_mem[67848] = 16'b0000000000000000;
	sram_mem[67849] = 16'b0000000000000000;
	sram_mem[67850] = 16'b0000000000000000;
	sram_mem[67851] = 16'b0000000000000000;
	sram_mem[67852] = 16'b0000000000000000;
	sram_mem[67853] = 16'b0000000000000000;
	sram_mem[67854] = 16'b0000000000000000;
	sram_mem[67855] = 16'b0000000000000000;
	sram_mem[67856] = 16'b0000000000000000;
	sram_mem[67857] = 16'b0000000000000000;
	sram_mem[67858] = 16'b0000000000000000;
	sram_mem[67859] = 16'b0000000000000000;
	sram_mem[67860] = 16'b0000000000000000;
	sram_mem[67861] = 16'b0000000000000000;
	sram_mem[67862] = 16'b0000000000000000;
	sram_mem[67863] = 16'b0000000000000000;
	sram_mem[67864] = 16'b0000000000000000;
	sram_mem[67865] = 16'b0000000000000000;
	sram_mem[67866] = 16'b0000000000000000;
	sram_mem[67867] = 16'b0000000000000000;
	sram_mem[67868] = 16'b0000000000000000;
	sram_mem[67869] = 16'b0000000000000000;
	sram_mem[67870] = 16'b0000000000000000;
	sram_mem[67871] = 16'b0000000000000000;
	sram_mem[67872] = 16'b0000000000000000;
	sram_mem[67873] = 16'b0000000000000000;
	sram_mem[67874] = 16'b0000000000000000;
	sram_mem[67875] = 16'b0000000000000000;
	sram_mem[67876] = 16'b0000000000000000;
	sram_mem[67877] = 16'b0000000000000000;
	sram_mem[67878] = 16'b0000000000000000;
	sram_mem[67879] = 16'b0000000000000000;
	sram_mem[67880] = 16'b0000000000000000;
	sram_mem[67881] = 16'b0000000000000000;
	sram_mem[67882] = 16'b0000000000000000;
	sram_mem[67883] = 16'b0000000000000000;
	sram_mem[67884] = 16'b0000000000000000;
	sram_mem[67885] = 16'b0000000000000000;
	sram_mem[67886] = 16'b0000000000000000;
	sram_mem[67887] = 16'b0000000000000000;
	sram_mem[67888] = 16'b0000000000000000;
	sram_mem[67889] = 16'b0000000000000000;
	sram_mem[67890] = 16'b0000000000000000;
	sram_mem[67891] = 16'b0000000000000000;
	sram_mem[67892] = 16'b0000000000000000;
	sram_mem[67893] = 16'b0000000000000000;
	sram_mem[67894] = 16'b0000000000000000;
	sram_mem[67895] = 16'b0000000000000000;
	sram_mem[67896] = 16'b0000000000000000;
	sram_mem[67897] = 16'b0000000000000000;
	sram_mem[67898] = 16'b0000000000000000;
	sram_mem[67899] = 16'b0000000000000000;
	sram_mem[67900] = 16'b0000000000000000;
	sram_mem[67901] = 16'b0000000000000000;
	sram_mem[67902] = 16'b0000000000000000;
	sram_mem[67903] = 16'b0000000000000000;
	sram_mem[67904] = 16'b0000000000000000;
	sram_mem[67905] = 16'b0000000000000000;
	sram_mem[67906] = 16'b0000000000000000;
	sram_mem[67907] = 16'b0000000000000000;
	sram_mem[67908] = 16'b0000000000000000;
	sram_mem[67909] = 16'b0000000000000000;
	sram_mem[67910] = 16'b0000000000000000;
	sram_mem[67911] = 16'b0000000000000000;
	sram_mem[67912] = 16'b0000000000000000;
	sram_mem[67913] = 16'b0000000000000000;
	sram_mem[67914] = 16'b0000000000000000;
	sram_mem[67915] = 16'b0000000000000000;
	sram_mem[67916] = 16'b0000000000000000;
	sram_mem[67917] = 16'b0000000000000000;
	sram_mem[67918] = 16'b0000000000000000;
	sram_mem[67919] = 16'b0000000000000000;
	sram_mem[67920] = 16'b0000000000000000;
	sram_mem[67921] = 16'b0000000000000000;
	sram_mem[67922] = 16'b0000000000000000;
	sram_mem[67923] = 16'b0000000000000000;
	sram_mem[67924] = 16'b0000000000000000;
	sram_mem[67925] = 16'b0000000000000000;
	sram_mem[67926] = 16'b0000000000000000;
	sram_mem[67927] = 16'b0000000000000000;
	sram_mem[67928] = 16'b0000000000000000;
	sram_mem[67929] = 16'b0000000000000000;
	sram_mem[67930] = 16'b0000000000000000;
	sram_mem[67931] = 16'b0000000000000000;
	sram_mem[67932] = 16'b0000000000000000;
	sram_mem[67933] = 16'b0000000000000000;
	sram_mem[67934] = 16'b0000000000000000;
	sram_mem[67935] = 16'b0000000000000000;
	sram_mem[67936] = 16'b0000000000000000;
	sram_mem[67937] = 16'b0000000000000000;
	sram_mem[67938] = 16'b0000000000000000;
	sram_mem[67939] = 16'b0000000000000000;
	sram_mem[67940] = 16'b0000000000000000;
	sram_mem[67941] = 16'b0000000000000000;
	sram_mem[67942] = 16'b0000000000000000;
	sram_mem[67943] = 16'b0000000000000000;
	sram_mem[67944] = 16'b0000000000000000;
	sram_mem[67945] = 16'b0000000000000000;
	sram_mem[67946] = 16'b0000000000000000;
	sram_mem[67947] = 16'b0000000000000000;
	sram_mem[67948] = 16'b0000000000000000;
	sram_mem[67949] = 16'b0000000000000000;
	sram_mem[67950] = 16'b0000000000000000;
	sram_mem[67951] = 16'b0000000000000000;
	sram_mem[67952] = 16'b0000000000000000;
	sram_mem[67953] = 16'b0000000000000000;
	sram_mem[67954] = 16'b0000000000000000;
	sram_mem[67955] = 16'b0000000000000000;
	sram_mem[67956] = 16'b0000000000000000;
	sram_mem[67957] = 16'b0000000000000000;
	sram_mem[67958] = 16'b0000000000000000;
	sram_mem[67959] = 16'b0000000000000000;
	sram_mem[67960] = 16'b0000000000000000;
	sram_mem[67961] = 16'b0000000000000000;
	sram_mem[67962] = 16'b0000000000000000;
	sram_mem[67963] = 16'b0000000000000000;
	sram_mem[67964] = 16'b0000000000000000;
	sram_mem[67965] = 16'b0000000000000000;
	sram_mem[67966] = 16'b0000000000000000;
	sram_mem[67967] = 16'b0000000000000000;
	sram_mem[67968] = 16'b0000000000000000;
	sram_mem[67969] = 16'b0000000000000000;
	sram_mem[67970] = 16'b0000000000000000;
	sram_mem[67971] = 16'b0000000000000000;
	sram_mem[67972] = 16'b0000000000000000;
	sram_mem[67973] = 16'b0000000000000000;
	sram_mem[67974] = 16'b0000000000000000;
	sram_mem[67975] = 16'b0000000000000000;
	sram_mem[67976] = 16'b0000000000000000;
	sram_mem[67977] = 16'b0000000000000000;
	sram_mem[67978] = 16'b0000000000000000;
	sram_mem[67979] = 16'b0000000000000000;
	sram_mem[67980] = 16'b0000000000000000;
	sram_mem[67981] = 16'b0000000000000000;
	sram_mem[67982] = 16'b0000000000000000;
	sram_mem[67983] = 16'b0000000000000000;
	sram_mem[67984] = 16'b0000000000000000;
	sram_mem[67985] = 16'b0000000000000000;
	sram_mem[67986] = 16'b0000000000000000;
	sram_mem[67987] = 16'b0000000000000000;
	sram_mem[67988] = 16'b0000000000000000;
	sram_mem[67989] = 16'b0000000000000000;
	sram_mem[67990] = 16'b0000000000000000;
	sram_mem[67991] = 16'b0000000000000000;
	sram_mem[67992] = 16'b0000000000000000;
	sram_mem[67993] = 16'b0000000000000000;
	sram_mem[67994] = 16'b0000000000000000;
	sram_mem[67995] = 16'b0000000000000000;
	sram_mem[67996] = 16'b0000000000000000;
	sram_mem[67997] = 16'b0000000000000000;
	sram_mem[67998] = 16'b0000000000000000;
	sram_mem[67999] = 16'b0000000000000000;
	sram_mem[68000] = 16'b0000000000000000;
	sram_mem[68001] = 16'b0000000000000000;
	sram_mem[68002] = 16'b0000000000000000;
	sram_mem[68003] = 16'b0000000000000000;
	sram_mem[68004] = 16'b0000000000000000;
	sram_mem[68005] = 16'b0000000000000000;
	sram_mem[68006] = 16'b0000000000000000;
	sram_mem[68007] = 16'b0000000000000000;
	sram_mem[68008] = 16'b0000000000000000;
	sram_mem[68009] = 16'b0000000000000000;
	sram_mem[68010] = 16'b0000000000000000;
	sram_mem[68011] = 16'b0000000000000000;
	sram_mem[68012] = 16'b0000000000000000;
	sram_mem[68013] = 16'b0000000000000000;
	sram_mem[68014] = 16'b0000000000000000;
	sram_mem[68015] = 16'b0000000000000000;
	sram_mem[68016] = 16'b0000000000000000;
	sram_mem[68017] = 16'b0000000000000000;
	sram_mem[68018] = 16'b0000000000000000;
	sram_mem[68019] = 16'b0000000000000000;
	sram_mem[68020] = 16'b0000000000000000;
	sram_mem[68021] = 16'b0000000000000000;
	sram_mem[68022] = 16'b0000000000000000;
	sram_mem[68023] = 16'b0000000000000000;
	sram_mem[68024] = 16'b0000000000000000;
	sram_mem[68025] = 16'b0000000000000000;
	sram_mem[68026] = 16'b0000000000000000;
	sram_mem[68027] = 16'b0000000000000000;
	sram_mem[68028] = 16'b0000000000000000;
	sram_mem[68029] = 16'b0000000000000000;
	sram_mem[68030] = 16'b0000000000000000;
	sram_mem[68031] = 16'b0000000000000000;
	sram_mem[68032] = 16'b0000000000000000;
	sram_mem[68033] = 16'b0000000000000000;
	sram_mem[68034] = 16'b0000000000000000;
	sram_mem[68035] = 16'b0000000000000000;
	sram_mem[68036] = 16'b0000000000000000;
	sram_mem[68037] = 16'b0000000000000000;
	sram_mem[68038] = 16'b0000000000000000;
	sram_mem[68039] = 16'b0000000000000000;
	sram_mem[68040] = 16'b0000000000000000;
	sram_mem[68041] = 16'b0000000000000000;
	sram_mem[68042] = 16'b0000000000000000;
	sram_mem[68043] = 16'b0000000000000000;
	sram_mem[68044] = 16'b0000000000000000;
	sram_mem[68045] = 16'b0000000000000000;
	sram_mem[68046] = 16'b0000000000000000;
	sram_mem[68047] = 16'b0000000000000000;
	sram_mem[68048] = 16'b0000000000000000;
	sram_mem[68049] = 16'b0000000000000000;
	sram_mem[68050] = 16'b0000000000000000;
	sram_mem[68051] = 16'b0000000000000000;
	sram_mem[68052] = 16'b0000000000000000;
	sram_mem[68053] = 16'b0000000000000000;
	sram_mem[68054] = 16'b0000000000000000;
	sram_mem[68055] = 16'b0000000000000000;
	sram_mem[68056] = 16'b0000000000000000;
	sram_mem[68057] = 16'b0000000000000000;
	sram_mem[68058] = 16'b0000000000000000;
	sram_mem[68059] = 16'b0000000000000000;
	sram_mem[68060] = 16'b0000000000000000;
	sram_mem[68061] = 16'b0000000000000000;
	sram_mem[68062] = 16'b0000000000000000;
	sram_mem[68063] = 16'b0000000000000000;
	sram_mem[68064] = 16'b0000000000000000;
	sram_mem[68065] = 16'b0000000000000000;
	sram_mem[68066] = 16'b0000000000000000;
	sram_mem[68067] = 16'b0000000000000000;
	sram_mem[68068] = 16'b0000000000000000;
	sram_mem[68069] = 16'b0000000000000000;
	sram_mem[68070] = 16'b0000000000000000;
	sram_mem[68071] = 16'b0000000000000000;
	sram_mem[68072] = 16'b0000000000000000;
	sram_mem[68073] = 16'b0000000000000000;
	sram_mem[68074] = 16'b0000000000000000;
	sram_mem[68075] = 16'b0000000000000000;
	sram_mem[68076] = 16'b0000000000000000;
	sram_mem[68077] = 16'b0000000000000000;
	sram_mem[68078] = 16'b0000000000000000;
	sram_mem[68079] = 16'b0000000000000000;
	sram_mem[68080] = 16'b0000000000000000;
	sram_mem[68081] = 16'b0000000000000000;
	sram_mem[68082] = 16'b0000000000000000;
	sram_mem[68083] = 16'b0000000000000000;
	sram_mem[68084] = 16'b0000000000000000;
	sram_mem[68085] = 16'b0000000000000000;
	sram_mem[68086] = 16'b0000000000000000;
	sram_mem[68087] = 16'b0000000000000000;
	sram_mem[68088] = 16'b0000000000000000;
	sram_mem[68089] = 16'b0000000000000000;
	sram_mem[68090] = 16'b0000000000000000;
	sram_mem[68091] = 16'b0000000000000000;
	sram_mem[68092] = 16'b0000000000000000;
	sram_mem[68093] = 16'b0000000000000000;
	sram_mem[68094] = 16'b0000000000000000;
	sram_mem[68095] = 16'b0000000000000000;
	sram_mem[68096] = 16'b0000000000000000;
	sram_mem[68097] = 16'b0000000000000000;
	sram_mem[68098] = 16'b0000000000000000;
	sram_mem[68099] = 16'b0000000000000000;
	sram_mem[68100] = 16'b0000000000000000;
	sram_mem[68101] = 16'b0000000000000000;
	sram_mem[68102] = 16'b0000000000000000;
	sram_mem[68103] = 16'b0000000000000000;
	sram_mem[68104] = 16'b0000000000000000;
	sram_mem[68105] = 16'b0000000000000000;
	sram_mem[68106] = 16'b0000000000000000;
	sram_mem[68107] = 16'b0000000000000000;
	sram_mem[68108] = 16'b0000000000000000;
	sram_mem[68109] = 16'b0000000000000000;
	sram_mem[68110] = 16'b0000000000000000;
	sram_mem[68111] = 16'b0000000000000000;
	sram_mem[68112] = 16'b0000000000000000;
	sram_mem[68113] = 16'b0000000000000000;
	sram_mem[68114] = 16'b0000000000000000;
	sram_mem[68115] = 16'b0000000000000000;
	sram_mem[68116] = 16'b0000000000000000;
	sram_mem[68117] = 16'b0000000000000000;
	sram_mem[68118] = 16'b0000000000000000;
	sram_mem[68119] = 16'b0000000000000000;
	sram_mem[68120] = 16'b0000000000000000;
	sram_mem[68121] = 16'b0000000000000000;
	sram_mem[68122] = 16'b0000000000000000;
	sram_mem[68123] = 16'b0000000000000000;
	sram_mem[68124] = 16'b0000000000000000;
	sram_mem[68125] = 16'b0000000000000000;
	sram_mem[68126] = 16'b0000000000000000;
	sram_mem[68127] = 16'b0000000000000000;
	sram_mem[68128] = 16'b0000000000000000;
	sram_mem[68129] = 16'b0000000000000000;
	sram_mem[68130] = 16'b0000000000000000;
	sram_mem[68131] = 16'b0000000000000000;
	sram_mem[68132] = 16'b0000000000000000;
	sram_mem[68133] = 16'b0000000000000000;
	sram_mem[68134] = 16'b0000000000000000;
	sram_mem[68135] = 16'b0000000000000000;
	sram_mem[68136] = 16'b0000000000000000;
	sram_mem[68137] = 16'b0000000000000000;
	sram_mem[68138] = 16'b0000000000000000;
	sram_mem[68139] = 16'b0000000000000000;
	sram_mem[68140] = 16'b0000000000000000;
	sram_mem[68141] = 16'b0000000000000000;
	sram_mem[68142] = 16'b0000000000000000;
	sram_mem[68143] = 16'b0000000000000000;
	sram_mem[68144] = 16'b0000000000000000;
	sram_mem[68145] = 16'b0000000000000000;
	sram_mem[68146] = 16'b0000000000000000;
	sram_mem[68147] = 16'b0000000000000000;
	sram_mem[68148] = 16'b0000000000000000;
	sram_mem[68149] = 16'b0000000000000000;
	sram_mem[68150] = 16'b0000000000000000;
	sram_mem[68151] = 16'b0000000000000000;
	sram_mem[68152] = 16'b0000000000000000;
	sram_mem[68153] = 16'b0000000000000000;
	sram_mem[68154] = 16'b0000000000000000;
	sram_mem[68155] = 16'b0000000000000000;
	sram_mem[68156] = 16'b0000000000000000;
	sram_mem[68157] = 16'b0000000000000000;
	sram_mem[68158] = 16'b0000000000000000;
	sram_mem[68159] = 16'b0000000000000000;
	sram_mem[68160] = 16'b0000000000000000;
	sram_mem[68161] = 16'b0000000000000000;
	sram_mem[68162] = 16'b0000000000000000;
	sram_mem[68163] = 16'b0000000000000000;
	sram_mem[68164] = 16'b0000000000000000;
	sram_mem[68165] = 16'b0000000000000000;
	sram_mem[68166] = 16'b0000000000000000;
	sram_mem[68167] = 16'b0000000000000000;
	sram_mem[68168] = 16'b0000000000000000;
	sram_mem[68169] = 16'b0000000000000000;
	sram_mem[68170] = 16'b0000000000000000;
	sram_mem[68171] = 16'b0000000000000000;
	sram_mem[68172] = 16'b0000000000000000;
	sram_mem[68173] = 16'b0000000000000000;
	sram_mem[68174] = 16'b0000000000000000;
	sram_mem[68175] = 16'b0000000000000000;
	sram_mem[68176] = 16'b0000000000000000;
	sram_mem[68177] = 16'b0000000000000000;
	sram_mem[68178] = 16'b0000000000000000;
	sram_mem[68179] = 16'b0000000000000000;
	sram_mem[68180] = 16'b0000000000000000;
	sram_mem[68181] = 16'b0000000000000000;
	sram_mem[68182] = 16'b0000000000000000;
	sram_mem[68183] = 16'b0000000000000000;
	sram_mem[68184] = 16'b0000000000000000;
	sram_mem[68185] = 16'b0000000000000000;
	sram_mem[68186] = 16'b0000000000000000;
	sram_mem[68187] = 16'b0000000000000000;
	sram_mem[68188] = 16'b0000000000000000;
	sram_mem[68189] = 16'b0000000000000000;
	sram_mem[68190] = 16'b0000000000000000;
	sram_mem[68191] = 16'b0000000000000000;
	sram_mem[68192] = 16'b0000000000000000;
	sram_mem[68193] = 16'b0000000000000000;
	sram_mem[68194] = 16'b0000000000000000;
	sram_mem[68195] = 16'b0000000000000000;
	sram_mem[68196] = 16'b0000000000000000;
	sram_mem[68197] = 16'b0000000000000000;
	sram_mem[68198] = 16'b0000000000000000;
	sram_mem[68199] = 16'b0000000000000000;
	sram_mem[68200] = 16'b0000000000000000;
	sram_mem[68201] = 16'b0000000000000000;
	sram_mem[68202] = 16'b0000000000000000;
	sram_mem[68203] = 16'b0000000000000000;
	sram_mem[68204] = 16'b0000000000000000;
	sram_mem[68205] = 16'b0000000000000000;
	sram_mem[68206] = 16'b0000000000000000;
	sram_mem[68207] = 16'b0000000000000000;
	sram_mem[68208] = 16'b0000000000000000;
	sram_mem[68209] = 16'b0000000000000000;
	sram_mem[68210] = 16'b0000000000000000;
	sram_mem[68211] = 16'b0000000000000000;
	sram_mem[68212] = 16'b0000000000000000;
	sram_mem[68213] = 16'b0000000000000000;
	sram_mem[68214] = 16'b0000000000000000;
	sram_mem[68215] = 16'b0000000000000000;
	sram_mem[68216] = 16'b0000000000000000;
	sram_mem[68217] = 16'b0000000000000000;
	sram_mem[68218] = 16'b0000000000000000;
	sram_mem[68219] = 16'b0000000000000000;
	sram_mem[68220] = 16'b0000000000000000;
	sram_mem[68221] = 16'b0000000000000000;
	sram_mem[68222] = 16'b0000000000000000;
	sram_mem[68223] = 16'b0000000000000000;
	sram_mem[68224] = 16'b0000000000000000;
	sram_mem[68225] = 16'b0000000000000000;
	sram_mem[68226] = 16'b0000000000000000;
	sram_mem[68227] = 16'b0000000000000000;
	sram_mem[68228] = 16'b0000000000000000;
	sram_mem[68229] = 16'b0000000000000000;
	sram_mem[68230] = 16'b0000000000000000;
	sram_mem[68231] = 16'b0000000000000000;
	sram_mem[68232] = 16'b0000000000000000;
	sram_mem[68233] = 16'b0000000000000000;
	sram_mem[68234] = 16'b0000000000000000;
	sram_mem[68235] = 16'b0000000000000000;
	sram_mem[68236] = 16'b0000000000000000;
	sram_mem[68237] = 16'b0000000000000000;
	sram_mem[68238] = 16'b0000000000000000;
	sram_mem[68239] = 16'b0000000000000000;
	sram_mem[68240] = 16'b0000000000000000;
	sram_mem[68241] = 16'b0000000000000000;
	sram_mem[68242] = 16'b0000000000000000;
	sram_mem[68243] = 16'b0000000000000000;
	sram_mem[68244] = 16'b0000000000000000;
	sram_mem[68245] = 16'b0000000000000000;
	sram_mem[68246] = 16'b0000000000000000;
	sram_mem[68247] = 16'b0000000000000000;
	sram_mem[68248] = 16'b0000000000000000;
	sram_mem[68249] = 16'b0000000000000000;
	sram_mem[68250] = 16'b0000000000000000;
	sram_mem[68251] = 16'b0000000000000000;
	sram_mem[68252] = 16'b0000000000000000;
	sram_mem[68253] = 16'b0000000000000000;
	sram_mem[68254] = 16'b0000000000000000;
	sram_mem[68255] = 16'b0000000000000000;
	sram_mem[68256] = 16'b0000000000000000;
	sram_mem[68257] = 16'b0000000000000000;
	sram_mem[68258] = 16'b0000000000000000;
	sram_mem[68259] = 16'b0000000000000000;
	sram_mem[68260] = 16'b0000000000000000;
	sram_mem[68261] = 16'b0000000000000000;
	sram_mem[68262] = 16'b0000000000000000;
	sram_mem[68263] = 16'b0000000000000000;
	sram_mem[68264] = 16'b0000000000000000;
	sram_mem[68265] = 16'b0000000000000000;
	sram_mem[68266] = 16'b0000000000000000;
	sram_mem[68267] = 16'b0000000000000000;
	sram_mem[68268] = 16'b0000000000000000;
	sram_mem[68269] = 16'b0000000000000000;
	sram_mem[68270] = 16'b0000000000000000;
	sram_mem[68271] = 16'b0000000000000000;
	sram_mem[68272] = 16'b0000000000000000;
	sram_mem[68273] = 16'b0000000000000000;
	sram_mem[68274] = 16'b0000000000000000;
	sram_mem[68275] = 16'b0000000000000000;
	sram_mem[68276] = 16'b0000000000000000;
	sram_mem[68277] = 16'b0000000000000000;
	sram_mem[68278] = 16'b0000000000000000;
	sram_mem[68279] = 16'b0000000000000000;
	sram_mem[68280] = 16'b0000000000000000;
	sram_mem[68281] = 16'b0000000000000000;
	sram_mem[68282] = 16'b0000000000000000;
	sram_mem[68283] = 16'b0000000000000000;
	sram_mem[68284] = 16'b0000000000000000;
	sram_mem[68285] = 16'b0000000000000000;
	sram_mem[68286] = 16'b0000000000000000;
	sram_mem[68287] = 16'b0000000000000000;
	sram_mem[68288] = 16'b0000000000000000;
	sram_mem[68289] = 16'b0000000000000000;
	sram_mem[68290] = 16'b0000000000000000;
	sram_mem[68291] = 16'b0000000000000000;
	sram_mem[68292] = 16'b0000000000000000;
	sram_mem[68293] = 16'b0000000000000000;
	sram_mem[68294] = 16'b0000000000000000;
	sram_mem[68295] = 16'b0000000000000000;
	sram_mem[68296] = 16'b0000000000000000;
	sram_mem[68297] = 16'b0000000000000000;
	sram_mem[68298] = 16'b0000000000000000;
	sram_mem[68299] = 16'b0000000000000000;
	sram_mem[68300] = 16'b0000000000000000;
	sram_mem[68301] = 16'b0000000000000000;
	sram_mem[68302] = 16'b0000000000000000;
	sram_mem[68303] = 16'b0000000000000000;
	sram_mem[68304] = 16'b0000000000000000;
	sram_mem[68305] = 16'b0000000000000000;
	sram_mem[68306] = 16'b0000000000000000;
	sram_mem[68307] = 16'b0000000000000000;
	sram_mem[68308] = 16'b0000000000000000;
	sram_mem[68309] = 16'b0000000000000000;
	sram_mem[68310] = 16'b0000000000000000;
	sram_mem[68311] = 16'b0000000000000000;
	sram_mem[68312] = 16'b0000000000000000;
	sram_mem[68313] = 16'b0000000000000000;
	sram_mem[68314] = 16'b0000000000000000;
	sram_mem[68315] = 16'b0000000000000000;
	sram_mem[68316] = 16'b0000000000000000;
	sram_mem[68317] = 16'b0000000000000000;
	sram_mem[68318] = 16'b0000000000000000;
	sram_mem[68319] = 16'b0000000000000000;
	sram_mem[68320] = 16'b0000000000000000;
	sram_mem[68321] = 16'b0000000000000000;
	sram_mem[68322] = 16'b0000000000000000;
	sram_mem[68323] = 16'b0000000000000000;
	sram_mem[68324] = 16'b0000000000000000;
	sram_mem[68325] = 16'b0000000000000000;
	sram_mem[68326] = 16'b0000000000000000;
	sram_mem[68327] = 16'b0000000000000000;
	sram_mem[68328] = 16'b0000000000000000;
	sram_mem[68329] = 16'b0000000000000000;
	sram_mem[68330] = 16'b0000000000000000;
	sram_mem[68331] = 16'b0000000000000000;
	sram_mem[68332] = 16'b0000000000000000;
	sram_mem[68333] = 16'b0000000000000000;
	sram_mem[68334] = 16'b0000000000000000;
	sram_mem[68335] = 16'b0000000000000000;
	sram_mem[68336] = 16'b0000000000000000;
	sram_mem[68337] = 16'b0000000000000000;
	sram_mem[68338] = 16'b0000000000000000;
	sram_mem[68339] = 16'b0000000000000000;
	sram_mem[68340] = 16'b0000000000000000;
	sram_mem[68341] = 16'b0000000000000000;
	sram_mem[68342] = 16'b0000000000000000;
	sram_mem[68343] = 16'b0000000000000000;
	sram_mem[68344] = 16'b0000000000000000;
	sram_mem[68345] = 16'b0000000000000000;
	sram_mem[68346] = 16'b0000000000000000;
	sram_mem[68347] = 16'b0000000000000000;
	sram_mem[68348] = 16'b0000000000000000;
	sram_mem[68349] = 16'b0000000000000000;
	sram_mem[68350] = 16'b0000000000000000;
	sram_mem[68351] = 16'b0000000000000000;
	sram_mem[68352] = 16'b0000000000000000;
	sram_mem[68353] = 16'b0000000000000000;
	sram_mem[68354] = 16'b0000000000000000;
	sram_mem[68355] = 16'b0000000000000000;
	sram_mem[68356] = 16'b0000000000000000;
	sram_mem[68357] = 16'b0000000000000000;
	sram_mem[68358] = 16'b0000000000000000;
	sram_mem[68359] = 16'b0000000000000000;
	sram_mem[68360] = 16'b0000000000000000;
	sram_mem[68361] = 16'b0000000000000000;
	sram_mem[68362] = 16'b0000000000000000;
	sram_mem[68363] = 16'b0000000000000000;
	sram_mem[68364] = 16'b0000000000000000;
	sram_mem[68365] = 16'b0000000000000000;
	sram_mem[68366] = 16'b0000000000000000;
	sram_mem[68367] = 16'b0000000000000000;
	sram_mem[68368] = 16'b0000000000000000;
	sram_mem[68369] = 16'b0000000000000000;
	sram_mem[68370] = 16'b0000000000000000;
	sram_mem[68371] = 16'b0000000000000000;
	sram_mem[68372] = 16'b0000000000000000;
	sram_mem[68373] = 16'b0000000000000000;
	sram_mem[68374] = 16'b0000000000000000;
	sram_mem[68375] = 16'b0000000000000000;
	sram_mem[68376] = 16'b0000000000000000;
	sram_mem[68377] = 16'b0000000000000000;
	sram_mem[68378] = 16'b0000000000000000;
	sram_mem[68379] = 16'b0000000000000000;
	sram_mem[68380] = 16'b0000000000000000;
	sram_mem[68381] = 16'b0000000000000000;
	sram_mem[68382] = 16'b0000000000000000;
	sram_mem[68383] = 16'b0000000000000000;
	sram_mem[68384] = 16'b0000000000000000;
	sram_mem[68385] = 16'b0000000000000000;
	sram_mem[68386] = 16'b0000000000000000;
	sram_mem[68387] = 16'b0000000000000000;
	sram_mem[68388] = 16'b0000000000000000;
	sram_mem[68389] = 16'b0000000000000000;
	sram_mem[68390] = 16'b0000000000000000;
	sram_mem[68391] = 16'b0000000000000000;
	sram_mem[68392] = 16'b0000000000000000;
	sram_mem[68393] = 16'b0000000000000000;
	sram_mem[68394] = 16'b0000000000000000;
	sram_mem[68395] = 16'b0000000000000000;
	sram_mem[68396] = 16'b0000000000000000;
	sram_mem[68397] = 16'b0000000000000000;
	sram_mem[68398] = 16'b0000000000000000;
	sram_mem[68399] = 16'b0000000000000000;
	sram_mem[68400] = 16'b0000000000000000;
	sram_mem[68401] = 16'b0000000000000000;
	sram_mem[68402] = 16'b0000000000000000;
	sram_mem[68403] = 16'b0000000000000000;
	sram_mem[68404] = 16'b0000000000000000;
	sram_mem[68405] = 16'b0000000000000000;
	sram_mem[68406] = 16'b0000000000000000;
	sram_mem[68407] = 16'b0000000000000000;
	sram_mem[68408] = 16'b0000000000000000;
	sram_mem[68409] = 16'b0000000000000000;
	sram_mem[68410] = 16'b0000000000000000;
	sram_mem[68411] = 16'b0000000000000000;
	sram_mem[68412] = 16'b0000000000000000;
	sram_mem[68413] = 16'b0000000000000000;
	sram_mem[68414] = 16'b0000000000000000;
	sram_mem[68415] = 16'b0000000000000000;
	sram_mem[68416] = 16'b0000000000000000;
	sram_mem[68417] = 16'b0000000000000000;
	sram_mem[68418] = 16'b0000000000000000;
	sram_mem[68419] = 16'b0000000000000000;
	sram_mem[68420] = 16'b0000000000000000;
	sram_mem[68421] = 16'b0000000000000000;
	sram_mem[68422] = 16'b0000000000000000;
	sram_mem[68423] = 16'b0000000000000000;
	sram_mem[68424] = 16'b0000000000000000;
	sram_mem[68425] = 16'b0000000000000000;
	sram_mem[68426] = 16'b0000000000000000;
	sram_mem[68427] = 16'b0000000000000000;
	sram_mem[68428] = 16'b0000000000000000;
	sram_mem[68429] = 16'b0000000000000000;
	sram_mem[68430] = 16'b0000000000000000;
	sram_mem[68431] = 16'b0000000000000000;
	sram_mem[68432] = 16'b0000000000000000;
	sram_mem[68433] = 16'b0000000000000000;
	sram_mem[68434] = 16'b0000000000000000;
	sram_mem[68435] = 16'b0000000000000000;
	sram_mem[68436] = 16'b0000000000000000;
	sram_mem[68437] = 16'b0000000000000000;
	sram_mem[68438] = 16'b0000000000000000;
	sram_mem[68439] = 16'b0000000000000000;
	sram_mem[68440] = 16'b0000000000000000;
	sram_mem[68441] = 16'b0000000000000000;
	sram_mem[68442] = 16'b0000000000000000;
	sram_mem[68443] = 16'b0000000000000000;
	sram_mem[68444] = 16'b0000000000000000;
	sram_mem[68445] = 16'b0000000000000000;
	sram_mem[68446] = 16'b0000000000000000;
	sram_mem[68447] = 16'b0000000000000000;
	sram_mem[68448] = 16'b0000000000000000;
	sram_mem[68449] = 16'b0000000000000000;
	sram_mem[68450] = 16'b0000000000000000;
	sram_mem[68451] = 16'b0000000000000000;
	sram_mem[68452] = 16'b0000000000000000;
	sram_mem[68453] = 16'b0000000000000000;
	sram_mem[68454] = 16'b0000000000000000;
	sram_mem[68455] = 16'b0000000000000000;
	sram_mem[68456] = 16'b0000000000000000;
	sram_mem[68457] = 16'b0000000000000000;
	sram_mem[68458] = 16'b0000000000000000;
	sram_mem[68459] = 16'b0000000000000000;
	sram_mem[68460] = 16'b0000000000000000;
	sram_mem[68461] = 16'b0000000000000000;
	sram_mem[68462] = 16'b0000000000000000;
	sram_mem[68463] = 16'b0000000000000000;
	sram_mem[68464] = 16'b0000000000000000;
	sram_mem[68465] = 16'b0000000000000000;
	sram_mem[68466] = 16'b0000000000000000;
	sram_mem[68467] = 16'b0000000000000000;
	sram_mem[68468] = 16'b0000000000000000;
	sram_mem[68469] = 16'b0000000000000000;
	sram_mem[68470] = 16'b0000000000000000;
	sram_mem[68471] = 16'b0000000000000000;
	sram_mem[68472] = 16'b0000000000000000;
	sram_mem[68473] = 16'b0000000000000000;
	sram_mem[68474] = 16'b0000000000000000;
	sram_mem[68475] = 16'b0000000000000000;
	sram_mem[68476] = 16'b0000000000000000;
	sram_mem[68477] = 16'b0000000000000000;
	sram_mem[68478] = 16'b0000000000000000;
	sram_mem[68479] = 16'b0000000000000000;
	sram_mem[68480] = 16'b0000000000000000;
	sram_mem[68481] = 16'b0000000000000000;
	sram_mem[68482] = 16'b0000000000000000;
	sram_mem[68483] = 16'b0000000000000000;
	sram_mem[68484] = 16'b0000000000000000;
	sram_mem[68485] = 16'b0000000000000000;
	sram_mem[68486] = 16'b0000000000000000;
	sram_mem[68487] = 16'b0000000000000000;
	sram_mem[68488] = 16'b0000000000000000;
	sram_mem[68489] = 16'b0000000000000000;
	sram_mem[68490] = 16'b0000000000000000;
	sram_mem[68491] = 16'b0000000000000000;
	sram_mem[68492] = 16'b0000000000000000;
	sram_mem[68493] = 16'b0000000000000000;
	sram_mem[68494] = 16'b0000000000000000;
	sram_mem[68495] = 16'b0000000000000000;
	sram_mem[68496] = 16'b0000000000000000;
	sram_mem[68497] = 16'b0000000000000000;
	sram_mem[68498] = 16'b0000000000000000;
	sram_mem[68499] = 16'b0000000000000000;
	sram_mem[68500] = 16'b0000000000000000;
	sram_mem[68501] = 16'b0000000000000000;
	sram_mem[68502] = 16'b0000000000000000;
	sram_mem[68503] = 16'b0000000000000000;
	sram_mem[68504] = 16'b0000000000000000;
	sram_mem[68505] = 16'b0000000000000000;
	sram_mem[68506] = 16'b0000000000000000;
	sram_mem[68507] = 16'b0000000000000000;
	sram_mem[68508] = 16'b0000000000000000;
	sram_mem[68509] = 16'b0000000000000000;
	sram_mem[68510] = 16'b0000000000000000;
	sram_mem[68511] = 16'b0000000000000000;
	sram_mem[68512] = 16'b0000000000000000;
	sram_mem[68513] = 16'b0000000000000000;
	sram_mem[68514] = 16'b0000000000000000;
	sram_mem[68515] = 16'b0000000000000000;
	sram_mem[68516] = 16'b0000000000000000;
	sram_mem[68517] = 16'b0000000000000000;
	sram_mem[68518] = 16'b0000000000000000;
	sram_mem[68519] = 16'b0000000000000000;
	sram_mem[68520] = 16'b0000000000000000;
	sram_mem[68521] = 16'b0000000000000000;
	sram_mem[68522] = 16'b0000000000000000;
	sram_mem[68523] = 16'b0000000000000000;
	sram_mem[68524] = 16'b0000000000000000;
	sram_mem[68525] = 16'b0000000000000000;
	sram_mem[68526] = 16'b0000000000000000;
	sram_mem[68527] = 16'b0000000000000000;
	sram_mem[68528] = 16'b0000000000000000;
	sram_mem[68529] = 16'b0000000000000000;
	sram_mem[68530] = 16'b0000000000000000;
	sram_mem[68531] = 16'b0000000000000000;
	sram_mem[68532] = 16'b0000000000000000;
	sram_mem[68533] = 16'b0000000000000000;
	sram_mem[68534] = 16'b0000000000000000;
	sram_mem[68535] = 16'b0000000000000000;
	sram_mem[68536] = 16'b0000000000000000;
	sram_mem[68537] = 16'b0000000000000000;
	sram_mem[68538] = 16'b0000000000000000;
	sram_mem[68539] = 16'b0000000000000000;
	sram_mem[68540] = 16'b0000000000000000;
	sram_mem[68541] = 16'b0000000000000000;
	sram_mem[68542] = 16'b0000000000000000;
	sram_mem[68543] = 16'b0000000000000000;
	sram_mem[68544] = 16'b0000000000000000;
	sram_mem[68545] = 16'b0000000000000000;
	sram_mem[68546] = 16'b0000000000000000;
	sram_mem[68547] = 16'b0000000000000000;
	sram_mem[68548] = 16'b0000000000000000;
	sram_mem[68549] = 16'b0000000000000000;
	sram_mem[68550] = 16'b0000000000000000;
	sram_mem[68551] = 16'b0000000000000000;
	sram_mem[68552] = 16'b0000000000000000;
	sram_mem[68553] = 16'b0000000000000000;
	sram_mem[68554] = 16'b0000000000000000;
	sram_mem[68555] = 16'b0000000000000000;
	sram_mem[68556] = 16'b0000000000000000;
	sram_mem[68557] = 16'b0000000000000000;
	sram_mem[68558] = 16'b0000000000000000;
	sram_mem[68559] = 16'b0000000000000000;
	sram_mem[68560] = 16'b0000000000000000;
	sram_mem[68561] = 16'b0000000000000000;
	sram_mem[68562] = 16'b0000000000000000;
	sram_mem[68563] = 16'b0000000000000000;
	sram_mem[68564] = 16'b0000000000000000;
	sram_mem[68565] = 16'b0000000000000000;
	sram_mem[68566] = 16'b0000000000000000;
	sram_mem[68567] = 16'b0000000000000000;
	sram_mem[68568] = 16'b0000000000000000;
	sram_mem[68569] = 16'b0000000000000000;
	sram_mem[68570] = 16'b0000000000000000;
	sram_mem[68571] = 16'b0000000000000000;
	sram_mem[68572] = 16'b0000000000000000;
	sram_mem[68573] = 16'b0000000000000000;
	sram_mem[68574] = 16'b0000000000000000;
	sram_mem[68575] = 16'b0000000000000000;
	sram_mem[68576] = 16'b0000000000000000;
	sram_mem[68577] = 16'b0000000000000000;
	sram_mem[68578] = 16'b0000000000000000;
	sram_mem[68579] = 16'b0000000000000000;
	sram_mem[68580] = 16'b0000000000000000;
	sram_mem[68581] = 16'b0000000000000000;
	sram_mem[68582] = 16'b0000000000000000;
	sram_mem[68583] = 16'b0000000000000000;
	sram_mem[68584] = 16'b0000000000000000;
	sram_mem[68585] = 16'b0000000000000000;
	sram_mem[68586] = 16'b0000000000000000;
	sram_mem[68587] = 16'b0000000000000000;
	sram_mem[68588] = 16'b0000000000000000;
	sram_mem[68589] = 16'b0000000000000000;
	sram_mem[68590] = 16'b0000000000000000;
	sram_mem[68591] = 16'b0000000000000000;
	sram_mem[68592] = 16'b0000000000000000;
	sram_mem[68593] = 16'b0000000000000000;
	sram_mem[68594] = 16'b0000000000000000;
	sram_mem[68595] = 16'b0000000000000000;
	sram_mem[68596] = 16'b0000000000000000;
	sram_mem[68597] = 16'b0000000000000000;
	sram_mem[68598] = 16'b0000000000000000;
	sram_mem[68599] = 16'b0000000000000000;
	sram_mem[68600] = 16'b0000000000000000;
	sram_mem[68601] = 16'b0000000000000000;
	sram_mem[68602] = 16'b0000000000000000;
	sram_mem[68603] = 16'b0000000000000000;
	sram_mem[68604] = 16'b0000000000000000;
	sram_mem[68605] = 16'b0000000000000000;
	sram_mem[68606] = 16'b0000000000000000;
	sram_mem[68607] = 16'b0000000000000000;
	sram_mem[68608] = 16'b0000000000000000;
	sram_mem[68609] = 16'b0000000000000000;
	sram_mem[68610] = 16'b0000000000000000;
	sram_mem[68611] = 16'b0000000000000000;
	sram_mem[68612] = 16'b0000000000000000;
	sram_mem[68613] = 16'b0000000000000000;
	sram_mem[68614] = 16'b0000000000000000;
	sram_mem[68615] = 16'b0000000000000000;
	sram_mem[68616] = 16'b0000000000000000;
	sram_mem[68617] = 16'b0000000000000000;
	sram_mem[68618] = 16'b0000000000000000;
	sram_mem[68619] = 16'b0000000000000000;
	sram_mem[68620] = 16'b0000000000000000;
	sram_mem[68621] = 16'b0000000000000000;
	sram_mem[68622] = 16'b0000000000000000;
	sram_mem[68623] = 16'b0000000000000000;
	sram_mem[68624] = 16'b0000000000000000;
	sram_mem[68625] = 16'b0000000000000000;
	sram_mem[68626] = 16'b0000000000000000;
	sram_mem[68627] = 16'b0000000000000000;
	sram_mem[68628] = 16'b0000000000000000;
	sram_mem[68629] = 16'b0000000000000000;
	sram_mem[68630] = 16'b0000000000000000;
	sram_mem[68631] = 16'b0000000000000000;
	sram_mem[68632] = 16'b0000000000000000;
	sram_mem[68633] = 16'b0000000000000000;
	sram_mem[68634] = 16'b0000000000000000;
	sram_mem[68635] = 16'b0000000000000000;
	sram_mem[68636] = 16'b0000000000000000;
	sram_mem[68637] = 16'b0000000000000000;
	sram_mem[68638] = 16'b0000000000000000;
	sram_mem[68639] = 16'b0000000000000000;
	sram_mem[68640] = 16'b0000000000000000;
	sram_mem[68641] = 16'b0000000000000000;
	sram_mem[68642] = 16'b0000000000000000;
	sram_mem[68643] = 16'b0000000000000000;
	sram_mem[68644] = 16'b0000000000000000;
	sram_mem[68645] = 16'b0000000000000000;
	sram_mem[68646] = 16'b0000000000000000;
	sram_mem[68647] = 16'b0000000000000000;
	sram_mem[68648] = 16'b0000000000000000;
	sram_mem[68649] = 16'b0000000000000000;
	sram_mem[68650] = 16'b0000000000000000;
	sram_mem[68651] = 16'b0000000000000000;
	sram_mem[68652] = 16'b0000000000000000;
	sram_mem[68653] = 16'b0000000000000000;
	sram_mem[68654] = 16'b0000000000000000;
	sram_mem[68655] = 16'b0000000000000000;
	sram_mem[68656] = 16'b0000000000000000;
	sram_mem[68657] = 16'b0000000000000000;
	sram_mem[68658] = 16'b0000000000000000;
	sram_mem[68659] = 16'b0000000000000000;
	sram_mem[68660] = 16'b0000000000000000;
	sram_mem[68661] = 16'b0000000000000000;
	sram_mem[68662] = 16'b0000000000000000;
	sram_mem[68663] = 16'b0000000000000000;
	sram_mem[68664] = 16'b0000000000000000;
	sram_mem[68665] = 16'b0000000000000000;
	sram_mem[68666] = 16'b0000000000000000;
	sram_mem[68667] = 16'b0000000000000000;
	sram_mem[68668] = 16'b0000000000000000;
	sram_mem[68669] = 16'b0000000000000000;
	sram_mem[68670] = 16'b0000000000000000;
	sram_mem[68671] = 16'b0000000000000000;
	sram_mem[68672] = 16'b0000000000000000;
	sram_mem[68673] = 16'b0000000000000000;
	sram_mem[68674] = 16'b0000000000000000;
	sram_mem[68675] = 16'b0000000000000000;
	sram_mem[68676] = 16'b0000000000000000;
	sram_mem[68677] = 16'b0000000000000000;
	sram_mem[68678] = 16'b0000000000000000;
	sram_mem[68679] = 16'b0000000000000000;
	sram_mem[68680] = 16'b0000000000000000;
	sram_mem[68681] = 16'b0000000000000000;
	sram_mem[68682] = 16'b0000000000000000;
	sram_mem[68683] = 16'b0000000000000000;
	sram_mem[68684] = 16'b0000000000000000;
	sram_mem[68685] = 16'b0000000000000000;
	sram_mem[68686] = 16'b0000000000000000;
	sram_mem[68687] = 16'b0000000000000000;
	sram_mem[68688] = 16'b0000000000000000;
	sram_mem[68689] = 16'b0000000000000000;
	sram_mem[68690] = 16'b0000000000000000;
	sram_mem[68691] = 16'b0000000000000000;
	sram_mem[68692] = 16'b0000000000000000;
	sram_mem[68693] = 16'b0000000000000000;
	sram_mem[68694] = 16'b0000000000000000;
	sram_mem[68695] = 16'b0000000000000000;
	sram_mem[68696] = 16'b0000000000000000;
	sram_mem[68697] = 16'b0000000000000000;
	sram_mem[68698] = 16'b0000000000000000;
	sram_mem[68699] = 16'b0000000000000000;
	sram_mem[68700] = 16'b0000000000000000;
	sram_mem[68701] = 16'b0000000000000000;
	sram_mem[68702] = 16'b0000000000000000;
	sram_mem[68703] = 16'b0000000000000000;
	sram_mem[68704] = 16'b0000000000000000;
	sram_mem[68705] = 16'b0000000000000000;
	sram_mem[68706] = 16'b0000000000000000;
	sram_mem[68707] = 16'b0000000000000000;
	sram_mem[68708] = 16'b0000000000000000;
	sram_mem[68709] = 16'b0000000000000000;
	sram_mem[68710] = 16'b0000000000000000;
	sram_mem[68711] = 16'b0000000000000000;
	sram_mem[68712] = 16'b0000000000000000;
	sram_mem[68713] = 16'b0000000000000000;
	sram_mem[68714] = 16'b0000000000000000;
	sram_mem[68715] = 16'b0000000000000000;
	sram_mem[68716] = 16'b0000000000000000;
	sram_mem[68717] = 16'b0000000000000000;
	sram_mem[68718] = 16'b0000000000000000;
	sram_mem[68719] = 16'b0000000000000000;
	sram_mem[68720] = 16'b0000000000000000;
	sram_mem[68721] = 16'b0000000000000000;
	sram_mem[68722] = 16'b0000000000000000;
	sram_mem[68723] = 16'b0000000000000000;
	sram_mem[68724] = 16'b0000000000000000;
	sram_mem[68725] = 16'b0000000000000000;
	sram_mem[68726] = 16'b0000000000000000;
	sram_mem[68727] = 16'b0000000000000000;
	sram_mem[68728] = 16'b0000000000000000;
	sram_mem[68729] = 16'b0000000000000000;
	sram_mem[68730] = 16'b0000000000000000;
	sram_mem[68731] = 16'b0000000000000000;
	sram_mem[68732] = 16'b0000000000000000;
	sram_mem[68733] = 16'b0000000000000000;
	sram_mem[68734] = 16'b0000000000000000;
	sram_mem[68735] = 16'b0000000000000000;
	sram_mem[68736] = 16'b0000000000000000;
	sram_mem[68737] = 16'b0000000000000000;
	sram_mem[68738] = 16'b0000000000000000;
	sram_mem[68739] = 16'b0000000000000000;
	sram_mem[68740] = 16'b0000000000000000;
	sram_mem[68741] = 16'b0000000000000000;
	sram_mem[68742] = 16'b0000000000000000;
	sram_mem[68743] = 16'b0000000000000000;
	sram_mem[68744] = 16'b0000000000000000;
	sram_mem[68745] = 16'b0000000000000000;
	sram_mem[68746] = 16'b0000000000000000;
	sram_mem[68747] = 16'b0000000000000000;
	sram_mem[68748] = 16'b0000000000000000;
	sram_mem[68749] = 16'b0000000000000000;
	sram_mem[68750] = 16'b0000000000000000;
	sram_mem[68751] = 16'b0000000000000000;
	sram_mem[68752] = 16'b0000000000000000;
	sram_mem[68753] = 16'b0000000000000000;
	sram_mem[68754] = 16'b0000000000000000;
	sram_mem[68755] = 16'b0000000000000000;
	sram_mem[68756] = 16'b0000000000000000;
	sram_mem[68757] = 16'b0000000000000000;
	sram_mem[68758] = 16'b0000000000000000;
	sram_mem[68759] = 16'b0000000000000000;
	sram_mem[68760] = 16'b0000000000000000;
	sram_mem[68761] = 16'b0000000000000000;
	sram_mem[68762] = 16'b0000000000000000;
	sram_mem[68763] = 16'b0000000000000000;
	sram_mem[68764] = 16'b0000000000000000;
	sram_mem[68765] = 16'b0000000000000000;
	sram_mem[68766] = 16'b0000000000000000;
	sram_mem[68767] = 16'b0000000000000000;
	sram_mem[68768] = 16'b0000000000000000;
	sram_mem[68769] = 16'b0000000000000000;
	sram_mem[68770] = 16'b0000000000000000;
	sram_mem[68771] = 16'b0000000000000000;
	sram_mem[68772] = 16'b0000000000000000;
	sram_mem[68773] = 16'b0000000000000000;
	sram_mem[68774] = 16'b0000000000000000;
	sram_mem[68775] = 16'b0000000000000000;
	sram_mem[68776] = 16'b0000000000000000;
	sram_mem[68777] = 16'b0000000000000000;
	sram_mem[68778] = 16'b0000000000000000;
	sram_mem[68779] = 16'b0000000000000000;
	sram_mem[68780] = 16'b0000000000000000;
	sram_mem[68781] = 16'b0000000000000000;
	sram_mem[68782] = 16'b0000000000000000;
	sram_mem[68783] = 16'b0000000000000000;
	sram_mem[68784] = 16'b0000000000000000;
	sram_mem[68785] = 16'b0000000000000000;
	sram_mem[68786] = 16'b0000000000000000;
	sram_mem[68787] = 16'b0000000000000000;
	sram_mem[68788] = 16'b0000000000000000;
	sram_mem[68789] = 16'b0000000000000000;
	sram_mem[68790] = 16'b0000000000000000;
	sram_mem[68791] = 16'b0000000000000000;
	sram_mem[68792] = 16'b0000000000000000;
	sram_mem[68793] = 16'b0000000000000000;
	sram_mem[68794] = 16'b0000000000000000;
	sram_mem[68795] = 16'b0000000000000000;
	sram_mem[68796] = 16'b0000000000000000;
	sram_mem[68797] = 16'b0000000000000000;
	sram_mem[68798] = 16'b0000000000000000;
	sram_mem[68799] = 16'b0000000000000000;
	sram_mem[68800] = 16'b0000000000000000;
	sram_mem[68801] = 16'b0000000000000000;
	sram_mem[68802] = 16'b0000000000000000;
	sram_mem[68803] = 16'b0000000000000000;
	sram_mem[68804] = 16'b0000000000000000;
	sram_mem[68805] = 16'b0000000000000000;
	sram_mem[68806] = 16'b0000000000000000;
	sram_mem[68807] = 16'b0000000000000000;
	sram_mem[68808] = 16'b0000000000000000;
	sram_mem[68809] = 16'b0000000000000000;
	sram_mem[68810] = 16'b0000000000000000;
	sram_mem[68811] = 16'b0000000000000000;
	sram_mem[68812] = 16'b0000000000000000;
	sram_mem[68813] = 16'b0000000000000000;
	sram_mem[68814] = 16'b0000000000000000;
	sram_mem[68815] = 16'b0000000000000000;
	sram_mem[68816] = 16'b0000000000000000;
	sram_mem[68817] = 16'b0000000000000000;
	sram_mem[68818] = 16'b0000000000000000;
	sram_mem[68819] = 16'b0000000000000000;
	sram_mem[68820] = 16'b0000000000000000;
	sram_mem[68821] = 16'b0000000000000000;
	sram_mem[68822] = 16'b0000000000000000;
	sram_mem[68823] = 16'b0000000000000000;
	sram_mem[68824] = 16'b0000000000000000;
	sram_mem[68825] = 16'b0000000000000000;
	sram_mem[68826] = 16'b0000000000000000;
	sram_mem[68827] = 16'b0000000000000000;
	sram_mem[68828] = 16'b0000000000000000;
	sram_mem[68829] = 16'b0000000000000000;
	sram_mem[68830] = 16'b0000000000000000;
	sram_mem[68831] = 16'b0000000000000000;
	sram_mem[68832] = 16'b0000000000000000;
	sram_mem[68833] = 16'b0000000000000000;
	sram_mem[68834] = 16'b0000000000000000;
	sram_mem[68835] = 16'b0000000000000000;
	sram_mem[68836] = 16'b0000000000000000;
	sram_mem[68837] = 16'b0000000000000000;
	sram_mem[68838] = 16'b0000000000000000;
	sram_mem[68839] = 16'b0000000000000000;
	sram_mem[68840] = 16'b0000000000000000;
	sram_mem[68841] = 16'b0000000000000000;
	sram_mem[68842] = 16'b0000000000000000;
	sram_mem[68843] = 16'b0000000000000000;
	sram_mem[68844] = 16'b0000000000000000;
	sram_mem[68845] = 16'b0000000000000000;
	sram_mem[68846] = 16'b0000000000000000;
	sram_mem[68847] = 16'b0000000000000000;
	sram_mem[68848] = 16'b0000000000000000;
	sram_mem[68849] = 16'b0000000000000000;
	sram_mem[68850] = 16'b0000000000000000;
	sram_mem[68851] = 16'b0000000000000000;
	sram_mem[68852] = 16'b0000000000000000;
	sram_mem[68853] = 16'b0000000000000000;
	sram_mem[68854] = 16'b0000000000000000;
	sram_mem[68855] = 16'b0000000000000000;
	sram_mem[68856] = 16'b0000000000000000;
	sram_mem[68857] = 16'b0000000000000000;
	sram_mem[68858] = 16'b0000000000000000;
	sram_mem[68859] = 16'b0000000000000000;
	sram_mem[68860] = 16'b0000000000000000;
	sram_mem[68861] = 16'b0000000000000000;
	sram_mem[68862] = 16'b0000000000000000;
	sram_mem[68863] = 16'b0000000000000000;
	sram_mem[68864] = 16'b0000000000000000;
	sram_mem[68865] = 16'b0000000000000000;
	sram_mem[68866] = 16'b0000000000000000;
	sram_mem[68867] = 16'b0000000000000000;
	sram_mem[68868] = 16'b0000000000000000;
	sram_mem[68869] = 16'b0000000000000000;
	sram_mem[68870] = 16'b0000000000000000;
	sram_mem[68871] = 16'b0000000000000000;
	sram_mem[68872] = 16'b0000000000000000;
	sram_mem[68873] = 16'b0000000000000000;
	sram_mem[68874] = 16'b0000000000000000;
	sram_mem[68875] = 16'b0000000000000000;
	sram_mem[68876] = 16'b0000000000000000;
	sram_mem[68877] = 16'b0000000000000000;
	sram_mem[68878] = 16'b0000000000000000;
	sram_mem[68879] = 16'b0000000000000000;
	sram_mem[68880] = 16'b0000000000000000;
	sram_mem[68881] = 16'b0000000000000000;
	sram_mem[68882] = 16'b0000000000000000;
	sram_mem[68883] = 16'b0000000000000000;
	sram_mem[68884] = 16'b0000000000000000;
	sram_mem[68885] = 16'b0000000000000000;
	sram_mem[68886] = 16'b0000000000000000;
	sram_mem[68887] = 16'b0000000000000000;
	sram_mem[68888] = 16'b0000000000000000;
	sram_mem[68889] = 16'b0000000000000000;
	sram_mem[68890] = 16'b0000000000000000;
	sram_mem[68891] = 16'b0000000000000000;
	sram_mem[68892] = 16'b0000000000000000;
	sram_mem[68893] = 16'b0000000000000000;
	sram_mem[68894] = 16'b0000000000000000;
	sram_mem[68895] = 16'b0000000000000000;
	sram_mem[68896] = 16'b0000000000000000;
	sram_mem[68897] = 16'b0000000000000000;
	sram_mem[68898] = 16'b0000000000000000;
	sram_mem[68899] = 16'b0000000000000000;
	sram_mem[68900] = 16'b0000000000000000;
	sram_mem[68901] = 16'b0000000000000000;
	sram_mem[68902] = 16'b0000000000000000;
	sram_mem[68903] = 16'b0000000000000000;
	sram_mem[68904] = 16'b0000000000000000;
	sram_mem[68905] = 16'b0000000000000000;
	sram_mem[68906] = 16'b0000000000000000;
	sram_mem[68907] = 16'b0000000000000000;
	sram_mem[68908] = 16'b0000000000000000;
	sram_mem[68909] = 16'b0000000000000000;
	sram_mem[68910] = 16'b0000000000000000;
	sram_mem[68911] = 16'b0000000000000000;
	sram_mem[68912] = 16'b0000000000000000;
	sram_mem[68913] = 16'b0000000000000000;
	sram_mem[68914] = 16'b0000000000000000;
	sram_mem[68915] = 16'b0000000000000000;
	sram_mem[68916] = 16'b0000000000000000;
	sram_mem[68917] = 16'b0000000000000000;
	sram_mem[68918] = 16'b0000000000000000;
	sram_mem[68919] = 16'b0000000000000000;
	sram_mem[68920] = 16'b0000000000000000;
	sram_mem[68921] = 16'b0000000000000000;
	sram_mem[68922] = 16'b0000000000000000;
	sram_mem[68923] = 16'b0000000000000000;
	sram_mem[68924] = 16'b0000000000000000;
	sram_mem[68925] = 16'b0000000000000000;
	sram_mem[68926] = 16'b0000000000000000;
	sram_mem[68927] = 16'b0000000000000000;
	sram_mem[68928] = 16'b0000000000000000;
	sram_mem[68929] = 16'b0000000000000000;
	sram_mem[68930] = 16'b0000000000000000;
	sram_mem[68931] = 16'b0000000000000000;
	sram_mem[68932] = 16'b0000000000000000;
	sram_mem[68933] = 16'b0000000000000000;
	sram_mem[68934] = 16'b0000000000000000;
	sram_mem[68935] = 16'b0000000000000000;
	sram_mem[68936] = 16'b0000000000000000;
	sram_mem[68937] = 16'b0000000000000000;
	sram_mem[68938] = 16'b0000000000000000;
	sram_mem[68939] = 16'b0000000000000000;
	sram_mem[68940] = 16'b0000000000000000;
	sram_mem[68941] = 16'b0000000000000000;
	sram_mem[68942] = 16'b0000000000000000;
	sram_mem[68943] = 16'b0000000000000000;
	sram_mem[68944] = 16'b0000000000000000;
	sram_mem[68945] = 16'b0000000000000000;
	sram_mem[68946] = 16'b0000000000000000;
	sram_mem[68947] = 16'b0000000000000000;
	sram_mem[68948] = 16'b0000000000000000;
	sram_mem[68949] = 16'b0000000000000000;
	sram_mem[68950] = 16'b0000000000000000;
	sram_mem[68951] = 16'b0000000000000000;
	sram_mem[68952] = 16'b0000000000000000;
	sram_mem[68953] = 16'b0000000000000000;
	sram_mem[68954] = 16'b0000000000000000;
	sram_mem[68955] = 16'b0000000000000000;
	sram_mem[68956] = 16'b0000000000000000;
	sram_mem[68957] = 16'b0000000000000000;
	sram_mem[68958] = 16'b0000000000000000;
	sram_mem[68959] = 16'b0000000000000000;
	sram_mem[68960] = 16'b0000000000000000;
	sram_mem[68961] = 16'b0000000000000000;
	sram_mem[68962] = 16'b0000000000000000;
	sram_mem[68963] = 16'b0000000000000000;
	sram_mem[68964] = 16'b0000000000000000;
	sram_mem[68965] = 16'b0000000000000000;
	sram_mem[68966] = 16'b0000000000000000;
	sram_mem[68967] = 16'b0000000000000000;
	sram_mem[68968] = 16'b0000000000000000;
	sram_mem[68969] = 16'b0000000000000000;
	sram_mem[68970] = 16'b0000000000000000;
	sram_mem[68971] = 16'b0000000000000000;
	sram_mem[68972] = 16'b0000000000000000;
	sram_mem[68973] = 16'b0000000000000000;
	sram_mem[68974] = 16'b0000000000000000;
	sram_mem[68975] = 16'b0000000000000000;
	sram_mem[68976] = 16'b0000000000000000;
	sram_mem[68977] = 16'b0000000000000000;
	sram_mem[68978] = 16'b0000000000000000;
	sram_mem[68979] = 16'b0000000000000000;
	sram_mem[68980] = 16'b0000000000000000;
	sram_mem[68981] = 16'b0000000000000000;
	sram_mem[68982] = 16'b0000000000000000;
	sram_mem[68983] = 16'b0000000000000000;
	sram_mem[68984] = 16'b0000000000000000;
	sram_mem[68985] = 16'b0000000000000000;
	sram_mem[68986] = 16'b0000000000000000;
	sram_mem[68987] = 16'b0000000000000000;
	sram_mem[68988] = 16'b0000000000000000;
	sram_mem[68989] = 16'b0000000000000000;
	sram_mem[68990] = 16'b0000000000000000;
	sram_mem[68991] = 16'b0000000000000000;
	sram_mem[68992] = 16'b0000000000000000;
	sram_mem[68993] = 16'b0000000000000000;
	sram_mem[68994] = 16'b0000000000000000;
	sram_mem[68995] = 16'b0000000000000000;
	sram_mem[68996] = 16'b0000000000000000;
	sram_mem[68997] = 16'b0000000000000000;
	sram_mem[68998] = 16'b0000000000000000;
	sram_mem[68999] = 16'b0000000000000000;
	sram_mem[69000] = 16'b0000000000000000;
	sram_mem[69001] = 16'b0000000000000000;
	sram_mem[69002] = 16'b0000000000000000;
	sram_mem[69003] = 16'b0000000000000000;
	sram_mem[69004] = 16'b0000000000000000;
	sram_mem[69005] = 16'b0000000000000000;
	sram_mem[69006] = 16'b0000000000000000;
	sram_mem[69007] = 16'b0000000000000000;
	sram_mem[69008] = 16'b0000000000000000;
	sram_mem[69009] = 16'b0000000000000000;
	sram_mem[69010] = 16'b0000000000000000;
	sram_mem[69011] = 16'b0000000000000000;
	sram_mem[69012] = 16'b0000000000000000;
	sram_mem[69013] = 16'b0000000000000000;
	sram_mem[69014] = 16'b0000000000000000;
	sram_mem[69015] = 16'b0000000000000000;
	sram_mem[69016] = 16'b0000000000000000;
	sram_mem[69017] = 16'b0000000000000000;
	sram_mem[69018] = 16'b0000000000000000;
	sram_mem[69019] = 16'b0000000000000000;
	sram_mem[69020] = 16'b0000000000000000;
	sram_mem[69021] = 16'b0000000000000000;
	sram_mem[69022] = 16'b0000000000000000;
	sram_mem[69023] = 16'b0000000000000000;
	sram_mem[69024] = 16'b0000000000000000;
	sram_mem[69025] = 16'b0000000000000000;
	sram_mem[69026] = 16'b0000000000000000;
	sram_mem[69027] = 16'b0000000000000000;
	sram_mem[69028] = 16'b0000000000000000;
	sram_mem[69029] = 16'b0000000000000000;
	sram_mem[69030] = 16'b0000000000000000;
	sram_mem[69031] = 16'b0000000000000000;
	sram_mem[69032] = 16'b0000000000000000;
	sram_mem[69033] = 16'b0000000000000000;
	sram_mem[69034] = 16'b0000000000000000;
	sram_mem[69035] = 16'b0000000000000000;
	sram_mem[69036] = 16'b0000000000000000;
	sram_mem[69037] = 16'b0000000000000000;
	sram_mem[69038] = 16'b0000000000000000;
	sram_mem[69039] = 16'b0000000000000000;
	sram_mem[69040] = 16'b0000000000000000;
	sram_mem[69041] = 16'b0000000000000000;
	sram_mem[69042] = 16'b0000000000000000;
	sram_mem[69043] = 16'b0000000000000000;
	sram_mem[69044] = 16'b0000000000000000;
	sram_mem[69045] = 16'b0000000000000000;
	sram_mem[69046] = 16'b0000000000000000;
	sram_mem[69047] = 16'b0000000000000000;
	sram_mem[69048] = 16'b0000000000000000;
	sram_mem[69049] = 16'b0000000000000000;
	sram_mem[69050] = 16'b0000000000000000;
	sram_mem[69051] = 16'b0000000000000000;
	sram_mem[69052] = 16'b0000000000000000;
	sram_mem[69053] = 16'b0000000000000000;
	sram_mem[69054] = 16'b0000000000000000;
	sram_mem[69055] = 16'b0000000000000000;
	sram_mem[69056] = 16'b0000000000000000;
	sram_mem[69057] = 16'b0000000000000000;
	sram_mem[69058] = 16'b0000000000000000;
	sram_mem[69059] = 16'b0000000000000000;
	sram_mem[69060] = 16'b0000000000000000;
	sram_mem[69061] = 16'b0000000000000000;
	sram_mem[69062] = 16'b0000000000000000;
	sram_mem[69063] = 16'b0000000000000000;
	sram_mem[69064] = 16'b0000000000000000;
	sram_mem[69065] = 16'b0000000000000000;
	sram_mem[69066] = 16'b0000000000000000;
	sram_mem[69067] = 16'b0000000000000000;
	sram_mem[69068] = 16'b0000000000000000;
	sram_mem[69069] = 16'b0000000000000000;
	sram_mem[69070] = 16'b0000000000000000;
	sram_mem[69071] = 16'b0000000000000000;
	sram_mem[69072] = 16'b0000000000000000;
	sram_mem[69073] = 16'b0000000000000000;
	sram_mem[69074] = 16'b0000000000000000;
	sram_mem[69075] = 16'b0000000000000000;
	sram_mem[69076] = 16'b0000000000000000;
	sram_mem[69077] = 16'b0000000000000000;
	sram_mem[69078] = 16'b0000000000000000;
	sram_mem[69079] = 16'b0000000000000000;
	sram_mem[69080] = 16'b0000000000000000;
	sram_mem[69081] = 16'b0000000000000000;
	sram_mem[69082] = 16'b0000000000000000;
	sram_mem[69083] = 16'b0000000000000000;
	sram_mem[69084] = 16'b0000000000000000;
	sram_mem[69085] = 16'b0000000000000000;
	sram_mem[69086] = 16'b0000000000000000;
	sram_mem[69087] = 16'b0000000000000000;
	sram_mem[69088] = 16'b0000000000000000;
	sram_mem[69089] = 16'b0000000000000000;
	sram_mem[69090] = 16'b0000000000000000;
	sram_mem[69091] = 16'b0000000000000000;
	sram_mem[69092] = 16'b0000000000000000;
	sram_mem[69093] = 16'b0000000000000000;
	sram_mem[69094] = 16'b0000000000000000;
	sram_mem[69095] = 16'b0000000000000000;
	sram_mem[69096] = 16'b0000000000000000;
	sram_mem[69097] = 16'b0000000000000000;
	sram_mem[69098] = 16'b0000000000000000;
	sram_mem[69099] = 16'b0000000000000000;
	sram_mem[69100] = 16'b0000000000000000;
	sram_mem[69101] = 16'b0000000000000000;
	sram_mem[69102] = 16'b0000000000000000;
	sram_mem[69103] = 16'b0000000000000000;
	sram_mem[69104] = 16'b0000000000000000;
	sram_mem[69105] = 16'b0000000000000000;
	sram_mem[69106] = 16'b0000000000000000;
	sram_mem[69107] = 16'b0000000000000000;
	sram_mem[69108] = 16'b0000000000000000;
	sram_mem[69109] = 16'b0000000000000000;
	sram_mem[69110] = 16'b0000000000000000;
	sram_mem[69111] = 16'b0000000000000000;
	sram_mem[69112] = 16'b0000000000000000;
	sram_mem[69113] = 16'b0000000000000000;
	sram_mem[69114] = 16'b0000000000000000;
	sram_mem[69115] = 16'b0000000000000000;
	sram_mem[69116] = 16'b0000000000000000;
	sram_mem[69117] = 16'b0000000000000000;
	sram_mem[69118] = 16'b0000000000000000;
	sram_mem[69119] = 16'b0000000000000000;
	sram_mem[69120] = 16'b0000000000000000;
	sram_mem[69121] = 16'b0000000000000000;
	sram_mem[69122] = 16'b0000000000000000;
	sram_mem[69123] = 16'b0000000000000000;
	sram_mem[69124] = 16'b0000000000000000;
	sram_mem[69125] = 16'b0000000000000000;
	sram_mem[69126] = 16'b0000000000000000;
	sram_mem[69127] = 16'b0000000000000000;
	sram_mem[69128] = 16'b0000000000000000;
	sram_mem[69129] = 16'b0000000000000000;
	sram_mem[69130] = 16'b0000000000000000;
	sram_mem[69131] = 16'b0000000000000000;
	sram_mem[69132] = 16'b0000000000000000;
	sram_mem[69133] = 16'b0000000000000000;
	sram_mem[69134] = 16'b0000000000000000;
	sram_mem[69135] = 16'b0000000000000000;
	sram_mem[69136] = 16'b0000000000000000;
	sram_mem[69137] = 16'b0000000000000000;
	sram_mem[69138] = 16'b0000000000000000;
	sram_mem[69139] = 16'b0000000000000000;
	sram_mem[69140] = 16'b0000000000000000;
	sram_mem[69141] = 16'b0000000000000000;
	sram_mem[69142] = 16'b0000000000000000;
	sram_mem[69143] = 16'b0000000000000000;
	sram_mem[69144] = 16'b0000000000000000;
	sram_mem[69145] = 16'b0000000000000000;
	sram_mem[69146] = 16'b0000000000000000;
	sram_mem[69147] = 16'b0000000000000000;
	sram_mem[69148] = 16'b0000000000000000;
	sram_mem[69149] = 16'b0000000000000000;
	sram_mem[69150] = 16'b0000000000000000;
	sram_mem[69151] = 16'b0000000000000000;
	sram_mem[69152] = 16'b0000000000000000;
	sram_mem[69153] = 16'b0000000000000000;
	sram_mem[69154] = 16'b0000000000000000;
	sram_mem[69155] = 16'b0000000000000000;
	sram_mem[69156] = 16'b0000000000000000;
	sram_mem[69157] = 16'b0000000000000000;
	sram_mem[69158] = 16'b0000000000000000;
	sram_mem[69159] = 16'b0000000000000000;
	sram_mem[69160] = 16'b0000000000000000;
	sram_mem[69161] = 16'b0000000000000000;
	sram_mem[69162] = 16'b0000000000000000;
	sram_mem[69163] = 16'b0000000000000000;
	sram_mem[69164] = 16'b0000000000000000;
	sram_mem[69165] = 16'b0000000000000000;
	sram_mem[69166] = 16'b0000000000000000;
	sram_mem[69167] = 16'b0000000000000000;
	sram_mem[69168] = 16'b0000000000000000;
	sram_mem[69169] = 16'b0000000000000000;
	sram_mem[69170] = 16'b0000000000000000;
	sram_mem[69171] = 16'b0000000000000000;
	sram_mem[69172] = 16'b0000000000000000;
	sram_mem[69173] = 16'b0000000000000000;
	sram_mem[69174] = 16'b0000000000000000;
	sram_mem[69175] = 16'b0000000000000000;
	sram_mem[69176] = 16'b0000000000000000;
	sram_mem[69177] = 16'b0000000000000000;
	sram_mem[69178] = 16'b0000000000000000;
	sram_mem[69179] = 16'b0000000000000000;
	sram_mem[69180] = 16'b0000000000000000;
	sram_mem[69181] = 16'b0000000000000000;
	sram_mem[69182] = 16'b0000000000000000;
	sram_mem[69183] = 16'b0000000000000000;
	sram_mem[69184] = 16'b0000000000000000;
	sram_mem[69185] = 16'b0000000000000000;
	sram_mem[69186] = 16'b0000000000000000;
	sram_mem[69187] = 16'b0000000000000000;
	sram_mem[69188] = 16'b0000000000000000;
	sram_mem[69189] = 16'b0000000000000000;
	sram_mem[69190] = 16'b0000000000000000;
	sram_mem[69191] = 16'b0000000000000000;
	sram_mem[69192] = 16'b0000000000000000;
	sram_mem[69193] = 16'b0000000000000000;
	sram_mem[69194] = 16'b0000000000000000;
	sram_mem[69195] = 16'b0000000000000000;
	sram_mem[69196] = 16'b0000000000000000;
	sram_mem[69197] = 16'b0000000000000000;
	sram_mem[69198] = 16'b0000000000000000;
	sram_mem[69199] = 16'b0000000000000000;
	sram_mem[69200] = 16'b0000000000000000;
	sram_mem[69201] = 16'b0000000000000000;
	sram_mem[69202] = 16'b0000000000000000;
	sram_mem[69203] = 16'b0000000000000000;
	sram_mem[69204] = 16'b0000000000000000;
	sram_mem[69205] = 16'b0000000000000000;
	sram_mem[69206] = 16'b0000000000000000;
	sram_mem[69207] = 16'b0000000000000000;
	sram_mem[69208] = 16'b0000000000000000;
	sram_mem[69209] = 16'b0000000000000000;
	sram_mem[69210] = 16'b0000000000000000;
	sram_mem[69211] = 16'b0000000000000000;
	sram_mem[69212] = 16'b0000000000000000;
	sram_mem[69213] = 16'b0000000000000000;
	sram_mem[69214] = 16'b0000000000000000;
	sram_mem[69215] = 16'b0000000000000000;
	sram_mem[69216] = 16'b0000000000000000;
	sram_mem[69217] = 16'b0000000000000000;
	sram_mem[69218] = 16'b0000000000000000;
	sram_mem[69219] = 16'b0000000000000000;
	sram_mem[69220] = 16'b0000000000000000;
	sram_mem[69221] = 16'b0000000000000000;
	sram_mem[69222] = 16'b0000000000000000;
	sram_mem[69223] = 16'b0000000000000000;
	sram_mem[69224] = 16'b0000000000000000;
	sram_mem[69225] = 16'b0000000000000000;
	sram_mem[69226] = 16'b0000000000000000;
	sram_mem[69227] = 16'b0000000000000000;
	sram_mem[69228] = 16'b0000000000000000;
	sram_mem[69229] = 16'b0000000000000000;
	sram_mem[69230] = 16'b0000000000000000;
	sram_mem[69231] = 16'b0000000000000000;
	sram_mem[69232] = 16'b0000000000000000;
	sram_mem[69233] = 16'b0000000000000000;
	sram_mem[69234] = 16'b0000000000000000;
	sram_mem[69235] = 16'b0000000000000000;
	sram_mem[69236] = 16'b0000000000000000;
	sram_mem[69237] = 16'b0000000000000000;
	sram_mem[69238] = 16'b0000000000000000;
	sram_mem[69239] = 16'b0000000000000000;
	sram_mem[69240] = 16'b0000000000000000;
	sram_mem[69241] = 16'b0000000000000000;
	sram_mem[69242] = 16'b0000000000000000;
	sram_mem[69243] = 16'b0000000000000000;
	sram_mem[69244] = 16'b0000000000000000;
	sram_mem[69245] = 16'b0000000000000000;
	sram_mem[69246] = 16'b0000000000000000;
	sram_mem[69247] = 16'b0000000000000000;
	sram_mem[69248] = 16'b0000000000000000;
	sram_mem[69249] = 16'b0000000000000000;
	sram_mem[69250] = 16'b0000000000000000;
	sram_mem[69251] = 16'b0000000000000000;
	sram_mem[69252] = 16'b0000000000000000;
	sram_mem[69253] = 16'b0000000000000000;
	sram_mem[69254] = 16'b0000000000000000;
	sram_mem[69255] = 16'b0000000000000000;
	sram_mem[69256] = 16'b0000000000000000;
	sram_mem[69257] = 16'b0000000000000000;
	sram_mem[69258] = 16'b0000000000000000;
	sram_mem[69259] = 16'b0000000000000000;
	sram_mem[69260] = 16'b0000000000000000;
	sram_mem[69261] = 16'b0000000000000000;
	sram_mem[69262] = 16'b0000000000000000;
	sram_mem[69263] = 16'b0000000000000000;
	sram_mem[69264] = 16'b0000000000000000;
	sram_mem[69265] = 16'b0000000000000000;
	sram_mem[69266] = 16'b0000000000000000;
	sram_mem[69267] = 16'b0000000000000000;
	sram_mem[69268] = 16'b0000000000000000;
	sram_mem[69269] = 16'b0000000000000000;
	sram_mem[69270] = 16'b0000000000000000;
	sram_mem[69271] = 16'b0000000000000000;
	sram_mem[69272] = 16'b0000000000000000;
	sram_mem[69273] = 16'b0000000000000000;
	sram_mem[69274] = 16'b0000000000000000;
	sram_mem[69275] = 16'b0000000000000000;
	sram_mem[69276] = 16'b0000000000000000;
	sram_mem[69277] = 16'b0000000000000000;
	sram_mem[69278] = 16'b0000000000000000;
	sram_mem[69279] = 16'b0000000000000000;
	sram_mem[69280] = 16'b0000000000000000;
	sram_mem[69281] = 16'b0000000000000000;
	sram_mem[69282] = 16'b0000000000000000;
	sram_mem[69283] = 16'b0000000000000000;
	sram_mem[69284] = 16'b0000000000000000;
	sram_mem[69285] = 16'b0000000000000000;
	sram_mem[69286] = 16'b0000000000000000;
	sram_mem[69287] = 16'b0000000000000000;
	sram_mem[69288] = 16'b0000000000000000;
	sram_mem[69289] = 16'b0000000000000000;
	sram_mem[69290] = 16'b0000000000000000;
	sram_mem[69291] = 16'b0000000000000000;
	sram_mem[69292] = 16'b0000000000000000;
	sram_mem[69293] = 16'b0000000000000000;
	sram_mem[69294] = 16'b0000000000000000;
	sram_mem[69295] = 16'b0000000000000000;
	sram_mem[69296] = 16'b0000000000000000;
	sram_mem[69297] = 16'b0000000000000000;
	sram_mem[69298] = 16'b0000000000000000;
	sram_mem[69299] = 16'b0000000000000000;
	sram_mem[69300] = 16'b0000000000000000;
	sram_mem[69301] = 16'b0000000000000000;
	sram_mem[69302] = 16'b0000000000000000;
	sram_mem[69303] = 16'b0000000000000000;
	sram_mem[69304] = 16'b0000000000000000;
	sram_mem[69305] = 16'b0000000000000000;
	sram_mem[69306] = 16'b0000000000000000;
	sram_mem[69307] = 16'b0000000000000000;
	sram_mem[69308] = 16'b0000000000000000;
	sram_mem[69309] = 16'b0000000000000000;
	sram_mem[69310] = 16'b0000000000000000;
	sram_mem[69311] = 16'b0000000000000000;
	sram_mem[69312] = 16'b0000000000000000;
	sram_mem[69313] = 16'b0000000000000000;
	sram_mem[69314] = 16'b0000000000000000;
	sram_mem[69315] = 16'b0000000000000000;
	sram_mem[69316] = 16'b0000000000000000;
	sram_mem[69317] = 16'b0000000000000000;
	sram_mem[69318] = 16'b0000000000000000;
	sram_mem[69319] = 16'b0000000000000000;
	sram_mem[69320] = 16'b0000000000000000;
	sram_mem[69321] = 16'b0000000000000000;
	sram_mem[69322] = 16'b0000000000000000;
	sram_mem[69323] = 16'b0000000000000000;
	sram_mem[69324] = 16'b0000000000000000;
	sram_mem[69325] = 16'b0000000000000000;
	sram_mem[69326] = 16'b0000000000000000;
	sram_mem[69327] = 16'b0000000000000000;
	sram_mem[69328] = 16'b0000000000000000;
	sram_mem[69329] = 16'b0000000000000000;
	sram_mem[69330] = 16'b0000000000000000;
	sram_mem[69331] = 16'b0000000000000000;
	sram_mem[69332] = 16'b0000000000000000;
	sram_mem[69333] = 16'b0000000000000000;
	sram_mem[69334] = 16'b0000000000000000;
	sram_mem[69335] = 16'b0000000000000000;
	sram_mem[69336] = 16'b0000000000000000;
	sram_mem[69337] = 16'b0000000000000000;
	sram_mem[69338] = 16'b0000000000000000;
	sram_mem[69339] = 16'b0000000000000000;
	sram_mem[69340] = 16'b0000000000000000;
	sram_mem[69341] = 16'b0000000000000000;
	sram_mem[69342] = 16'b0000000000000000;
	sram_mem[69343] = 16'b0000000000000000;
	sram_mem[69344] = 16'b0000000000000000;
	sram_mem[69345] = 16'b0000000000000000;
	sram_mem[69346] = 16'b0000000000000000;
	sram_mem[69347] = 16'b0000000000000000;
	sram_mem[69348] = 16'b0000000000000000;
	sram_mem[69349] = 16'b0000000000000000;
	sram_mem[69350] = 16'b0000000000000000;
	sram_mem[69351] = 16'b0000000000000000;
	sram_mem[69352] = 16'b0000000000000000;
	sram_mem[69353] = 16'b0000000000000000;
	sram_mem[69354] = 16'b0000000000000000;
	sram_mem[69355] = 16'b0000000000000000;
	sram_mem[69356] = 16'b0000000000000000;
	sram_mem[69357] = 16'b0000000000000000;
	sram_mem[69358] = 16'b0000000000000000;
	sram_mem[69359] = 16'b0000000000000000;
	sram_mem[69360] = 16'b0000000000000000;
	sram_mem[69361] = 16'b0000000000000000;
	sram_mem[69362] = 16'b0000000000000000;
	sram_mem[69363] = 16'b0000000000000000;
	sram_mem[69364] = 16'b0000000000000000;
	sram_mem[69365] = 16'b0000000000000000;
	sram_mem[69366] = 16'b0000000000000000;
	sram_mem[69367] = 16'b0000000000000000;
	sram_mem[69368] = 16'b0000000000000000;
	sram_mem[69369] = 16'b0000000000000000;
	sram_mem[69370] = 16'b0000000000000000;
	sram_mem[69371] = 16'b0000000000000000;
	sram_mem[69372] = 16'b0000000000000000;
	sram_mem[69373] = 16'b0000000000000000;
	sram_mem[69374] = 16'b0000000000000000;
	sram_mem[69375] = 16'b0000000000000000;
	sram_mem[69376] = 16'b0000000000000000;
	sram_mem[69377] = 16'b0000000000000000;
	sram_mem[69378] = 16'b0000000000000000;
	sram_mem[69379] = 16'b0000000000000000;
	sram_mem[69380] = 16'b0000000000000000;
	sram_mem[69381] = 16'b0000000000000000;
	sram_mem[69382] = 16'b0000000000000000;
	sram_mem[69383] = 16'b0000000000000000;
	sram_mem[69384] = 16'b0000000000000000;
	sram_mem[69385] = 16'b0000000000000000;
	sram_mem[69386] = 16'b0000000000000000;
	sram_mem[69387] = 16'b0000000000000000;
	sram_mem[69388] = 16'b0000000000000000;
	sram_mem[69389] = 16'b0000000000000000;
	sram_mem[69390] = 16'b0000000000000000;
	sram_mem[69391] = 16'b0000000000000000;
	sram_mem[69392] = 16'b0000000000000000;
	sram_mem[69393] = 16'b0000000000000000;
	sram_mem[69394] = 16'b0000000000000000;
	sram_mem[69395] = 16'b0000000000000000;
	sram_mem[69396] = 16'b0000000000000000;
	sram_mem[69397] = 16'b0000000000000000;
	sram_mem[69398] = 16'b0000000000000000;
	sram_mem[69399] = 16'b0000000000000000;
	sram_mem[69400] = 16'b0000000000000000;
	sram_mem[69401] = 16'b0000000000000000;
	sram_mem[69402] = 16'b0000000000000000;
	sram_mem[69403] = 16'b0000000000000000;
	sram_mem[69404] = 16'b0000000000000000;
	sram_mem[69405] = 16'b0000000000000000;
	sram_mem[69406] = 16'b0000000000000000;
	sram_mem[69407] = 16'b0000000000000000;
	sram_mem[69408] = 16'b0000000000000000;
	sram_mem[69409] = 16'b0000000000000000;
	sram_mem[69410] = 16'b0000000000000000;
	sram_mem[69411] = 16'b0000000000000000;
	sram_mem[69412] = 16'b0000000000000000;
	sram_mem[69413] = 16'b0000000000000000;
	sram_mem[69414] = 16'b0000000000000000;
	sram_mem[69415] = 16'b0000000000000000;
	sram_mem[69416] = 16'b0000000000000000;
	sram_mem[69417] = 16'b0000000000000000;
	sram_mem[69418] = 16'b0000000000000000;
	sram_mem[69419] = 16'b0000000000000000;
	sram_mem[69420] = 16'b0000000000000000;
	sram_mem[69421] = 16'b0000000000000000;
	sram_mem[69422] = 16'b0000000000000000;
	sram_mem[69423] = 16'b0000000000000000;
	sram_mem[69424] = 16'b0000000000000000;
	sram_mem[69425] = 16'b0000000000000000;
	sram_mem[69426] = 16'b0000000000000000;
	sram_mem[69427] = 16'b0000000000000000;
	sram_mem[69428] = 16'b0000000000000000;
	sram_mem[69429] = 16'b0000000000000000;
	sram_mem[69430] = 16'b0000000000000000;
	sram_mem[69431] = 16'b0000000000000000;
	sram_mem[69432] = 16'b0000000000000000;
	sram_mem[69433] = 16'b0000000000000000;
	sram_mem[69434] = 16'b0000000000000000;
	sram_mem[69435] = 16'b0000000000000000;
	sram_mem[69436] = 16'b0000000000000000;
	sram_mem[69437] = 16'b0000000000000000;
	sram_mem[69438] = 16'b0000000000000000;
	sram_mem[69439] = 16'b0000000000000000;
	sram_mem[69440] = 16'b0000000000000000;
	sram_mem[69441] = 16'b0000000000000000;
	sram_mem[69442] = 16'b0000000000000000;
	sram_mem[69443] = 16'b0000000000000000;
	sram_mem[69444] = 16'b0000000000000000;
	sram_mem[69445] = 16'b0000000000000000;
	sram_mem[69446] = 16'b0000000000000000;
	sram_mem[69447] = 16'b0000000000000000;
	sram_mem[69448] = 16'b0000000000000000;
	sram_mem[69449] = 16'b0000000000000000;
	sram_mem[69450] = 16'b0000000000000000;
	sram_mem[69451] = 16'b0000000000000000;
	sram_mem[69452] = 16'b0000000000000000;
	sram_mem[69453] = 16'b0000000000000000;
	sram_mem[69454] = 16'b0000000000000000;
	sram_mem[69455] = 16'b0000000000000000;
	sram_mem[69456] = 16'b0000000000000000;
	sram_mem[69457] = 16'b0000000000000000;
	sram_mem[69458] = 16'b0000000000000000;
	sram_mem[69459] = 16'b0000000000000000;
	sram_mem[69460] = 16'b0000000000000000;
	sram_mem[69461] = 16'b0000000000000000;
	sram_mem[69462] = 16'b0000000000000000;
	sram_mem[69463] = 16'b0000000000000000;
	sram_mem[69464] = 16'b0000000000000000;
	sram_mem[69465] = 16'b0000000000000000;
	sram_mem[69466] = 16'b0000000000000000;
	sram_mem[69467] = 16'b0000000000000000;
	sram_mem[69468] = 16'b0000000000000000;
	sram_mem[69469] = 16'b0000000000000000;
	sram_mem[69470] = 16'b0000000000000000;
	sram_mem[69471] = 16'b0000000000000000;
	sram_mem[69472] = 16'b0000000000000000;
	sram_mem[69473] = 16'b0000000000000000;
	sram_mem[69474] = 16'b0000000000000000;
	sram_mem[69475] = 16'b0000000000000000;
	sram_mem[69476] = 16'b0000000000000000;
	sram_mem[69477] = 16'b0000000000000000;
	sram_mem[69478] = 16'b0000000000000000;
	sram_mem[69479] = 16'b0000000000000000;
	sram_mem[69480] = 16'b0000000000000000;
	sram_mem[69481] = 16'b0000000000000000;
	sram_mem[69482] = 16'b0000000000000000;
	sram_mem[69483] = 16'b0000000000000000;
	sram_mem[69484] = 16'b0000000000000000;
	sram_mem[69485] = 16'b0000000000000000;
	sram_mem[69486] = 16'b0000000000000000;
	sram_mem[69487] = 16'b0000000000000000;
	sram_mem[69488] = 16'b0000000000000000;
	sram_mem[69489] = 16'b0000000000000000;
	sram_mem[69490] = 16'b0000000000000000;
	sram_mem[69491] = 16'b0000000000000000;
	sram_mem[69492] = 16'b0000000000000000;
	sram_mem[69493] = 16'b0000000000000000;
	sram_mem[69494] = 16'b0000000000000000;
	sram_mem[69495] = 16'b0000000000000000;
	sram_mem[69496] = 16'b0000000000000000;
	sram_mem[69497] = 16'b0000000000000000;
	sram_mem[69498] = 16'b0000000000000000;
	sram_mem[69499] = 16'b0000000000000000;
	sram_mem[69500] = 16'b0000000000000000;
	sram_mem[69501] = 16'b0000000000000000;
	sram_mem[69502] = 16'b0000000000000000;
	sram_mem[69503] = 16'b0000000000000000;
	sram_mem[69504] = 16'b0000000000000000;
	sram_mem[69505] = 16'b0000000000000000;
	sram_mem[69506] = 16'b0000000000000000;
	sram_mem[69507] = 16'b0000000000000000;
	sram_mem[69508] = 16'b0000000000000000;
	sram_mem[69509] = 16'b0000000000000000;
	sram_mem[69510] = 16'b0000000000000000;
	sram_mem[69511] = 16'b0000000000000000;
	sram_mem[69512] = 16'b0000000000000000;
	sram_mem[69513] = 16'b0000000000000000;
	sram_mem[69514] = 16'b0000000000000000;
	sram_mem[69515] = 16'b0000000000000000;
	sram_mem[69516] = 16'b0000000000000000;
	sram_mem[69517] = 16'b0000000000000000;
	sram_mem[69518] = 16'b0000000000000000;
	sram_mem[69519] = 16'b0000000000000000;
	sram_mem[69520] = 16'b0000000000000000;
	sram_mem[69521] = 16'b0000000000000000;
	sram_mem[69522] = 16'b0000000000000000;
	sram_mem[69523] = 16'b0000000000000000;
	sram_mem[69524] = 16'b0000000000000000;
	sram_mem[69525] = 16'b0000000000000000;
	sram_mem[69526] = 16'b0000000000000000;
	sram_mem[69527] = 16'b0000000000000000;
	sram_mem[69528] = 16'b0000000000000000;
	sram_mem[69529] = 16'b0000000000000000;
	sram_mem[69530] = 16'b0000000000000000;
	sram_mem[69531] = 16'b0000000000000000;
	sram_mem[69532] = 16'b0000000000000000;
	sram_mem[69533] = 16'b0000000000000000;
	sram_mem[69534] = 16'b0000000000000000;
	sram_mem[69535] = 16'b0000000000000000;
	sram_mem[69536] = 16'b0000000000000000;
	sram_mem[69537] = 16'b0000000000000000;
	sram_mem[69538] = 16'b0000000000000000;
	sram_mem[69539] = 16'b0000000000000000;
	sram_mem[69540] = 16'b0000000000000000;
	sram_mem[69541] = 16'b0000000000000000;
	sram_mem[69542] = 16'b0000000000000000;
	sram_mem[69543] = 16'b0000000000000000;
	sram_mem[69544] = 16'b0000000000000000;
	sram_mem[69545] = 16'b0000000000000000;
	sram_mem[69546] = 16'b0000000000000000;
	sram_mem[69547] = 16'b0000000000000000;
	sram_mem[69548] = 16'b0000000000000000;
	sram_mem[69549] = 16'b0000000000000000;
	sram_mem[69550] = 16'b0000000000000000;
	sram_mem[69551] = 16'b0000000000000000;
	sram_mem[69552] = 16'b0000000000000000;
	sram_mem[69553] = 16'b0000000000000000;
	sram_mem[69554] = 16'b0000000000000000;
	sram_mem[69555] = 16'b0000000000000000;
	sram_mem[69556] = 16'b0000000000000000;
	sram_mem[69557] = 16'b0000000000000000;
	sram_mem[69558] = 16'b0000000000000000;
	sram_mem[69559] = 16'b0000000000000000;
	sram_mem[69560] = 16'b0000000000000000;
	sram_mem[69561] = 16'b0000000000000000;
	sram_mem[69562] = 16'b0000000000000000;
	sram_mem[69563] = 16'b0000000000000000;
	sram_mem[69564] = 16'b0000000000000000;
	sram_mem[69565] = 16'b0000000000000000;
	sram_mem[69566] = 16'b0000000000000000;
	sram_mem[69567] = 16'b0000000000000000;
	sram_mem[69568] = 16'b0000000000000000;
	sram_mem[69569] = 16'b0000000000000000;
	sram_mem[69570] = 16'b0000000000000000;
	sram_mem[69571] = 16'b0000000000000000;
	sram_mem[69572] = 16'b0000000000000000;
	sram_mem[69573] = 16'b0000000000000000;
	sram_mem[69574] = 16'b0000000000000000;
	sram_mem[69575] = 16'b0000000000000000;
	sram_mem[69576] = 16'b0000000000000000;
	sram_mem[69577] = 16'b0000000000000000;
	sram_mem[69578] = 16'b0000000000000000;
	sram_mem[69579] = 16'b0000000000000000;
	sram_mem[69580] = 16'b0000000000000000;
	sram_mem[69581] = 16'b0000000000000000;
	sram_mem[69582] = 16'b0000000000000000;
	sram_mem[69583] = 16'b0000000000000000;
	sram_mem[69584] = 16'b0000000000000000;
	sram_mem[69585] = 16'b0000000000000000;
	sram_mem[69586] = 16'b0000000000000000;
	sram_mem[69587] = 16'b0000000000000000;
	sram_mem[69588] = 16'b0000000000000000;
	sram_mem[69589] = 16'b0000000000000000;
	sram_mem[69590] = 16'b0000000000000000;
	sram_mem[69591] = 16'b0000000000000000;
	sram_mem[69592] = 16'b0000000000000000;
	sram_mem[69593] = 16'b0000000000000000;
	sram_mem[69594] = 16'b0000000000000000;
	sram_mem[69595] = 16'b0000000000000000;
	sram_mem[69596] = 16'b0000000000000000;
	sram_mem[69597] = 16'b0000000000000000;
	sram_mem[69598] = 16'b0000000000000000;
	sram_mem[69599] = 16'b0000000000000000;
	sram_mem[69600] = 16'b0000000000000000;
	sram_mem[69601] = 16'b0000000000000000;
	sram_mem[69602] = 16'b0000000000000000;
	sram_mem[69603] = 16'b0000000000000000;
	sram_mem[69604] = 16'b0000000000000000;
	sram_mem[69605] = 16'b0000000000000000;
	sram_mem[69606] = 16'b0000000000000000;
	sram_mem[69607] = 16'b0000000000000000;
	sram_mem[69608] = 16'b0000000000000000;
	sram_mem[69609] = 16'b0000000000000000;
	sram_mem[69610] = 16'b0000000000000000;
	sram_mem[69611] = 16'b0000000000000000;
	sram_mem[69612] = 16'b0000000000000000;
	sram_mem[69613] = 16'b0000000000000000;
	sram_mem[69614] = 16'b0000000000000000;
	sram_mem[69615] = 16'b0000000000000000;
	sram_mem[69616] = 16'b0000000000000000;
	sram_mem[69617] = 16'b0000000000000000;
	sram_mem[69618] = 16'b0000000000000000;
	sram_mem[69619] = 16'b0000000000000000;
	sram_mem[69620] = 16'b0000000000000000;
	sram_mem[69621] = 16'b0000000000000000;
	sram_mem[69622] = 16'b0000000000000000;
	sram_mem[69623] = 16'b0000000000000000;
	sram_mem[69624] = 16'b0000000000000000;
	sram_mem[69625] = 16'b0000000000000000;
	sram_mem[69626] = 16'b0000000000000000;
	sram_mem[69627] = 16'b0000000000000000;
	sram_mem[69628] = 16'b0000000000000000;
	sram_mem[69629] = 16'b0000000000000000;
	sram_mem[69630] = 16'b0000000000000000;
	sram_mem[69631] = 16'b0000000000000000;
	sram_mem[69632] = 16'b0000000000000000;
	sram_mem[69633] = 16'b0000000000000000;
	sram_mem[69634] = 16'b0000000000000000;
	sram_mem[69635] = 16'b0000000000000000;
	sram_mem[69636] = 16'b0000000000000000;
	sram_mem[69637] = 16'b0000000000000000;
	sram_mem[69638] = 16'b0000000000000000;
	sram_mem[69639] = 16'b0000000000000000;
	sram_mem[69640] = 16'b0000000000000000;
	sram_mem[69641] = 16'b0000000000000000;
	sram_mem[69642] = 16'b0000000000000000;
	sram_mem[69643] = 16'b0000000000000000;
	sram_mem[69644] = 16'b0000000000000000;
	sram_mem[69645] = 16'b0000000000000000;
	sram_mem[69646] = 16'b0000000000000000;
	sram_mem[69647] = 16'b0000000000000000;
	sram_mem[69648] = 16'b0000000000000000;
	sram_mem[69649] = 16'b0000000000000000;
	sram_mem[69650] = 16'b0000000000000000;
	sram_mem[69651] = 16'b0000000000000000;
	sram_mem[69652] = 16'b0000000000000000;
	sram_mem[69653] = 16'b0000000000000000;
	sram_mem[69654] = 16'b0000000000000000;
	sram_mem[69655] = 16'b0000000000000000;
	sram_mem[69656] = 16'b0000000000000000;
	sram_mem[69657] = 16'b0000000000000000;
	sram_mem[69658] = 16'b0000000000000000;
	sram_mem[69659] = 16'b0000000000000000;
	sram_mem[69660] = 16'b0000000000000000;
	sram_mem[69661] = 16'b0000000000000000;
	sram_mem[69662] = 16'b0000000000000000;
	sram_mem[69663] = 16'b0000000000000000;
	sram_mem[69664] = 16'b0000000000000000;
	sram_mem[69665] = 16'b0000000000000000;
	sram_mem[69666] = 16'b0000000000000000;
	sram_mem[69667] = 16'b0000000000000000;
	sram_mem[69668] = 16'b0000000000000000;
	sram_mem[69669] = 16'b0000000000000000;
	sram_mem[69670] = 16'b0000000000000000;
	sram_mem[69671] = 16'b0000000000000000;
	sram_mem[69672] = 16'b0000000000000000;
	sram_mem[69673] = 16'b0000000000000000;
	sram_mem[69674] = 16'b0000000000000000;
	sram_mem[69675] = 16'b0000000000000000;
	sram_mem[69676] = 16'b0000000000000000;
	sram_mem[69677] = 16'b0000000000000000;
	sram_mem[69678] = 16'b0000000000000000;
	sram_mem[69679] = 16'b0000000000000000;
	sram_mem[69680] = 16'b0000000000000000;
	sram_mem[69681] = 16'b0000000000000000;
	sram_mem[69682] = 16'b0000000000000000;
	sram_mem[69683] = 16'b0000000000000000;
	sram_mem[69684] = 16'b0000000000000000;
	sram_mem[69685] = 16'b0000000000000000;
	sram_mem[69686] = 16'b0000000000000000;
	sram_mem[69687] = 16'b0000000000000000;
	sram_mem[69688] = 16'b0000000000000000;
	sram_mem[69689] = 16'b0000000000000000;
	sram_mem[69690] = 16'b0000000000000000;
	sram_mem[69691] = 16'b0000000000000000;
	sram_mem[69692] = 16'b0000000000000000;
	sram_mem[69693] = 16'b0000000000000000;
	sram_mem[69694] = 16'b0000000000000000;
	sram_mem[69695] = 16'b0000000000000000;
	sram_mem[69696] = 16'b0000000000000000;
	sram_mem[69697] = 16'b0000000000000000;
	sram_mem[69698] = 16'b0000000000000000;
	sram_mem[69699] = 16'b0000000000000000;
	sram_mem[69700] = 16'b0000000000000000;
	sram_mem[69701] = 16'b0000000000000000;
	sram_mem[69702] = 16'b0000000000000000;
	sram_mem[69703] = 16'b0000000000000000;
	sram_mem[69704] = 16'b0000000000000000;
	sram_mem[69705] = 16'b0000000000000000;
	sram_mem[69706] = 16'b0000000000000000;
	sram_mem[69707] = 16'b0000000000000000;
	sram_mem[69708] = 16'b0000000000000000;
	sram_mem[69709] = 16'b0000000000000000;
	sram_mem[69710] = 16'b0000000000000000;
	sram_mem[69711] = 16'b0000000000000000;
	sram_mem[69712] = 16'b0000000000000000;
	sram_mem[69713] = 16'b0000000000000000;
	sram_mem[69714] = 16'b0000000000000000;
	sram_mem[69715] = 16'b0000000000000000;
	sram_mem[69716] = 16'b0000000000000000;
	sram_mem[69717] = 16'b0000000000000000;
	sram_mem[69718] = 16'b0000000000000000;
	sram_mem[69719] = 16'b0000000000000000;
	sram_mem[69720] = 16'b0000000000000000;
	sram_mem[69721] = 16'b0000000000000000;
	sram_mem[69722] = 16'b0000000000000000;
	sram_mem[69723] = 16'b0000000000000000;
	sram_mem[69724] = 16'b0000000000000000;
	sram_mem[69725] = 16'b0000000000000000;
	sram_mem[69726] = 16'b0000000000000000;
	sram_mem[69727] = 16'b0000000000000000;
	sram_mem[69728] = 16'b0000000000000000;
	sram_mem[69729] = 16'b0000000000000000;
	sram_mem[69730] = 16'b0000000000000000;
	sram_mem[69731] = 16'b0000000000000000;
	sram_mem[69732] = 16'b0000000000000000;
	sram_mem[69733] = 16'b0000000000000000;
	sram_mem[69734] = 16'b0000000000000000;
	sram_mem[69735] = 16'b0000000000000000;
	sram_mem[69736] = 16'b0000000000000000;
	sram_mem[69737] = 16'b0000000000000000;
	sram_mem[69738] = 16'b0000000000000000;
	sram_mem[69739] = 16'b0000000000000000;
	sram_mem[69740] = 16'b0000000000000000;
	sram_mem[69741] = 16'b0000000000000000;
	sram_mem[69742] = 16'b0000000000000000;
	sram_mem[69743] = 16'b0000000000000000;
	sram_mem[69744] = 16'b0000000000000000;
	sram_mem[69745] = 16'b0000000000000000;
	sram_mem[69746] = 16'b0000000000000000;
	sram_mem[69747] = 16'b0000000000000000;
	sram_mem[69748] = 16'b0000000000000000;
	sram_mem[69749] = 16'b0000000000000000;
	sram_mem[69750] = 16'b0000000000000000;
	sram_mem[69751] = 16'b0000000000000000;
	sram_mem[69752] = 16'b0000000000000000;
	sram_mem[69753] = 16'b0000000000000000;
	sram_mem[69754] = 16'b0000000000000000;
	sram_mem[69755] = 16'b0000000000000000;
	sram_mem[69756] = 16'b0000000000000000;
	sram_mem[69757] = 16'b0000000000000000;
	sram_mem[69758] = 16'b0000000000000000;
	sram_mem[69759] = 16'b0000000000000000;
	sram_mem[69760] = 16'b0000000000000000;
	sram_mem[69761] = 16'b0000000000000000;
	sram_mem[69762] = 16'b0000000000000000;
	sram_mem[69763] = 16'b0000000000000000;
	sram_mem[69764] = 16'b0000000000000000;
	sram_mem[69765] = 16'b0000000000000000;
	sram_mem[69766] = 16'b0000000000000000;
	sram_mem[69767] = 16'b0000000000000000;
	sram_mem[69768] = 16'b0000000000000000;
	sram_mem[69769] = 16'b0000000000000000;
	sram_mem[69770] = 16'b0000000000000000;
	sram_mem[69771] = 16'b0000000000000000;
	sram_mem[69772] = 16'b0000000000000000;
	sram_mem[69773] = 16'b0000000000000000;
	sram_mem[69774] = 16'b0000000000000000;
	sram_mem[69775] = 16'b0000000000000000;
	sram_mem[69776] = 16'b0000000000000000;
	sram_mem[69777] = 16'b0000000000000000;
	sram_mem[69778] = 16'b0000000000000000;
	sram_mem[69779] = 16'b0000000000000000;
	sram_mem[69780] = 16'b0000000000000000;
	sram_mem[69781] = 16'b0000000000000000;
	sram_mem[69782] = 16'b0000000000000000;
	sram_mem[69783] = 16'b0000000000000000;
	sram_mem[69784] = 16'b0000000000000000;
	sram_mem[69785] = 16'b0000000000000000;
	sram_mem[69786] = 16'b0000000000000000;
	sram_mem[69787] = 16'b0000000000000000;
	sram_mem[69788] = 16'b0000000000000000;
	sram_mem[69789] = 16'b0000000000000000;
	sram_mem[69790] = 16'b0000000000000000;
	sram_mem[69791] = 16'b0000000000000000;
	sram_mem[69792] = 16'b0000000000000000;
	sram_mem[69793] = 16'b0000000000000000;
	sram_mem[69794] = 16'b0000000000000000;
	sram_mem[69795] = 16'b0000000000000000;
	sram_mem[69796] = 16'b0000000000000000;
	sram_mem[69797] = 16'b0000000000000000;
	sram_mem[69798] = 16'b0000000000000000;
	sram_mem[69799] = 16'b0000000000000000;
	sram_mem[69800] = 16'b0000000000000000;
	sram_mem[69801] = 16'b0000000000000000;
	sram_mem[69802] = 16'b0000000000000000;
	sram_mem[69803] = 16'b0000000000000000;
	sram_mem[69804] = 16'b0000000000000000;
	sram_mem[69805] = 16'b0000000000000000;
	sram_mem[69806] = 16'b0000000000000000;
	sram_mem[69807] = 16'b0000000000000000;
	sram_mem[69808] = 16'b0000000000000000;
	sram_mem[69809] = 16'b0000000000000000;
	sram_mem[69810] = 16'b0000000000000000;
	sram_mem[69811] = 16'b0000000000000000;
	sram_mem[69812] = 16'b0000000000000000;
	sram_mem[69813] = 16'b0000000000000000;
	sram_mem[69814] = 16'b0000000000000000;
	sram_mem[69815] = 16'b0000000000000000;
	sram_mem[69816] = 16'b0000000000000000;
	sram_mem[69817] = 16'b0000000000000000;
	sram_mem[69818] = 16'b0000000000000000;
	sram_mem[69819] = 16'b0000000000000000;
	sram_mem[69820] = 16'b0000000000000000;
	sram_mem[69821] = 16'b0000000000000000;
	sram_mem[69822] = 16'b0000000000000000;
	sram_mem[69823] = 16'b0000000000000000;
	sram_mem[69824] = 16'b0000000000000000;
	sram_mem[69825] = 16'b0000000000000000;
	sram_mem[69826] = 16'b0000000000000000;
	sram_mem[69827] = 16'b0000000000000000;
	sram_mem[69828] = 16'b0000000000000000;
	sram_mem[69829] = 16'b0000000000000000;
	sram_mem[69830] = 16'b0000000000000000;
	sram_mem[69831] = 16'b0000000000000000;
	sram_mem[69832] = 16'b0000000000000000;
	sram_mem[69833] = 16'b0000000000000000;
	sram_mem[69834] = 16'b0000000000000000;
	sram_mem[69835] = 16'b0000000000000000;
	sram_mem[69836] = 16'b0000000000000000;
	sram_mem[69837] = 16'b0000000000000000;
	sram_mem[69838] = 16'b0000000000000000;
	sram_mem[69839] = 16'b0000000000000000;
	sram_mem[69840] = 16'b0000000000000000;
	sram_mem[69841] = 16'b0000000000000000;
	sram_mem[69842] = 16'b0000000000000000;
	sram_mem[69843] = 16'b0000000000000000;
	sram_mem[69844] = 16'b0000000000000000;
	sram_mem[69845] = 16'b0000000000000000;
	sram_mem[69846] = 16'b0000000000000000;
	sram_mem[69847] = 16'b0000000000000000;
	sram_mem[69848] = 16'b0000000000000000;
	sram_mem[69849] = 16'b0000000000000000;
	sram_mem[69850] = 16'b0000000000000000;
	sram_mem[69851] = 16'b0000000000000000;
	sram_mem[69852] = 16'b0000000000000000;
	sram_mem[69853] = 16'b0000000000000000;
	sram_mem[69854] = 16'b0000000000000000;
	sram_mem[69855] = 16'b0000000000000000;
	sram_mem[69856] = 16'b0000000000000000;
	sram_mem[69857] = 16'b0000000000000000;
	sram_mem[69858] = 16'b0000000000000000;
	sram_mem[69859] = 16'b0000000000000000;
	sram_mem[69860] = 16'b0000000000000000;
	sram_mem[69861] = 16'b0000000000000000;
	sram_mem[69862] = 16'b0000000000000000;
	sram_mem[69863] = 16'b0000000000000000;
	sram_mem[69864] = 16'b0000000000000000;
	sram_mem[69865] = 16'b0000000000000000;
	sram_mem[69866] = 16'b0000000000000000;
	sram_mem[69867] = 16'b0000000000000000;
	sram_mem[69868] = 16'b0000000000000000;
	sram_mem[69869] = 16'b0000000000000000;
	sram_mem[69870] = 16'b0000000000000000;
	sram_mem[69871] = 16'b0000000000000000;
	sram_mem[69872] = 16'b0000000000000000;
	sram_mem[69873] = 16'b0000000000000000;
	sram_mem[69874] = 16'b0000000000000000;
	sram_mem[69875] = 16'b0000000000000000;
	sram_mem[69876] = 16'b0000000000000000;
	sram_mem[69877] = 16'b0000000000000000;
	sram_mem[69878] = 16'b0000000000000000;
	sram_mem[69879] = 16'b0000000000000000;
	sram_mem[69880] = 16'b0000000000000000;
	sram_mem[69881] = 16'b0000000000000000;
	sram_mem[69882] = 16'b0000000000000000;
	sram_mem[69883] = 16'b0000000000000000;
	sram_mem[69884] = 16'b0000000000000000;
	sram_mem[69885] = 16'b0000000000000000;
	sram_mem[69886] = 16'b0000000000000000;
	sram_mem[69887] = 16'b0000000000000000;
	sram_mem[69888] = 16'b0000000000000000;
	sram_mem[69889] = 16'b0000000000000000;
	sram_mem[69890] = 16'b0000000000000000;
	sram_mem[69891] = 16'b0000000000000000;
	sram_mem[69892] = 16'b0000000000000000;
	sram_mem[69893] = 16'b0000000000000000;
	sram_mem[69894] = 16'b0000000000000000;
	sram_mem[69895] = 16'b0000000000000000;
	sram_mem[69896] = 16'b0000000000000000;
	sram_mem[69897] = 16'b0000000000000000;
	sram_mem[69898] = 16'b0000000000000000;
	sram_mem[69899] = 16'b0000000000000000;
	sram_mem[69900] = 16'b0000000000000000;
	sram_mem[69901] = 16'b0000000000000000;
	sram_mem[69902] = 16'b0000000000000000;
	sram_mem[69903] = 16'b0000000000000000;
	sram_mem[69904] = 16'b0000000000000000;
	sram_mem[69905] = 16'b0000000000000000;
	sram_mem[69906] = 16'b0000000000000000;
	sram_mem[69907] = 16'b0000000000000000;
	sram_mem[69908] = 16'b0000000000000000;
	sram_mem[69909] = 16'b0000000000000000;
	sram_mem[69910] = 16'b0000000000000000;
	sram_mem[69911] = 16'b0000000000000000;
	sram_mem[69912] = 16'b0000000000000000;
	sram_mem[69913] = 16'b0000000000000000;
	sram_mem[69914] = 16'b0000000000000000;
	sram_mem[69915] = 16'b0000000000000000;
	sram_mem[69916] = 16'b0000000000000000;
	sram_mem[69917] = 16'b0000000000000000;
	sram_mem[69918] = 16'b0000000000000000;
	sram_mem[69919] = 16'b0000000000000000;
	sram_mem[69920] = 16'b0000000000000000;
	sram_mem[69921] = 16'b0000000000000000;
	sram_mem[69922] = 16'b0000000000000000;
	sram_mem[69923] = 16'b0000000000000000;
	sram_mem[69924] = 16'b0000000000000000;
	sram_mem[69925] = 16'b0000000000000000;
	sram_mem[69926] = 16'b0000000000000000;
	sram_mem[69927] = 16'b0000000000000000;
	sram_mem[69928] = 16'b0000000000000000;
	sram_mem[69929] = 16'b0000000000000000;
	sram_mem[69930] = 16'b0000000000000000;
	sram_mem[69931] = 16'b0000000000000000;
	sram_mem[69932] = 16'b0000000000000000;
	sram_mem[69933] = 16'b0000000000000000;
	sram_mem[69934] = 16'b0000000000000000;
	sram_mem[69935] = 16'b0000000000000000;
	sram_mem[69936] = 16'b0000000000000000;
	sram_mem[69937] = 16'b0000000000000000;
	sram_mem[69938] = 16'b0000000000000000;
	sram_mem[69939] = 16'b0000000000000000;
	sram_mem[69940] = 16'b0000000000000000;
	sram_mem[69941] = 16'b0000000000000000;
	sram_mem[69942] = 16'b0000000000000000;
	sram_mem[69943] = 16'b0000000000000000;
	sram_mem[69944] = 16'b0000000000000000;
	sram_mem[69945] = 16'b0000000000000000;
	sram_mem[69946] = 16'b0000000000000000;
	sram_mem[69947] = 16'b0000000000000000;
	sram_mem[69948] = 16'b0000000000000000;
	sram_mem[69949] = 16'b0000000000000000;
	sram_mem[69950] = 16'b0000000000000000;
	sram_mem[69951] = 16'b0000000000000000;
	sram_mem[69952] = 16'b0000000000000000;
	sram_mem[69953] = 16'b0000000000000000;
	sram_mem[69954] = 16'b0000000000000000;
	sram_mem[69955] = 16'b0000000000000000;
	sram_mem[69956] = 16'b0000000000000000;
	sram_mem[69957] = 16'b0000000000000000;
	sram_mem[69958] = 16'b0000000000000000;
	sram_mem[69959] = 16'b0000000000000000;
	sram_mem[69960] = 16'b0000000000000000;
	sram_mem[69961] = 16'b0000000000000000;
	sram_mem[69962] = 16'b0000000000000000;
	sram_mem[69963] = 16'b0000000000000000;
	sram_mem[69964] = 16'b0000000000000000;
	sram_mem[69965] = 16'b0000000000000000;
	sram_mem[69966] = 16'b0000000000000000;
	sram_mem[69967] = 16'b0000000000000000;
	sram_mem[69968] = 16'b0000000000000000;
	sram_mem[69969] = 16'b0000000000000000;
	sram_mem[69970] = 16'b0000000000000000;
	sram_mem[69971] = 16'b0000000000000000;
	sram_mem[69972] = 16'b0000000000000000;
	sram_mem[69973] = 16'b0000000000000000;
	sram_mem[69974] = 16'b0000000000000000;
	sram_mem[69975] = 16'b0000000000000000;
	sram_mem[69976] = 16'b0000000000000000;
	sram_mem[69977] = 16'b0000000000000000;
	sram_mem[69978] = 16'b0000000000000000;
	sram_mem[69979] = 16'b0000000000000000;
	sram_mem[69980] = 16'b0000000000000000;
	sram_mem[69981] = 16'b0000000000000000;
	sram_mem[69982] = 16'b0000000000000000;
	sram_mem[69983] = 16'b0000000000000000;
	sram_mem[69984] = 16'b0000000000000000;
	sram_mem[69985] = 16'b0000000000000000;
	sram_mem[69986] = 16'b0000000000000000;
	sram_mem[69987] = 16'b0000000000000000;
	sram_mem[69988] = 16'b0000000000000000;
	sram_mem[69989] = 16'b0000000000000000;
	sram_mem[69990] = 16'b0000000000000000;
	sram_mem[69991] = 16'b0000000000000000;
	sram_mem[69992] = 16'b0000000000000000;
	sram_mem[69993] = 16'b0000000000000000;
	sram_mem[69994] = 16'b0000000000000000;
	sram_mem[69995] = 16'b0000000000000000;
	sram_mem[69996] = 16'b0000000000000000;
	sram_mem[69997] = 16'b0000000000000000;
	sram_mem[69998] = 16'b0000000000000000;
	sram_mem[69999] = 16'b0000000000000000;
	sram_mem[70000] = 16'b0000000000000000;
	sram_mem[70001] = 16'b0000000000000000;
	sram_mem[70002] = 16'b0000000000000000;
	sram_mem[70003] = 16'b0000000000000000;
	sram_mem[70004] = 16'b0000000000000000;
	sram_mem[70005] = 16'b0000000000000000;
	sram_mem[70006] = 16'b0000000000000000;
	sram_mem[70007] = 16'b0000000000000000;
	sram_mem[70008] = 16'b0000000000000000;
	sram_mem[70009] = 16'b0000000000000000;
	sram_mem[70010] = 16'b0000000000000000;
	sram_mem[70011] = 16'b0000000000000000;
	sram_mem[70012] = 16'b0000000000000000;
	sram_mem[70013] = 16'b0000000000000000;
	sram_mem[70014] = 16'b0000000000000000;
	sram_mem[70015] = 16'b0000000000000000;
	sram_mem[70016] = 16'b0000000000000000;
	sram_mem[70017] = 16'b0000000000000000;
	sram_mem[70018] = 16'b0000000000000000;
	sram_mem[70019] = 16'b0000000000000000;
	sram_mem[70020] = 16'b0000000000000000;
	sram_mem[70021] = 16'b0000000000000000;
	sram_mem[70022] = 16'b0000000000000000;
	sram_mem[70023] = 16'b0000000000000000;
	sram_mem[70024] = 16'b0000000000000000;
	sram_mem[70025] = 16'b0000000000000000;
	sram_mem[70026] = 16'b0000000000000000;
	sram_mem[70027] = 16'b0000000000000000;
	sram_mem[70028] = 16'b0000000000000000;
	sram_mem[70029] = 16'b0000000000000000;
	sram_mem[70030] = 16'b0000000000000000;
	sram_mem[70031] = 16'b0000000000000000;
	sram_mem[70032] = 16'b0000000000000000;
	sram_mem[70033] = 16'b0000000000000000;
	sram_mem[70034] = 16'b0000000000000000;
	sram_mem[70035] = 16'b0000000000000000;
	sram_mem[70036] = 16'b0000000000000000;
	sram_mem[70037] = 16'b0000000000000000;
	sram_mem[70038] = 16'b0000000000000000;
	sram_mem[70039] = 16'b0000000000000000;
	sram_mem[70040] = 16'b0000000000000000;
	sram_mem[70041] = 16'b0000000000000000;
	sram_mem[70042] = 16'b0000000000000000;
	sram_mem[70043] = 16'b0000000000000000;
	sram_mem[70044] = 16'b0000000000000000;
	sram_mem[70045] = 16'b0000000000000000;
	sram_mem[70046] = 16'b0000000000000000;
	sram_mem[70047] = 16'b0000000000000000;
	sram_mem[70048] = 16'b0000000000000000;
	sram_mem[70049] = 16'b0000000000000000;
	sram_mem[70050] = 16'b0000000000000000;
	sram_mem[70051] = 16'b0000000000000000;
	sram_mem[70052] = 16'b0000000000000000;
	sram_mem[70053] = 16'b0000000000000000;
	sram_mem[70054] = 16'b0000000000000000;
	sram_mem[70055] = 16'b0000000000000000;
	sram_mem[70056] = 16'b0000000000000000;
	sram_mem[70057] = 16'b0000000000000000;
	sram_mem[70058] = 16'b0000000000000000;
	sram_mem[70059] = 16'b0000000000000000;
	sram_mem[70060] = 16'b0000000000000000;
	sram_mem[70061] = 16'b0000000000000000;
	sram_mem[70062] = 16'b0000000000000000;
	sram_mem[70063] = 16'b0000000000000000;
	sram_mem[70064] = 16'b0000000000000000;
	sram_mem[70065] = 16'b0000000000000000;
	sram_mem[70066] = 16'b0000000000000000;
	sram_mem[70067] = 16'b0000000000000000;
	sram_mem[70068] = 16'b0000000000000000;
	sram_mem[70069] = 16'b0000000000000000;
	sram_mem[70070] = 16'b0000000000000000;
	sram_mem[70071] = 16'b0000000000000000;
	sram_mem[70072] = 16'b0000000000000000;
	sram_mem[70073] = 16'b0000000000000000;
	sram_mem[70074] = 16'b0000000000000000;
	sram_mem[70075] = 16'b0000000000000000;
	sram_mem[70076] = 16'b0000000000000000;
	sram_mem[70077] = 16'b0000000000000000;
	sram_mem[70078] = 16'b0000000000000000;
	sram_mem[70079] = 16'b0000000000000000;
	sram_mem[70080] = 16'b0000000000000000;
	sram_mem[70081] = 16'b0000000000000000;
	sram_mem[70082] = 16'b0000000000000000;
	sram_mem[70083] = 16'b0000000000000000;
	sram_mem[70084] = 16'b0000000000000000;
	sram_mem[70085] = 16'b0000000000000000;
	sram_mem[70086] = 16'b0000000000000000;
	sram_mem[70087] = 16'b0000000000000000;
	sram_mem[70088] = 16'b0000000000000000;
	sram_mem[70089] = 16'b0000000000000000;
	sram_mem[70090] = 16'b0000000000000000;
	sram_mem[70091] = 16'b0000000000000000;
	sram_mem[70092] = 16'b0000000000000000;
	sram_mem[70093] = 16'b0000000000000000;
	sram_mem[70094] = 16'b0000000000000000;
	sram_mem[70095] = 16'b0000000000000000;
	sram_mem[70096] = 16'b0000000000000000;
	sram_mem[70097] = 16'b0000000000000000;
	sram_mem[70098] = 16'b0000000000000000;
	sram_mem[70099] = 16'b0000000000000000;
	sram_mem[70100] = 16'b0000000000000000;
	sram_mem[70101] = 16'b0000000000000000;
	sram_mem[70102] = 16'b0000000000000000;
	sram_mem[70103] = 16'b0000000000000000;
	sram_mem[70104] = 16'b0000000000000000;
	sram_mem[70105] = 16'b0000000000000000;
	sram_mem[70106] = 16'b0000000000000000;
	sram_mem[70107] = 16'b0000000000000000;
	sram_mem[70108] = 16'b0000000000000000;
	sram_mem[70109] = 16'b0000000000000000;
	sram_mem[70110] = 16'b0000000000000000;
	sram_mem[70111] = 16'b0000000000000000;
	sram_mem[70112] = 16'b0000000000000000;
	sram_mem[70113] = 16'b0000000000000000;
	sram_mem[70114] = 16'b0000000000000000;
	sram_mem[70115] = 16'b0000000000000000;
	sram_mem[70116] = 16'b0000000000000000;
	sram_mem[70117] = 16'b0000000000000000;
	sram_mem[70118] = 16'b0000000000000000;
	sram_mem[70119] = 16'b0000000000000000;
	sram_mem[70120] = 16'b0000000000000000;
	sram_mem[70121] = 16'b0000000000000000;
	sram_mem[70122] = 16'b0000000000000000;
	sram_mem[70123] = 16'b0000000000000000;
	sram_mem[70124] = 16'b0000000000000000;
	sram_mem[70125] = 16'b0000000000000000;
	sram_mem[70126] = 16'b0000000000000000;
	sram_mem[70127] = 16'b0000000000000000;
	sram_mem[70128] = 16'b0000000000000000;
	sram_mem[70129] = 16'b0000000000000000;
	sram_mem[70130] = 16'b0000000000000000;
	sram_mem[70131] = 16'b0000000000000000;
	sram_mem[70132] = 16'b0000000000000000;
	sram_mem[70133] = 16'b0000000000000000;
	sram_mem[70134] = 16'b0000000000000000;
	sram_mem[70135] = 16'b0000000000000000;
	sram_mem[70136] = 16'b0000000000000000;
	sram_mem[70137] = 16'b0000000000000000;
	sram_mem[70138] = 16'b0000000000000000;
	sram_mem[70139] = 16'b0000000000000000;
	sram_mem[70140] = 16'b0000000000000000;
	sram_mem[70141] = 16'b0000000000000000;
	sram_mem[70142] = 16'b0000000000000000;
	sram_mem[70143] = 16'b0000000000000000;
	sram_mem[70144] = 16'b0000000000000000;
	sram_mem[70145] = 16'b0000000000000000;
	sram_mem[70146] = 16'b0000000000000000;
	sram_mem[70147] = 16'b0000000000000000;
	sram_mem[70148] = 16'b0000000000000000;
	sram_mem[70149] = 16'b0000000000000000;
	sram_mem[70150] = 16'b0000000000000000;
	sram_mem[70151] = 16'b0000000000000000;
	sram_mem[70152] = 16'b0000000000000000;
	sram_mem[70153] = 16'b0000000000000000;
	sram_mem[70154] = 16'b0000000000000000;
	sram_mem[70155] = 16'b0000000000000000;
	sram_mem[70156] = 16'b0000000000000000;
	sram_mem[70157] = 16'b0000000000000000;
	sram_mem[70158] = 16'b0000000000000000;
	sram_mem[70159] = 16'b0000000000000000;
	sram_mem[70160] = 16'b0000000000000000;
	sram_mem[70161] = 16'b0000000000000000;
	sram_mem[70162] = 16'b0000000000000000;
	sram_mem[70163] = 16'b0000000000000000;
	sram_mem[70164] = 16'b0000000000000000;
	sram_mem[70165] = 16'b0000000000000000;
	sram_mem[70166] = 16'b0000000000000000;
	sram_mem[70167] = 16'b0000000000000000;
	sram_mem[70168] = 16'b0000000000000000;
	sram_mem[70169] = 16'b0000000000000000;
	sram_mem[70170] = 16'b0000000000000000;
	sram_mem[70171] = 16'b0000000000000000;
	sram_mem[70172] = 16'b0000000000000000;
	sram_mem[70173] = 16'b0000000000000000;
	sram_mem[70174] = 16'b0000000000000000;
	sram_mem[70175] = 16'b0000000000000000;
	sram_mem[70176] = 16'b0000000000000000;
	sram_mem[70177] = 16'b0000000000000000;
	sram_mem[70178] = 16'b0000000000000000;
	sram_mem[70179] = 16'b0000000000000000;
	sram_mem[70180] = 16'b0000000000000000;
	sram_mem[70181] = 16'b0000000000000000;
	sram_mem[70182] = 16'b0000000000000000;
	sram_mem[70183] = 16'b0000000000000000;
	sram_mem[70184] = 16'b0000000000000000;
	sram_mem[70185] = 16'b0000000000000000;
	sram_mem[70186] = 16'b0000000000000000;
	sram_mem[70187] = 16'b0000000000000000;
	sram_mem[70188] = 16'b0000000000000000;
	sram_mem[70189] = 16'b0000000000000000;
	sram_mem[70190] = 16'b0000000000000000;
	sram_mem[70191] = 16'b0000000000000000;
	sram_mem[70192] = 16'b0000000000000000;
	sram_mem[70193] = 16'b0000000000000000;
	sram_mem[70194] = 16'b0000000000000000;
	sram_mem[70195] = 16'b0000000000000000;
	sram_mem[70196] = 16'b0000000000000000;
	sram_mem[70197] = 16'b0000000000000000;
	sram_mem[70198] = 16'b0000000000000000;
	sram_mem[70199] = 16'b0000000000000000;
	sram_mem[70200] = 16'b0000000000000000;
	sram_mem[70201] = 16'b0000000000000000;
	sram_mem[70202] = 16'b0000000000000000;
	sram_mem[70203] = 16'b0000000000000000;
	sram_mem[70204] = 16'b0000000000000000;
	sram_mem[70205] = 16'b0000000000000000;
	sram_mem[70206] = 16'b0000000000000000;
	sram_mem[70207] = 16'b0000000000000000;
	sram_mem[70208] = 16'b0000000000000000;
	sram_mem[70209] = 16'b0000000000000000;
	sram_mem[70210] = 16'b0000000000000000;
	sram_mem[70211] = 16'b0000000000000000;
	sram_mem[70212] = 16'b0000000000000000;
	sram_mem[70213] = 16'b0000000000000000;
	sram_mem[70214] = 16'b0000000000000000;
	sram_mem[70215] = 16'b0000000000000000;
	sram_mem[70216] = 16'b0000000000000000;
	sram_mem[70217] = 16'b0000000000000000;
	sram_mem[70218] = 16'b0000000000000000;
	sram_mem[70219] = 16'b0000000000000000;
	sram_mem[70220] = 16'b0000000000000000;
	sram_mem[70221] = 16'b0000000000000000;
	sram_mem[70222] = 16'b0000000000000000;
	sram_mem[70223] = 16'b0000000000000000;
	sram_mem[70224] = 16'b0000000000000000;
	sram_mem[70225] = 16'b0000000000000000;
	sram_mem[70226] = 16'b0000000000000000;
	sram_mem[70227] = 16'b0000000000000000;
	sram_mem[70228] = 16'b0000000000000000;
	sram_mem[70229] = 16'b0000000000000000;
	sram_mem[70230] = 16'b0000000000000000;
	sram_mem[70231] = 16'b0000000000000000;
	sram_mem[70232] = 16'b0000000000000000;
	sram_mem[70233] = 16'b0000000000000000;
	sram_mem[70234] = 16'b0000000000000000;
	sram_mem[70235] = 16'b0000000000000000;
	sram_mem[70236] = 16'b0000000000000000;
	sram_mem[70237] = 16'b0000000000000000;
	sram_mem[70238] = 16'b0000000000000000;
	sram_mem[70239] = 16'b0000000000000000;
	sram_mem[70240] = 16'b0000000000000000;
	sram_mem[70241] = 16'b0000000000000000;
	sram_mem[70242] = 16'b0000000000000000;
	sram_mem[70243] = 16'b0000000000000000;
	sram_mem[70244] = 16'b0000000000000000;
	sram_mem[70245] = 16'b0000000000000000;
	sram_mem[70246] = 16'b0000000000000000;
	sram_mem[70247] = 16'b0000000000000000;
	sram_mem[70248] = 16'b0000000000000000;
	sram_mem[70249] = 16'b0000000000000000;
	sram_mem[70250] = 16'b0000000000000000;
	sram_mem[70251] = 16'b0000000000000000;
	sram_mem[70252] = 16'b0000000000000000;
	sram_mem[70253] = 16'b0000000000000000;
	sram_mem[70254] = 16'b0000000000000000;
	sram_mem[70255] = 16'b0000000000000000;
	sram_mem[70256] = 16'b0000000000000000;
	sram_mem[70257] = 16'b0000000000000000;
	sram_mem[70258] = 16'b0000000000000000;
	sram_mem[70259] = 16'b0000000000000000;
	sram_mem[70260] = 16'b0000000000000000;
	sram_mem[70261] = 16'b0000000000000000;
	sram_mem[70262] = 16'b0000000000000000;
	sram_mem[70263] = 16'b0000000000000000;
	sram_mem[70264] = 16'b0000000000000000;
	sram_mem[70265] = 16'b0000000000000000;
	sram_mem[70266] = 16'b0000000000000000;
	sram_mem[70267] = 16'b0000000000000000;
	sram_mem[70268] = 16'b0000000000000000;
	sram_mem[70269] = 16'b0000000000000000;
	sram_mem[70270] = 16'b0000000000000000;
	sram_mem[70271] = 16'b0000000000000000;
	sram_mem[70272] = 16'b0000000000000000;
	sram_mem[70273] = 16'b0000000000000000;
	sram_mem[70274] = 16'b0000000000000000;
	sram_mem[70275] = 16'b0000000000000000;
	sram_mem[70276] = 16'b0000000000000000;
	sram_mem[70277] = 16'b0000000000000000;
	sram_mem[70278] = 16'b0000000000000000;
	sram_mem[70279] = 16'b0000000000000000;
	sram_mem[70280] = 16'b0000000000000000;
	sram_mem[70281] = 16'b0000000000000000;
	sram_mem[70282] = 16'b0000000000000000;
	sram_mem[70283] = 16'b0000000000000000;
	sram_mem[70284] = 16'b0000000000000000;
	sram_mem[70285] = 16'b0000000000000000;
	sram_mem[70286] = 16'b0000000000000000;
	sram_mem[70287] = 16'b0000000000000000;
	sram_mem[70288] = 16'b0000000000000000;
	sram_mem[70289] = 16'b0000000000000000;
	sram_mem[70290] = 16'b0000000000000000;
	sram_mem[70291] = 16'b0000000000000000;
	sram_mem[70292] = 16'b0000000000000000;
	sram_mem[70293] = 16'b0000000000000000;
	sram_mem[70294] = 16'b0000000000000000;
	sram_mem[70295] = 16'b0000000000000000;
	sram_mem[70296] = 16'b0000000000000000;
	sram_mem[70297] = 16'b0000000000000000;
	sram_mem[70298] = 16'b0000000000000000;
	sram_mem[70299] = 16'b0000000000000000;
	sram_mem[70300] = 16'b0000000000000000;
	sram_mem[70301] = 16'b0000000000000000;
	sram_mem[70302] = 16'b0000000000000000;
	sram_mem[70303] = 16'b0000000000000000;
	sram_mem[70304] = 16'b0000000000000000;
	sram_mem[70305] = 16'b0000000000000000;
	sram_mem[70306] = 16'b0000000000000000;
	sram_mem[70307] = 16'b0000000000000000;
	sram_mem[70308] = 16'b0000000000000000;
	sram_mem[70309] = 16'b0000000000000000;
	sram_mem[70310] = 16'b0000000000000000;
	sram_mem[70311] = 16'b0000000000000000;
	sram_mem[70312] = 16'b0000000000000000;
	sram_mem[70313] = 16'b0000000000000000;
	sram_mem[70314] = 16'b0000000000000000;
	sram_mem[70315] = 16'b0000000000000000;
	sram_mem[70316] = 16'b0000000000000000;
	sram_mem[70317] = 16'b0000000000000000;
	sram_mem[70318] = 16'b0000000000000000;
	sram_mem[70319] = 16'b0000000000000000;
	sram_mem[70320] = 16'b0000000000000000;
	sram_mem[70321] = 16'b0000000000000000;
	sram_mem[70322] = 16'b0000000000000000;
	sram_mem[70323] = 16'b0000000000000000;
	sram_mem[70324] = 16'b0000000000000000;
	sram_mem[70325] = 16'b0000000000000000;
	sram_mem[70326] = 16'b0000000000000000;
	sram_mem[70327] = 16'b0000000000000000;
	sram_mem[70328] = 16'b0000000000000000;
	sram_mem[70329] = 16'b0000000000000000;
	sram_mem[70330] = 16'b0000000000000000;
	sram_mem[70331] = 16'b0000000000000000;
	sram_mem[70332] = 16'b0000000000000000;
	sram_mem[70333] = 16'b0000000000000000;
	sram_mem[70334] = 16'b0000000000000000;
	sram_mem[70335] = 16'b0000000000000000;
	sram_mem[70336] = 16'b0000000000000000;
	sram_mem[70337] = 16'b0000000000000000;
	sram_mem[70338] = 16'b0000000000000000;
	sram_mem[70339] = 16'b0000000000000000;
	sram_mem[70340] = 16'b0000000000000000;
	sram_mem[70341] = 16'b0000000000000000;
	sram_mem[70342] = 16'b0000000000000000;
	sram_mem[70343] = 16'b0000000000000000;
	sram_mem[70344] = 16'b0000000000000000;
	sram_mem[70345] = 16'b0000000000000000;
	sram_mem[70346] = 16'b0000000000000000;
	sram_mem[70347] = 16'b0000000000000000;
	sram_mem[70348] = 16'b0000000000000000;
	sram_mem[70349] = 16'b0000000000000000;
	sram_mem[70350] = 16'b0000000000000000;
	sram_mem[70351] = 16'b0000000000000000;
	sram_mem[70352] = 16'b0000000000000000;
	sram_mem[70353] = 16'b0000000000000000;
	sram_mem[70354] = 16'b0000000000000000;
	sram_mem[70355] = 16'b0000000000000000;
	sram_mem[70356] = 16'b0000000000000000;
	sram_mem[70357] = 16'b0000000000000000;
	sram_mem[70358] = 16'b0000000000000000;
	sram_mem[70359] = 16'b0000000000000000;
	sram_mem[70360] = 16'b0000000000000000;
	sram_mem[70361] = 16'b0000000000000000;
	sram_mem[70362] = 16'b0000000000000000;
	sram_mem[70363] = 16'b0000000000000000;
	sram_mem[70364] = 16'b0000000000000000;
	sram_mem[70365] = 16'b0000000000000000;
	sram_mem[70366] = 16'b0000000000000000;
	sram_mem[70367] = 16'b0000000000000000;
	sram_mem[70368] = 16'b0000000000000000;
	sram_mem[70369] = 16'b0000000000000000;
	sram_mem[70370] = 16'b0000000000000000;
	sram_mem[70371] = 16'b0000000000000000;
	sram_mem[70372] = 16'b0000000000000000;
	sram_mem[70373] = 16'b0000000000000000;
	sram_mem[70374] = 16'b0000000000000000;
	sram_mem[70375] = 16'b0000000000000000;
	sram_mem[70376] = 16'b0000000000000000;
	sram_mem[70377] = 16'b0000000000000000;
	sram_mem[70378] = 16'b0000000000000000;
	sram_mem[70379] = 16'b0000000000000000;
	sram_mem[70380] = 16'b0000000000000000;
	sram_mem[70381] = 16'b0000000000000000;
	sram_mem[70382] = 16'b0000000000000000;
	sram_mem[70383] = 16'b0000000000000000;
	sram_mem[70384] = 16'b0000000000000000;
	sram_mem[70385] = 16'b0000000000000000;
	sram_mem[70386] = 16'b0000000000000000;
	sram_mem[70387] = 16'b0000000000000000;
	sram_mem[70388] = 16'b0000000000000000;
	sram_mem[70389] = 16'b0000000000000000;
	sram_mem[70390] = 16'b0000000000000000;
	sram_mem[70391] = 16'b0000000000000000;
	sram_mem[70392] = 16'b0000000000000000;
	sram_mem[70393] = 16'b0000000000000000;
	sram_mem[70394] = 16'b0000000000000000;
	sram_mem[70395] = 16'b0000000000000000;
	sram_mem[70396] = 16'b0000000000000000;
	sram_mem[70397] = 16'b0000000000000000;
	sram_mem[70398] = 16'b0000000000000000;
	sram_mem[70399] = 16'b0000000000000000;
	sram_mem[70400] = 16'b0000000000000000;
	sram_mem[70401] = 16'b0000000000000000;
	sram_mem[70402] = 16'b0000000000000000;
	sram_mem[70403] = 16'b0000000000000000;
	sram_mem[70404] = 16'b0000000000000000;
	sram_mem[70405] = 16'b0000000000000000;
	sram_mem[70406] = 16'b0000000000000000;
	sram_mem[70407] = 16'b0000000000000000;
	sram_mem[70408] = 16'b0000000000000000;
	sram_mem[70409] = 16'b0000000000000000;
	sram_mem[70410] = 16'b0000000000000000;
	sram_mem[70411] = 16'b0000000000000000;
	sram_mem[70412] = 16'b0000000000000000;
	sram_mem[70413] = 16'b0000000000000000;
	sram_mem[70414] = 16'b0000000000000000;
	sram_mem[70415] = 16'b0000000000000000;
	sram_mem[70416] = 16'b0000000000000000;
	sram_mem[70417] = 16'b0000000000000000;
	sram_mem[70418] = 16'b0000000000000000;
	sram_mem[70419] = 16'b0000000000000000;
	sram_mem[70420] = 16'b0000000000000000;
	sram_mem[70421] = 16'b0000000000000000;
	sram_mem[70422] = 16'b0000000000000000;
	sram_mem[70423] = 16'b0000000000000000;
	sram_mem[70424] = 16'b0000000000000000;
	sram_mem[70425] = 16'b0000000000000000;
	sram_mem[70426] = 16'b0000000000000000;
	sram_mem[70427] = 16'b0000000000000000;
	sram_mem[70428] = 16'b0000000000000000;
	sram_mem[70429] = 16'b0000000000000000;
	sram_mem[70430] = 16'b0000000000000000;
	sram_mem[70431] = 16'b0000000000000000;
	sram_mem[70432] = 16'b0000000000000000;
	sram_mem[70433] = 16'b0000000000000000;
	sram_mem[70434] = 16'b0000000000000000;
	sram_mem[70435] = 16'b0000000000000000;
	sram_mem[70436] = 16'b0000000000000000;
	sram_mem[70437] = 16'b0000000000000000;
	sram_mem[70438] = 16'b0000000000000000;
	sram_mem[70439] = 16'b0000000000000000;
	sram_mem[70440] = 16'b0000000000000000;
	sram_mem[70441] = 16'b0000000000000000;
	sram_mem[70442] = 16'b0000000000000000;
	sram_mem[70443] = 16'b0000000000000000;
	sram_mem[70444] = 16'b0000000000000000;
	sram_mem[70445] = 16'b0000000000000000;
	sram_mem[70446] = 16'b0000000000000000;
	sram_mem[70447] = 16'b0000000000000000;
	sram_mem[70448] = 16'b0000000000000000;
	sram_mem[70449] = 16'b0000000000000000;
	sram_mem[70450] = 16'b0000000000000000;
	sram_mem[70451] = 16'b0000000000000000;
	sram_mem[70452] = 16'b0000000000000000;
	sram_mem[70453] = 16'b0000000000000000;
	sram_mem[70454] = 16'b0000000000000000;
	sram_mem[70455] = 16'b0000000000000000;
	sram_mem[70456] = 16'b0000000000000000;
	sram_mem[70457] = 16'b0000000000000000;
	sram_mem[70458] = 16'b0000000000000000;
	sram_mem[70459] = 16'b0000000000000000;
	sram_mem[70460] = 16'b0000000000000000;
	sram_mem[70461] = 16'b0000000000000000;
	sram_mem[70462] = 16'b0000000000000000;
	sram_mem[70463] = 16'b0000000000000000;
	sram_mem[70464] = 16'b0000000000000000;
	sram_mem[70465] = 16'b0000000000000000;
	sram_mem[70466] = 16'b0000000000000000;
	sram_mem[70467] = 16'b0000000000000000;
	sram_mem[70468] = 16'b0000000000000000;
	sram_mem[70469] = 16'b0000000000000000;
	sram_mem[70470] = 16'b0000000000000000;
	sram_mem[70471] = 16'b0000000000000000;
	sram_mem[70472] = 16'b0000000000000000;
	sram_mem[70473] = 16'b0000000000000000;
	sram_mem[70474] = 16'b0000000000000000;
	sram_mem[70475] = 16'b0000000000000000;
	sram_mem[70476] = 16'b0000000000000000;
	sram_mem[70477] = 16'b0000000000000000;
	sram_mem[70478] = 16'b0000000000000000;
	sram_mem[70479] = 16'b0000000000000000;
	sram_mem[70480] = 16'b0000000000000000;
	sram_mem[70481] = 16'b0000000000000000;
	sram_mem[70482] = 16'b0000000000000000;
	sram_mem[70483] = 16'b0000000000000000;
	sram_mem[70484] = 16'b0000000000000000;
	sram_mem[70485] = 16'b0000000000000000;
	sram_mem[70486] = 16'b0000000000000000;
	sram_mem[70487] = 16'b0000000000000000;
	sram_mem[70488] = 16'b0000000000000000;
	sram_mem[70489] = 16'b0000000000000000;
	sram_mem[70490] = 16'b0000000000000000;
	sram_mem[70491] = 16'b0000000000000000;
	sram_mem[70492] = 16'b0000000000000000;
	sram_mem[70493] = 16'b0000000000000000;
	sram_mem[70494] = 16'b0000000000000000;
	sram_mem[70495] = 16'b0000000000000000;
	sram_mem[70496] = 16'b0000000000000000;
	sram_mem[70497] = 16'b0000000000000000;
	sram_mem[70498] = 16'b0000000000000000;
	sram_mem[70499] = 16'b0000000000000000;
	sram_mem[70500] = 16'b0000000000000000;
	sram_mem[70501] = 16'b0000000000000000;
	sram_mem[70502] = 16'b0000000000000000;
	sram_mem[70503] = 16'b0000000000000000;
	sram_mem[70504] = 16'b0000000000000000;
	sram_mem[70505] = 16'b0000000000000000;
	sram_mem[70506] = 16'b0000000000000000;
	sram_mem[70507] = 16'b0000000000000000;
	sram_mem[70508] = 16'b0000000000000000;
	sram_mem[70509] = 16'b0000000000000000;
	sram_mem[70510] = 16'b0000000000000000;
	sram_mem[70511] = 16'b0000000000000000;
	sram_mem[70512] = 16'b0000000000000000;
	sram_mem[70513] = 16'b0000000000000000;
	sram_mem[70514] = 16'b0000000000000000;
	sram_mem[70515] = 16'b0000000000000000;
	sram_mem[70516] = 16'b0000000000000000;
	sram_mem[70517] = 16'b0000000000000000;
	sram_mem[70518] = 16'b0000000000000000;
	sram_mem[70519] = 16'b0000000000000000;
	sram_mem[70520] = 16'b0000000000000000;
	sram_mem[70521] = 16'b0000000000000000;
	sram_mem[70522] = 16'b0000000000000000;
	sram_mem[70523] = 16'b0000000000000000;
	sram_mem[70524] = 16'b0000000000000000;
	sram_mem[70525] = 16'b0000000000000000;
	sram_mem[70526] = 16'b0000000000000000;
	sram_mem[70527] = 16'b0000000000000000;
	sram_mem[70528] = 16'b0000000000000000;
	sram_mem[70529] = 16'b0000000000000000;
	sram_mem[70530] = 16'b0000000000000000;
	sram_mem[70531] = 16'b0000000000000000;
	sram_mem[70532] = 16'b0000000000000000;
	sram_mem[70533] = 16'b0000000000000000;
	sram_mem[70534] = 16'b0000000000000000;
	sram_mem[70535] = 16'b0000000000000000;
	sram_mem[70536] = 16'b0000000000000000;
	sram_mem[70537] = 16'b0000000000000000;
	sram_mem[70538] = 16'b0000000000000000;
	sram_mem[70539] = 16'b0000000000000000;
	sram_mem[70540] = 16'b0000000000000000;
	sram_mem[70541] = 16'b0000000000000000;
	sram_mem[70542] = 16'b0000000000000000;
	sram_mem[70543] = 16'b0000000000000000;
	sram_mem[70544] = 16'b0000000000000000;
	sram_mem[70545] = 16'b0000000000000000;
	sram_mem[70546] = 16'b0000000000000000;
	sram_mem[70547] = 16'b0000000000000000;
	sram_mem[70548] = 16'b0000000000000000;
	sram_mem[70549] = 16'b0000000000000000;
	sram_mem[70550] = 16'b0000000000000000;
	sram_mem[70551] = 16'b0000000000000000;
	sram_mem[70552] = 16'b0000000000000000;
	sram_mem[70553] = 16'b0000000000000000;
	sram_mem[70554] = 16'b0000000000000000;
	sram_mem[70555] = 16'b0000000000000000;
	sram_mem[70556] = 16'b0000000000000000;
	sram_mem[70557] = 16'b0000000000000000;
	sram_mem[70558] = 16'b0000000000000000;
	sram_mem[70559] = 16'b0000000000000000;
	sram_mem[70560] = 16'b0000000000000000;
	sram_mem[70561] = 16'b0000000000000000;
	sram_mem[70562] = 16'b0000000000000000;
	sram_mem[70563] = 16'b0000000000000000;
	sram_mem[70564] = 16'b0000000000000000;
	sram_mem[70565] = 16'b0000000000000000;
	sram_mem[70566] = 16'b0000000000000000;
	sram_mem[70567] = 16'b0000000000000000;
	sram_mem[70568] = 16'b0000000000000000;
	sram_mem[70569] = 16'b0000000000000000;
	sram_mem[70570] = 16'b0000000000000000;
	sram_mem[70571] = 16'b0000000000000000;
	sram_mem[70572] = 16'b0000000000000000;
	sram_mem[70573] = 16'b0000000000000000;
	sram_mem[70574] = 16'b0000000000000000;
	sram_mem[70575] = 16'b0000000000000000;
	sram_mem[70576] = 16'b0000000000000000;
	sram_mem[70577] = 16'b0000000000000000;
	sram_mem[70578] = 16'b0000000000000000;
	sram_mem[70579] = 16'b0000000000000000;
	sram_mem[70580] = 16'b0000000000000000;
	sram_mem[70581] = 16'b0000000000000000;
	sram_mem[70582] = 16'b0000000000000000;
	sram_mem[70583] = 16'b0000000000000000;
	sram_mem[70584] = 16'b0000000000000000;
	sram_mem[70585] = 16'b0000000000000000;
	sram_mem[70586] = 16'b0000000000000000;
	sram_mem[70587] = 16'b0000000000000000;
	sram_mem[70588] = 16'b0000000000000000;
	sram_mem[70589] = 16'b0000000000000000;
	sram_mem[70590] = 16'b0000000000000000;
	sram_mem[70591] = 16'b0000000000000000;
	sram_mem[70592] = 16'b0000000000000000;
	sram_mem[70593] = 16'b0000000000000000;
	sram_mem[70594] = 16'b0000000000000000;
	sram_mem[70595] = 16'b0000000000000000;
	sram_mem[70596] = 16'b0000000000000000;
	sram_mem[70597] = 16'b0000000000000000;
	sram_mem[70598] = 16'b0000000000000000;
	sram_mem[70599] = 16'b0000000000000000;
	sram_mem[70600] = 16'b0000000000000000;
	sram_mem[70601] = 16'b0000000000000000;
	sram_mem[70602] = 16'b0000000000000000;
	sram_mem[70603] = 16'b0000000000000000;
	sram_mem[70604] = 16'b0000000000000000;
	sram_mem[70605] = 16'b0000000000000000;
	sram_mem[70606] = 16'b0000000000000000;
	sram_mem[70607] = 16'b0000000000000000;
	sram_mem[70608] = 16'b0000000000000000;
	sram_mem[70609] = 16'b0000000000000000;
	sram_mem[70610] = 16'b0000000000000000;
	sram_mem[70611] = 16'b0000000000000000;
	sram_mem[70612] = 16'b0000000000000000;
	sram_mem[70613] = 16'b0000000000000000;
	sram_mem[70614] = 16'b0000000000000000;
	sram_mem[70615] = 16'b0000000000000000;
	sram_mem[70616] = 16'b0000000000000000;
	sram_mem[70617] = 16'b0000000000000000;
	sram_mem[70618] = 16'b0000000000000000;
	sram_mem[70619] = 16'b0000000000000000;
	sram_mem[70620] = 16'b0000000000000000;
	sram_mem[70621] = 16'b0000000000000000;
	sram_mem[70622] = 16'b0000000000000000;
	sram_mem[70623] = 16'b0000000000000000;
	sram_mem[70624] = 16'b0000000000000000;
	sram_mem[70625] = 16'b0000000000000000;
	sram_mem[70626] = 16'b0000000000000000;
	sram_mem[70627] = 16'b0000000000000000;
	sram_mem[70628] = 16'b0000000000000000;
	sram_mem[70629] = 16'b0000000000000000;
	sram_mem[70630] = 16'b0000000000000000;
	sram_mem[70631] = 16'b0000000000000000;
	sram_mem[70632] = 16'b0000000000000000;
	sram_mem[70633] = 16'b0000000000000000;
	sram_mem[70634] = 16'b0000000000000000;
	sram_mem[70635] = 16'b0000000000000000;
	sram_mem[70636] = 16'b0000000000000000;
	sram_mem[70637] = 16'b0000000000000000;
	sram_mem[70638] = 16'b0000000000000000;
	sram_mem[70639] = 16'b0000000000000000;
	sram_mem[70640] = 16'b0000000000000000;
	sram_mem[70641] = 16'b0000000000000000;
	sram_mem[70642] = 16'b0000000000000000;
	sram_mem[70643] = 16'b0000000000000000;
	sram_mem[70644] = 16'b0000000000000000;
	sram_mem[70645] = 16'b0000000000000000;
	sram_mem[70646] = 16'b0000000000000000;
	sram_mem[70647] = 16'b0000000000000000;
	sram_mem[70648] = 16'b0000000000000000;
	sram_mem[70649] = 16'b0000000000000000;
	sram_mem[70650] = 16'b0000000000000000;
	sram_mem[70651] = 16'b0000000000000000;
	sram_mem[70652] = 16'b0000000000000000;
	sram_mem[70653] = 16'b0000000000000000;
	sram_mem[70654] = 16'b0000000000000000;
	sram_mem[70655] = 16'b0000000000000000;
	sram_mem[70656] = 16'b0000000000000000;
	sram_mem[70657] = 16'b0000000000000000;
	sram_mem[70658] = 16'b0000000000000000;
	sram_mem[70659] = 16'b0000000000000000;
	sram_mem[70660] = 16'b0000000000000000;
	sram_mem[70661] = 16'b0000000000000000;
	sram_mem[70662] = 16'b0000000000000000;
	sram_mem[70663] = 16'b0000000000000000;
	sram_mem[70664] = 16'b0000000000000000;
	sram_mem[70665] = 16'b0000000000000000;
	sram_mem[70666] = 16'b0000000000000000;
	sram_mem[70667] = 16'b0000000000000000;
	sram_mem[70668] = 16'b0000000000000000;
	sram_mem[70669] = 16'b0000000000000000;
	sram_mem[70670] = 16'b0000000000000000;
	sram_mem[70671] = 16'b0000000000000000;
	sram_mem[70672] = 16'b0000000000000000;
	sram_mem[70673] = 16'b0000000000000000;
	sram_mem[70674] = 16'b0000000000000000;
	sram_mem[70675] = 16'b0000000000000000;
	sram_mem[70676] = 16'b0000000000000000;
	sram_mem[70677] = 16'b0000000000000000;
	sram_mem[70678] = 16'b0000000000000000;
	sram_mem[70679] = 16'b0000000000000000;
	sram_mem[70680] = 16'b0000000000000000;
	sram_mem[70681] = 16'b0000000000000000;
	sram_mem[70682] = 16'b0000000000000000;
	sram_mem[70683] = 16'b0000000000000000;
	sram_mem[70684] = 16'b0000000000000000;
	sram_mem[70685] = 16'b0000000000000000;
	sram_mem[70686] = 16'b0000000000000000;
	sram_mem[70687] = 16'b0000000000000000;
	sram_mem[70688] = 16'b0000000000000000;
	sram_mem[70689] = 16'b0000000000000000;
	sram_mem[70690] = 16'b0000000000000000;
	sram_mem[70691] = 16'b0000000000000000;
	sram_mem[70692] = 16'b0000000000000000;
	sram_mem[70693] = 16'b0000000000000000;
	sram_mem[70694] = 16'b0000000000000000;
	sram_mem[70695] = 16'b0000000000000000;
	sram_mem[70696] = 16'b0000000000000000;
	sram_mem[70697] = 16'b0000000000000000;
	sram_mem[70698] = 16'b0000000000000000;
	sram_mem[70699] = 16'b0000000000000000;
	sram_mem[70700] = 16'b0000000000000000;
	sram_mem[70701] = 16'b0000000000000000;
	sram_mem[70702] = 16'b0000000000000000;
	sram_mem[70703] = 16'b0000000000000000;
	sram_mem[70704] = 16'b0000000000000000;
	sram_mem[70705] = 16'b0000000000000000;
	sram_mem[70706] = 16'b0000000000000000;
	sram_mem[70707] = 16'b0000000000000000;
	sram_mem[70708] = 16'b0000000000000000;
	sram_mem[70709] = 16'b0000000000000000;
	sram_mem[70710] = 16'b0000000000000000;
	sram_mem[70711] = 16'b0000000000000000;
	sram_mem[70712] = 16'b0000000000000000;
	sram_mem[70713] = 16'b0000000000000000;
	sram_mem[70714] = 16'b0000000000000000;
	sram_mem[70715] = 16'b0000000000000000;
	sram_mem[70716] = 16'b0000000000000000;
	sram_mem[70717] = 16'b0000000000000000;
	sram_mem[70718] = 16'b0000000000000000;
	sram_mem[70719] = 16'b0000000000000000;
	sram_mem[70720] = 16'b0000000000000000;
	sram_mem[70721] = 16'b0000000000000000;
	sram_mem[70722] = 16'b0000000000000000;
	sram_mem[70723] = 16'b0000000000000000;
	sram_mem[70724] = 16'b0000000000000000;
	sram_mem[70725] = 16'b0000000000000000;
	sram_mem[70726] = 16'b0000000000000000;
	sram_mem[70727] = 16'b0000000000000000;
	sram_mem[70728] = 16'b0000000000000000;
	sram_mem[70729] = 16'b0000000000000000;
	sram_mem[70730] = 16'b0000000000000000;
	sram_mem[70731] = 16'b0000000000000000;
	sram_mem[70732] = 16'b0000000000000000;
	sram_mem[70733] = 16'b0000000000000000;
	sram_mem[70734] = 16'b0000000000000000;
	sram_mem[70735] = 16'b0000000000000000;
	sram_mem[70736] = 16'b0000000000000000;
	sram_mem[70737] = 16'b0000000000000000;
	sram_mem[70738] = 16'b0000000000000000;
	sram_mem[70739] = 16'b0000000000000000;
	sram_mem[70740] = 16'b0000000000000000;
	sram_mem[70741] = 16'b0000000000000000;
	sram_mem[70742] = 16'b0000000000000000;
	sram_mem[70743] = 16'b0000000000000000;
	sram_mem[70744] = 16'b0000000000000000;
	sram_mem[70745] = 16'b0000000000000000;
	sram_mem[70746] = 16'b0000000000000000;
	sram_mem[70747] = 16'b0000000000000000;
	sram_mem[70748] = 16'b0000000000000000;
	sram_mem[70749] = 16'b0000000000000000;
	sram_mem[70750] = 16'b0000000000000000;
	sram_mem[70751] = 16'b0000000000000000;
	sram_mem[70752] = 16'b0000000000000000;
	sram_mem[70753] = 16'b0000000000000000;
	sram_mem[70754] = 16'b0000000000000000;
	sram_mem[70755] = 16'b0000000000000000;
	sram_mem[70756] = 16'b0000000000000000;
	sram_mem[70757] = 16'b0000000000000000;
	sram_mem[70758] = 16'b0000000000000000;
	sram_mem[70759] = 16'b0000000000000000;
	sram_mem[70760] = 16'b0000000000000000;
	sram_mem[70761] = 16'b0000000000000000;
	sram_mem[70762] = 16'b0000000000000000;
	sram_mem[70763] = 16'b0000000000000000;
	sram_mem[70764] = 16'b0000000000000000;
	sram_mem[70765] = 16'b0000000000000000;
	sram_mem[70766] = 16'b0000000000000000;
	sram_mem[70767] = 16'b0000000000000000;
	sram_mem[70768] = 16'b0000000000000000;
	sram_mem[70769] = 16'b0000000000000000;
	sram_mem[70770] = 16'b0000000000000000;
	sram_mem[70771] = 16'b0000000000000000;
	sram_mem[70772] = 16'b0000000000000000;
	sram_mem[70773] = 16'b0000000000000000;
	sram_mem[70774] = 16'b0000000000000000;
	sram_mem[70775] = 16'b0000000000000000;
	sram_mem[70776] = 16'b0000000000000000;
	sram_mem[70777] = 16'b0000000000000000;
	sram_mem[70778] = 16'b0000000000000000;
	sram_mem[70779] = 16'b0000000000000000;
	sram_mem[70780] = 16'b0000000000000000;
	sram_mem[70781] = 16'b0000000000000000;
	sram_mem[70782] = 16'b0000000000000000;
	sram_mem[70783] = 16'b0000000000000000;
	sram_mem[70784] = 16'b0000000000000000;
	sram_mem[70785] = 16'b0000000000000000;
	sram_mem[70786] = 16'b0000000000000000;
	sram_mem[70787] = 16'b0000000000000000;
	sram_mem[70788] = 16'b0000000000000000;
	sram_mem[70789] = 16'b0000000000000000;
	sram_mem[70790] = 16'b0000000000000000;
	sram_mem[70791] = 16'b0000000000000000;
	sram_mem[70792] = 16'b0000000000000000;
	sram_mem[70793] = 16'b0000000000000000;
	sram_mem[70794] = 16'b0000000000000000;
	sram_mem[70795] = 16'b0000000000000000;
	sram_mem[70796] = 16'b0000000000000000;
	sram_mem[70797] = 16'b0000000000000000;
	sram_mem[70798] = 16'b0000000000000000;
	sram_mem[70799] = 16'b0000000000000000;
	sram_mem[70800] = 16'b0000000000000000;
	sram_mem[70801] = 16'b0000000000000000;
	sram_mem[70802] = 16'b0000000000000000;
	sram_mem[70803] = 16'b0000000000000000;
	sram_mem[70804] = 16'b0000000000000000;
	sram_mem[70805] = 16'b0000000000000000;
	sram_mem[70806] = 16'b0000000000000000;
	sram_mem[70807] = 16'b0000000000000000;
	sram_mem[70808] = 16'b0000000000000000;
	sram_mem[70809] = 16'b0000000000000000;
	sram_mem[70810] = 16'b0000000000000000;
	sram_mem[70811] = 16'b0000000000000000;
	sram_mem[70812] = 16'b0000000000000000;
	sram_mem[70813] = 16'b0000000000000000;
	sram_mem[70814] = 16'b0000000000000000;
	sram_mem[70815] = 16'b0000000000000000;
	sram_mem[70816] = 16'b0000000000000000;
	sram_mem[70817] = 16'b0000000000000000;
	sram_mem[70818] = 16'b0000000000000000;
	sram_mem[70819] = 16'b0000000000000000;
	sram_mem[70820] = 16'b0000000000000000;
	sram_mem[70821] = 16'b0000000000000000;
	sram_mem[70822] = 16'b0000000000000000;
	sram_mem[70823] = 16'b0000000000000000;
	sram_mem[70824] = 16'b0000000000000000;
	sram_mem[70825] = 16'b0000000000000000;
	sram_mem[70826] = 16'b0000000000000000;
	sram_mem[70827] = 16'b0000000000000000;
	sram_mem[70828] = 16'b0000000000000000;
	sram_mem[70829] = 16'b0000000000000000;
	sram_mem[70830] = 16'b0000000000000000;
	sram_mem[70831] = 16'b0000000000000000;
	sram_mem[70832] = 16'b0000000000000000;
	sram_mem[70833] = 16'b0000000000000000;
	sram_mem[70834] = 16'b0000000000000000;
	sram_mem[70835] = 16'b0000000000000000;
	sram_mem[70836] = 16'b0000000000000000;
	sram_mem[70837] = 16'b0000000000000000;
	sram_mem[70838] = 16'b0000000000000000;
	sram_mem[70839] = 16'b0000000000000000;
	sram_mem[70840] = 16'b0000000000000000;
	sram_mem[70841] = 16'b0000000000000000;
	sram_mem[70842] = 16'b0000000000000000;
	sram_mem[70843] = 16'b0000000000000000;
	sram_mem[70844] = 16'b0000000000000000;
	sram_mem[70845] = 16'b0000000000000000;
	sram_mem[70846] = 16'b0000000000000000;
	sram_mem[70847] = 16'b0000000000000000;
	sram_mem[70848] = 16'b0000000000000000;
	sram_mem[70849] = 16'b0000000000000000;
	sram_mem[70850] = 16'b0000000000000000;
	sram_mem[70851] = 16'b0000000000000000;
	sram_mem[70852] = 16'b0000000000000000;
	sram_mem[70853] = 16'b0000000000000000;
	sram_mem[70854] = 16'b0000000000000000;
	sram_mem[70855] = 16'b0000000000000000;
	sram_mem[70856] = 16'b0000000000000000;
	sram_mem[70857] = 16'b0000000000000000;
	sram_mem[70858] = 16'b0000000000000000;
	sram_mem[70859] = 16'b0000000000000000;
	sram_mem[70860] = 16'b0000000000000000;
	sram_mem[70861] = 16'b0000000000000000;
	sram_mem[70862] = 16'b0000000000000000;
	sram_mem[70863] = 16'b0000000000000000;
	sram_mem[70864] = 16'b0000000000000000;
	sram_mem[70865] = 16'b0000000000000000;
	sram_mem[70866] = 16'b0000000000000000;
	sram_mem[70867] = 16'b0000000000000000;
	sram_mem[70868] = 16'b0000000000000000;
	sram_mem[70869] = 16'b0000000000000000;
	sram_mem[70870] = 16'b0000000000000000;
	sram_mem[70871] = 16'b0000000000000000;
	sram_mem[70872] = 16'b0000000000000000;
	sram_mem[70873] = 16'b0000000000000000;
	sram_mem[70874] = 16'b0000000000000000;
	sram_mem[70875] = 16'b0000000000000000;
	sram_mem[70876] = 16'b0000000000000000;
	sram_mem[70877] = 16'b0000000000000000;
	sram_mem[70878] = 16'b0000000000000000;
	sram_mem[70879] = 16'b0000000000000000;
	sram_mem[70880] = 16'b0000000000000000;
	sram_mem[70881] = 16'b0000000000000000;
	sram_mem[70882] = 16'b0000000000000000;
	sram_mem[70883] = 16'b0000000000000000;
	sram_mem[70884] = 16'b0000000000000000;
	sram_mem[70885] = 16'b0000000000000000;
	sram_mem[70886] = 16'b0000000000000000;
	sram_mem[70887] = 16'b0000000000000000;
	sram_mem[70888] = 16'b0000000000000000;
	sram_mem[70889] = 16'b0000000000000000;
	sram_mem[70890] = 16'b0000000000000000;
	sram_mem[70891] = 16'b0000000000000000;
	sram_mem[70892] = 16'b0000000000000000;
	sram_mem[70893] = 16'b0000000000000000;
	sram_mem[70894] = 16'b0000000000000000;
	sram_mem[70895] = 16'b0000000000000000;
	sram_mem[70896] = 16'b0000000000000000;
	sram_mem[70897] = 16'b0000000000000000;
	sram_mem[70898] = 16'b0000000000000000;
	sram_mem[70899] = 16'b0000000000000000;
	sram_mem[70900] = 16'b0000000000000000;
	sram_mem[70901] = 16'b0000000000000000;
	sram_mem[70902] = 16'b0000000000000000;
	sram_mem[70903] = 16'b0000000000000000;
	sram_mem[70904] = 16'b0000000000000000;
	sram_mem[70905] = 16'b0000000000000000;
	sram_mem[70906] = 16'b0000000000000000;
	sram_mem[70907] = 16'b0000000000000000;
	sram_mem[70908] = 16'b0000000000000000;
	sram_mem[70909] = 16'b0000000000000000;
	sram_mem[70910] = 16'b0000000000000000;
	sram_mem[70911] = 16'b0000000000000000;
	sram_mem[70912] = 16'b0000000000000000;
	sram_mem[70913] = 16'b0000000000000000;
	sram_mem[70914] = 16'b0000000000000000;
	sram_mem[70915] = 16'b0000000000000000;
	sram_mem[70916] = 16'b0000000000000000;
	sram_mem[70917] = 16'b0000000000000000;
	sram_mem[70918] = 16'b0000000000000000;
	sram_mem[70919] = 16'b0000000000000000;
	sram_mem[70920] = 16'b0000000000000000;
	sram_mem[70921] = 16'b0000000000000000;
	sram_mem[70922] = 16'b0000000000000000;
	sram_mem[70923] = 16'b0000000000000000;
	sram_mem[70924] = 16'b0000000000000000;
	sram_mem[70925] = 16'b0000000000000000;
	sram_mem[70926] = 16'b0000000000000000;
	sram_mem[70927] = 16'b0000000000000000;
	sram_mem[70928] = 16'b0000000000000000;
	sram_mem[70929] = 16'b0000000000000000;
	sram_mem[70930] = 16'b0000000000000000;
	sram_mem[70931] = 16'b0000000000000000;
	sram_mem[70932] = 16'b0000000000000000;
	sram_mem[70933] = 16'b0000000000000000;
	sram_mem[70934] = 16'b0000000000000000;
	sram_mem[70935] = 16'b0000000000000000;
	sram_mem[70936] = 16'b0000000000000000;
	sram_mem[70937] = 16'b0000000000000000;
	sram_mem[70938] = 16'b0000000000000000;
	sram_mem[70939] = 16'b0000000000000000;
	sram_mem[70940] = 16'b0000000000000000;
	sram_mem[70941] = 16'b0000000000000000;
	sram_mem[70942] = 16'b0000000000000000;
	sram_mem[70943] = 16'b0000000000000000;
	sram_mem[70944] = 16'b0000000000000000;
	sram_mem[70945] = 16'b0000000000000000;
	sram_mem[70946] = 16'b0000000000000000;
	sram_mem[70947] = 16'b0000000000000000;
	sram_mem[70948] = 16'b0000000000000000;
	sram_mem[70949] = 16'b0000000000000000;
	sram_mem[70950] = 16'b0000000000000000;
	sram_mem[70951] = 16'b0000000000000000;
	sram_mem[70952] = 16'b0000000000000000;
	sram_mem[70953] = 16'b0000000000000000;
	sram_mem[70954] = 16'b0000000000000000;
	sram_mem[70955] = 16'b0000000000000000;
	sram_mem[70956] = 16'b0000000000000000;
	sram_mem[70957] = 16'b0000000000000000;
	sram_mem[70958] = 16'b0000000000000000;
	sram_mem[70959] = 16'b0000000000000000;
	sram_mem[70960] = 16'b0000000000000000;
	sram_mem[70961] = 16'b0000000000000000;
	sram_mem[70962] = 16'b0000000000000000;
	sram_mem[70963] = 16'b0000000000000000;
	sram_mem[70964] = 16'b0000000000000000;
	sram_mem[70965] = 16'b0000000000000000;
	sram_mem[70966] = 16'b0000000000000000;
	sram_mem[70967] = 16'b0000000000000000;
	sram_mem[70968] = 16'b0000000000000000;
	sram_mem[70969] = 16'b0000000000000000;
	sram_mem[70970] = 16'b0000000000000000;
	sram_mem[70971] = 16'b0000000000000000;
	sram_mem[70972] = 16'b0000000000000000;
	sram_mem[70973] = 16'b0000000000000000;
	sram_mem[70974] = 16'b0000000000000000;
	sram_mem[70975] = 16'b0000000000000000;
	sram_mem[70976] = 16'b0000000000000000;
	sram_mem[70977] = 16'b0000000000000000;
	sram_mem[70978] = 16'b0000000000000000;
	sram_mem[70979] = 16'b0000000000000000;
	sram_mem[70980] = 16'b0000000000000000;
	sram_mem[70981] = 16'b0000000000000000;
	sram_mem[70982] = 16'b0000000000000000;
	sram_mem[70983] = 16'b0000000000000000;
	sram_mem[70984] = 16'b0000000000000000;
	sram_mem[70985] = 16'b0000000000000000;
	sram_mem[70986] = 16'b0000000000000000;
	sram_mem[70987] = 16'b0000000000000000;
	sram_mem[70988] = 16'b0000000000000000;
	sram_mem[70989] = 16'b0000000000000000;
	sram_mem[70990] = 16'b0000000000000000;
	sram_mem[70991] = 16'b0000000000000000;
	sram_mem[70992] = 16'b0000000000000000;
	sram_mem[70993] = 16'b0000000000000000;
	sram_mem[70994] = 16'b0000000000000000;
	sram_mem[70995] = 16'b0000000000000000;
	sram_mem[70996] = 16'b0000000000000000;
	sram_mem[70997] = 16'b0000000000000000;
	sram_mem[70998] = 16'b0000000000000000;
	sram_mem[70999] = 16'b0000000000000000;
	sram_mem[71000] = 16'b0000000000000000;
	sram_mem[71001] = 16'b0000000000000000;
	sram_mem[71002] = 16'b0000000000000000;
	sram_mem[71003] = 16'b0000000000000000;
	sram_mem[71004] = 16'b0000000000000000;
	sram_mem[71005] = 16'b0000000000000000;
	sram_mem[71006] = 16'b0000000000000000;
	sram_mem[71007] = 16'b0000000000000000;
	sram_mem[71008] = 16'b0000000000000000;
	sram_mem[71009] = 16'b0000000000000000;
	sram_mem[71010] = 16'b0000000000000000;
	sram_mem[71011] = 16'b0000000000000000;
	sram_mem[71012] = 16'b0000000000000000;
	sram_mem[71013] = 16'b0000000000000000;
	sram_mem[71014] = 16'b0000000000000000;
	sram_mem[71015] = 16'b0000000000000000;
	sram_mem[71016] = 16'b0000000000000000;
	sram_mem[71017] = 16'b0000000000000000;
	sram_mem[71018] = 16'b0000000000000000;
	sram_mem[71019] = 16'b0000000000000000;
	sram_mem[71020] = 16'b0000000000000000;
	sram_mem[71021] = 16'b0000000000000000;
	sram_mem[71022] = 16'b0000000000000000;
	sram_mem[71023] = 16'b0000000000000000;
	sram_mem[71024] = 16'b0000000000000000;
	sram_mem[71025] = 16'b0000000000000000;
	sram_mem[71026] = 16'b0000000000000000;
	sram_mem[71027] = 16'b0000000000000000;
	sram_mem[71028] = 16'b0000000000000000;
	sram_mem[71029] = 16'b0000000000000000;
	sram_mem[71030] = 16'b0000000000000000;
	sram_mem[71031] = 16'b0000000000000000;
	sram_mem[71032] = 16'b0000000000000000;
	sram_mem[71033] = 16'b0000000000000000;
	sram_mem[71034] = 16'b0000000000000000;
	sram_mem[71035] = 16'b0000000000000000;
	sram_mem[71036] = 16'b0000000000000000;
	sram_mem[71037] = 16'b0000000000000000;
	sram_mem[71038] = 16'b0000000000000000;
	sram_mem[71039] = 16'b0000000000000000;
	sram_mem[71040] = 16'b0000000000000000;
	sram_mem[71041] = 16'b0000000000000000;
	sram_mem[71042] = 16'b0000000000000000;
	sram_mem[71043] = 16'b0000000000000000;
	sram_mem[71044] = 16'b0000000000000000;
	sram_mem[71045] = 16'b0000000000000000;
	sram_mem[71046] = 16'b0000000000000000;
	sram_mem[71047] = 16'b0000000000000000;
	sram_mem[71048] = 16'b0000000000000000;
	sram_mem[71049] = 16'b0000000000000000;
	sram_mem[71050] = 16'b0000000000000000;
	sram_mem[71051] = 16'b0000000000000000;
	sram_mem[71052] = 16'b0000000000000000;
	sram_mem[71053] = 16'b0000000000000000;
	sram_mem[71054] = 16'b0000000000000000;
	sram_mem[71055] = 16'b0000000000000000;
	sram_mem[71056] = 16'b0000000000000000;
	sram_mem[71057] = 16'b0000000000000000;
	sram_mem[71058] = 16'b0000000000000000;
	sram_mem[71059] = 16'b0000000000000000;
	sram_mem[71060] = 16'b0000000000000000;
	sram_mem[71061] = 16'b0000000000000000;
	sram_mem[71062] = 16'b0000000000000000;
	sram_mem[71063] = 16'b0000000000000000;
	sram_mem[71064] = 16'b0000000000000000;
	sram_mem[71065] = 16'b0000000000000000;
	sram_mem[71066] = 16'b0000000000000000;
	sram_mem[71067] = 16'b0000000000000000;
	sram_mem[71068] = 16'b0000000000000000;
	sram_mem[71069] = 16'b0000000000000000;
	sram_mem[71070] = 16'b0000000000000000;
	sram_mem[71071] = 16'b0000000000000000;
	sram_mem[71072] = 16'b0000000000000000;
	sram_mem[71073] = 16'b0000000000000000;
	sram_mem[71074] = 16'b0000000000000000;
	sram_mem[71075] = 16'b0000000000000000;
	sram_mem[71076] = 16'b0000000000000000;
	sram_mem[71077] = 16'b0000000000000000;
	sram_mem[71078] = 16'b0000000000000000;
	sram_mem[71079] = 16'b0000000000000000;
	sram_mem[71080] = 16'b0000000000000000;
	sram_mem[71081] = 16'b0000000000000000;
	sram_mem[71082] = 16'b0000000000000000;
	sram_mem[71083] = 16'b0000000000000000;
	sram_mem[71084] = 16'b0000000000000000;
	sram_mem[71085] = 16'b0000000000000000;
	sram_mem[71086] = 16'b0000000000000000;
	sram_mem[71087] = 16'b0000000000000000;
	sram_mem[71088] = 16'b0000000000000000;
	sram_mem[71089] = 16'b0000000000000000;
	sram_mem[71090] = 16'b0000000000000000;
	sram_mem[71091] = 16'b0000000000000000;
	sram_mem[71092] = 16'b0000000000000000;
	sram_mem[71093] = 16'b0000000000000000;
	sram_mem[71094] = 16'b0000000000000000;
	sram_mem[71095] = 16'b0000000000000000;
	sram_mem[71096] = 16'b0000000000000000;
	sram_mem[71097] = 16'b0000000000000000;
	sram_mem[71098] = 16'b0000000000000000;
	sram_mem[71099] = 16'b0000000000000000;
	sram_mem[71100] = 16'b0000000000000000;
	sram_mem[71101] = 16'b0000000000000000;
	sram_mem[71102] = 16'b0000000000000000;
	sram_mem[71103] = 16'b0000000000000000;
	sram_mem[71104] = 16'b0000000000000000;
	sram_mem[71105] = 16'b0000000000000000;
	sram_mem[71106] = 16'b0000000000000000;
	sram_mem[71107] = 16'b0000000000000000;
	sram_mem[71108] = 16'b0000000000000000;
	sram_mem[71109] = 16'b0000000000000000;
	sram_mem[71110] = 16'b0000000000000000;
	sram_mem[71111] = 16'b0000000000000000;
	sram_mem[71112] = 16'b0000000000000000;
	sram_mem[71113] = 16'b0000000000000000;
	sram_mem[71114] = 16'b0000000000000000;
	sram_mem[71115] = 16'b0000000000000000;
	sram_mem[71116] = 16'b0000000000000000;
	sram_mem[71117] = 16'b0000000000000000;
	sram_mem[71118] = 16'b0000000000000000;
	sram_mem[71119] = 16'b0000000000000000;
	sram_mem[71120] = 16'b0000000000000000;
	sram_mem[71121] = 16'b0000000000000000;
	sram_mem[71122] = 16'b0000000000000000;
	sram_mem[71123] = 16'b0000000000000000;
	sram_mem[71124] = 16'b0000000000000000;
	sram_mem[71125] = 16'b0000000000000000;
	sram_mem[71126] = 16'b0000000000000000;
	sram_mem[71127] = 16'b0000000000000000;
	sram_mem[71128] = 16'b0000000000000000;
	sram_mem[71129] = 16'b0000000000000000;
	sram_mem[71130] = 16'b0000000000000000;
	sram_mem[71131] = 16'b0000000000000000;
	sram_mem[71132] = 16'b0000000000000000;
	sram_mem[71133] = 16'b0000000000000000;
	sram_mem[71134] = 16'b0000000000000000;
	sram_mem[71135] = 16'b0000000000000000;
	sram_mem[71136] = 16'b0000000000000000;
	sram_mem[71137] = 16'b0000000000000000;
	sram_mem[71138] = 16'b0000000000000000;
	sram_mem[71139] = 16'b0000000000000000;
	sram_mem[71140] = 16'b0000000000000000;
	sram_mem[71141] = 16'b0000000000000000;
	sram_mem[71142] = 16'b0000000000000000;
	sram_mem[71143] = 16'b0000000000000000;
	sram_mem[71144] = 16'b0000000000000000;
	sram_mem[71145] = 16'b0000000000000000;
	sram_mem[71146] = 16'b0000000000000000;
	sram_mem[71147] = 16'b0000000000000000;
	sram_mem[71148] = 16'b0000000000000000;
	sram_mem[71149] = 16'b0000000000000000;
	sram_mem[71150] = 16'b0000000000000000;
	sram_mem[71151] = 16'b0000000000000000;
	sram_mem[71152] = 16'b0000000000000000;
	sram_mem[71153] = 16'b0000000000000000;
	sram_mem[71154] = 16'b0000000000000000;
	sram_mem[71155] = 16'b0000000000000000;
	sram_mem[71156] = 16'b0000000000000000;
	sram_mem[71157] = 16'b0000000000000000;
	sram_mem[71158] = 16'b0000000000000000;
	sram_mem[71159] = 16'b0000000000000000;
	sram_mem[71160] = 16'b0000000000000000;
	sram_mem[71161] = 16'b0000000000000000;
	sram_mem[71162] = 16'b0000000000000000;
	sram_mem[71163] = 16'b0000000000000000;
	sram_mem[71164] = 16'b0000000000000000;
	sram_mem[71165] = 16'b0000000000000000;
	sram_mem[71166] = 16'b0000000000000000;
	sram_mem[71167] = 16'b0000000000000000;
	sram_mem[71168] = 16'b0000000000000000;
	sram_mem[71169] = 16'b0000000000000000;
	sram_mem[71170] = 16'b0000000000000000;
	sram_mem[71171] = 16'b0000000000000000;
	sram_mem[71172] = 16'b0000000000000000;
	sram_mem[71173] = 16'b0000000000000000;
	sram_mem[71174] = 16'b0000000000000000;
	sram_mem[71175] = 16'b0000000000000000;
	sram_mem[71176] = 16'b0000000000000000;
	sram_mem[71177] = 16'b0000000000000000;
	sram_mem[71178] = 16'b0000000000000000;
	sram_mem[71179] = 16'b0000000000000000;
	sram_mem[71180] = 16'b0000000000000000;
	sram_mem[71181] = 16'b0000000000000000;
	sram_mem[71182] = 16'b0000000000000000;
	sram_mem[71183] = 16'b0000000000000000;
	sram_mem[71184] = 16'b0000000000000000;
	sram_mem[71185] = 16'b0000000000000000;
	sram_mem[71186] = 16'b0000000000000000;
	sram_mem[71187] = 16'b0000000000000000;
	sram_mem[71188] = 16'b0000000000000000;
	sram_mem[71189] = 16'b0000000000000000;
	sram_mem[71190] = 16'b0000000000000000;
	sram_mem[71191] = 16'b0000000000000000;
	sram_mem[71192] = 16'b0000000000000000;
	sram_mem[71193] = 16'b0000000000000000;
	sram_mem[71194] = 16'b0000000000000000;
	sram_mem[71195] = 16'b0000000000000000;
	sram_mem[71196] = 16'b0000000000000000;
	sram_mem[71197] = 16'b0000000000000000;
	sram_mem[71198] = 16'b0000000000000000;
	sram_mem[71199] = 16'b0000000000000000;
	sram_mem[71200] = 16'b0000000000000000;
	sram_mem[71201] = 16'b0000000000000000;
	sram_mem[71202] = 16'b0000000000000000;
	sram_mem[71203] = 16'b0000000000000000;
	sram_mem[71204] = 16'b0000000000000000;
	sram_mem[71205] = 16'b0000000000000000;
	sram_mem[71206] = 16'b0000000000000000;
	sram_mem[71207] = 16'b0000000000000000;
	sram_mem[71208] = 16'b0000000000000000;
	sram_mem[71209] = 16'b0000000000000000;
	sram_mem[71210] = 16'b0000000000000000;
	sram_mem[71211] = 16'b0000000000000000;
	sram_mem[71212] = 16'b0000000000000000;
	sram_mem[71213] = 16'b0000000000000000;
	sram_mem[71214] = 16'b0000000000000000;
	sram_mem[71215] = 16'b0000000000000000;
	sram_mem[71216] = 16'b0000000000000000;
	sram_mem[71217] = 16'b0000000000000000;
	sram_mem[71218] = 16'b0000000000000000;
	sram_mem[71219] = 16'b0000000000000000;
	sram_mem[71220] = 16'b0000000000000000;
	sram_mem[71221] = 16'b0000000000000000;
	sram_mem[71222] = 16'b0000000000000000;
	sram_mem[71223] = 16'b0000000000000000;
	sram_mem[71224] = 16'b0000000000000000;
	sram_mem[71225] = 16'b0000000000000000;
	sram_mem[71226] = 16'b0000000000000000;
	sram_mem[71227] = 16'b0000000000000000;
	sram_mem[71228] = 16'b0000000000000000;
	sram_mem[71229] = 16'b0000000000000000;
	sram_mem[71230] = 16'b0000000000000000;
	sram_mem[71231] = 16'b0000000000000000;
	sram_mem[71232] = 16'b0000000000000000;
	sram_mem[71233] = 16'b0000000000000000;
	sram_mem[71234] = 16'b0000000000000000;
	sram_mem[71235] = 16'b0000000000000000;
	sram_mem[71236] = 16'b0000000000000000;
	sram_mem[71237] = 16'b0000000000000000;
	sram_mem[71238] = 16'b0000000000000000;
	sram_mem[71239] = 16'b0000000000000000;
	sram_mem[71240] = 16'b0000000000000000;
	sram_mem[71241] = 16'b0000000000000000;
	sram_mem[71242] = 16'b0000000000000000;
	sram_mem[71243] = 16'b0000000000000000;
	sram_mem[71244] = 16'b0000000000000000;
	sram_mem[71245] = 16'b0000000000000000;
	sram_mem[71246] = 16'b0000000000000000;
	sram_mem[71247] = 16'b0000000000000000;
	sram_mem[71248] = 16'b0000000000000000;
	sram_mem[71249] = 16'b0000000000000000;
	sram_mem[71250] = 16'b0000000000000000;
	sram_mem[71251] = 16'b0000000000000000;
	sram_mem[71252] = 16'b0000000000000000;
	sram_mem[71253] = 16'b0000000000000000;
	sram_mem[71254] = 16'b0000000000000000;
	sram_mem[71255] = 16'b0000000000000000;
	sram_mem[71256] = 16'b0000000000000000;
	sram_mem[71257] = 16'b0000000000000000;
	sram_mem[71258] = 16'b0000000000000000;
	sram_mem[71259] = 16'b0000000000000000;
	sram_mem[71260] = 16'b0000000000000000;
	sram_mem[71261] = 16'b0000000000000000;
	sram_mem[71262] = 16'b0000000000000000;
	sram_mem[71263] = 16'b0000000000000000;
	sram_mem[71264] = 16'b0000000000000000;
	sram_mem[71265] = 16'b0000000000000000;
	sram_mem[71266] = 16'b0000000000000000;
	sram_mem[71267] = 16'b0000000000000000;
	sram_mem[71268] = 16'b0000000000000000;
	sram_mem[71269] = 16'b0000000000000000;
	sram_mem[71270] = 16'b0000000000000000;
	sram_mem[71271] = 16'b0000000000000000;
	sram_mem[71272] = 16'b0000000000000000;
	sram_mem[71273] = 16'b0000000000000000;
	sram_mem[71274] = 16'b0000000000000000;
	sram_mem[71275] = 16'b0000000000000000;
	sram_mem[71276] = 16'b0000000000000000;
	sram_mem[71277] = 16'b0000000000000000;
	sram_mem[71278] = 16'b0000000000000000;
	sram_mem[71279] = 16'b0000000000000000;
	sram_mem[71280] = 16'b0000000000000000;
	sram_mem[71281] = 16'b0000000000000000;
	sram_mem[71282] = 16'b0000000000000000;
	sram_mem[71283] = 16'b0000000000000000;
	sram_mem[71284] = 16'b0000000000000000;
	sram_mem[71285] = 16'b0000000000000000;
	sram_mem[71286] = 16'b0000000000000000;
	sram_mem[71287] = 16'b0000000000000000;
	sram_mem[71288] = 16'b0000000000000000;
	sram_mem[71289] = 16'b0000000000000000;
	sram_mem[71290] = 16'b0000000000000000;
	sram_mem[71291] = 16'b0000000000000000;
	sram_mem[71292] = 16'b0000000000000000;
	sram_mem[71293] = 16'b0000000000000000;
	sram_mem[71294] = 16'b0000000000000000;
	sram_mem[71295] = 16'b0000000000000000;
	sram_mem[71296] = 16'b0000000000000000;
	sram_mem[71297] = 16'b0000000000000000;
	sram_mem[71298] = 16'b0000000000000000;
	sram_mem[71299] = 16'b0000000000000000;
	sram_mem[71300] = 16'b0000000000000000;
	sram_mem[71301] = 16'b0000000000000000;
	sram_mem[71302] = 16'b0000000000000000;
	sram_mem[71303] = 16'b0000000000000000;
	sram_mem[71304] = 16'b0000000000000000;
	sram_mem[71305] = 16'b0000000000000000;
	sram_mem[71306] = 16'b0000000000000000;
	sram_mem[71307] = 16'b0000000000000000;
	sram_mem[71308] = 16'b0000000000000000;
	sram_mem[71309] = 16'b0000000000000000;
	sram_mem[71310] = 16'b0000000000000000;
	sram_mem[71311] = 16'b0000000000000000;
	sram_mem[71312] = 16'b0000000000000000;
	sram_mem[71313] = 16'b0000000000000000;
	sram_mem[71314] = 16'b0000000000000000;
	sram_mem[71315] = 16'b0000000000000000;
	sram_mem[71316] = 16'b0000000000000000;
	sram_mem[71317] = 16'b0000000000000000;
	sram_mem[71318] = 16'b0000000000000000;
	sram_mem[71319] = 16'b0000000000000000;
	sram_mem[71320] = 16'b0000000000000000;
	sram_mem[71321] = 16'b0000000000000000;
	sram_mem[71322] = 16'b0000000000000000;
	sram_mem[71323] = 16'b0000000000000000;
	sram_mem[71324] = 16'b0000000000000000;
	sram_mem[71325] = 16'b0000000000000000;
	sram_mem[71326] = 16'b0000000000000000;
	sram_mem[71327] = 16'b0000000000000000;
	sram_mem[71328] = 16'b0000000000000000;
	sram_mem[71329] = 16'b0000000000000000;
	sram_mem[71330] = 16'b0000000000000000;
	sram_mem[71331] = 16'b0000000000000000;
	sram_mem[71332] = 16'b0000000000000000;
	sram_mem[71333] = 16'b0000000000000000;
	sram_mem[71334] = 16'b0000000000000000;
	sram_mem[71335] = 16'b0000000000000000;
	sram_mem[71336] = 16'b0000000000000000;
	sram_mem[71337] = 16'b0000000000000000;
	sram_mem[71338] = 16'b0000000000000000;
	sram_mem[71339] = 16'b0000000000000000;
	sram_mem[71340] = 16'b0000000000000000;
	sram_mem[71341] = 16'b0000000000000000;
	sram_mem[71342] = 16'b0000000000000000;
	sram_mem[71343] = 16'b0000000000000000;
	sram_mem[71344] = 16'b0000000000000000;
	sram_mem[71345] = 16'b0000000000000000;
	sram_mem[71346] = 16'b0000000000000000;
	sram_mem[71347] = 16'b0000000000000000;
	sram_mem[71348] = 16'b0000000000000000;
	sram_mem[71349] = 16'b0000000000000000;
	sram_mem[71350] = 16'b0000000000000000;
	sram_mem[71351] = 16'b0000000000000000;
	sram_mem[71352] = 16'b0000000000000000;
	sram_mem[71353] = 16'b0000000000000000;
	sram_mem[71354] = 16'b0000000000000000;
	sram_mem[71355] = 16'b0000000000000000;
	sram_mem[71356] = 16'b0000000000000000;
	sram_mem[71357] = 16'b0000000000000000;
	sram_mem[71358] = 16'b0000000000000000;
	sram_mem[71359] = 16'b0000000000000000;
	sram_mem[71360] = 16'b0000000000000000;
	sram_mem[71361] = 16'b0000000000000000;
	sram_mem[71362] = 16'b0000000000000000;
	sram_mem[71363] = 16'b0000000000000000;
	sram_mem[71364] = 16'b0000000000000000;
	sram_mem[71365] = 16'b0000000000000000;
	sram_mem[71366] = 16'b0000000000000000;
	sram_mem[71367] = 16'b0000000000000000;
	sram_mem[71368] = 16'b0000000000000000;
	sram_mem[71369] = 16'b0000000000000000;
	sram_mem[71370] = 16'b0000000000000000;
	sram_mem[71371] = 16'b0000000000000000;
	sram_mem[71372] = 16'b0000000000000000;
	sram_mem[71373] = 16'b0000000000000000;
	sram_mem[71374] = 16'b0000000000000000;
	sram_mem[71375] = 16'b0000000000000000;
	sram_mem[71376] = 16'b0000000000000000;
	sram_mem[71377] = 16'b0000000000000000;
	sram_mem[71378] = 16'b0000000000000000;
	sram_mem[71379] = 16'b0000000000000000;
	sram_mem[71380] = 16'b0000000000000000;
	sram_mem[71381] = 16'b0000000000000000;
	sram_mem[71382] = 16'b0000000000000000;
	sram_mem[71383] = 16'b0000000000000000;
	sram_mem[71384] = 16'b0000000000000000;
	sram_mem[71385] = 16'b0000000000000000;
	sram_mem[71386] = 16'b0000000000000000;
	sram_mem[71387] = 16'b0000000000000000;
	sram_mem[71388] = 16'b0000000000000000;
	sram_mem[71389] = 16'b0000000000000000;
	sram_mem[71390] = 16'b0000000000000000;
	sram_mem[71391] = 16'b0000000000000000;
	sram_mem[71392] = 16'b0000000000000000;
	sram_mem[71393] = 16'b0000000000000000;
	sram_mem[71394] = 16'b0000000000000000;
	sram_mem[71395] = 16'b0000000000000000;
	sram_mem[71396] = 16'b0000000000000000;
	sram_mem[71397] = 16'b0000000000000000;
	sram_mem[71398] = 16'b0000000000000000;
	sram_mem[71399] = 16'b0000000000000000;
	sram_mem[71400] = 16'b0000000000000000;
	sram_mem[71401] = 16'b0000000000000000;
	sram_mem[71402] = 16'b0000000000000000;
	sram_mem[71403] = 16'b0000000000000000;
	sram_mem[71404] = 16'b0000000000000000;
	sram_mem[71405] = 16'b0000000000000000;
	sram_mem[71406] = 16'b0000000000000000;
	sram_mem[71407] = 16'b0000000000000000;
	sram_mem[71408] = 16'b0000000000000000;
	sram_mem[71409] = 16'b0000000000000000;
	sram_mem[71410] = 16'b0000000000000000;
	sram_mem[71411] = 16'b0000000000000000;
	sram_mem[71412] = 16'b0000000000000000;
	sram_mem[71413] = 16'b0000000000000000;
	sram_mem[71414] = 16'b0000000000000000;
	sram_mem[71415] = 16'b0000000000000000;
	sram_mem[71416] = 16'b0000000000000000;
	sram_mem[71417] = 16'b0000000000000000;
	sram_mem[71418] = 16'b0000000000000000;
	sram_mem[71419] = 16'b0000000000000000;
	sram_mem[71420] = 16'b0000000000000000;
	sram_mem[71421] = 16'b0000000000000000;
	sram_mem[71422] = 16'b0000000000000000;
	sram_mem[71423] = 16'b0000000000000000;
	sram_mem[71424] = 16'b0000000000000000;
	sram_mem[71425] = 16'b0000000000000000;
	sram_mem[71426] = 16'b0000000000000000;
	sram_mem[71427] = 16'b0000000000000000;
	sram_mem[71428] = 16'b0000000000000000;
	sram_mem[71429] = 16'b0000000000000000;
	sram_mem[71430] = 16'b0000000000000000;
	sram_mem[71431] = 16'b0000000000000000;
	sram_mem[71432] = 16'b0000000000000000;
	sram_mem[71433] = 16'b0000000000000000;
	sram_mem[71434] = 16'b0000000000000000;
	sram_mem[71435] = 16'b0000000000000000;
	sram_mem[71436] = 16'b0000000000000000;
	sram_mem[71437] = 16'b0000000000000000;
	sram_mem[71438] = 16'b0000000000000000;
	sram_mem[71439] = 16'b0000000000000000;
	sram_mem[71440] = 16'b0000000000000000;
	sram_mem[71441] = 16'b0000000000000000;
	sram_mem[71442] = 16'b0000000000000000;
	sram_mem[71443] = 16'b0000000000000000;
	sram_mem[71444] = 16'b0000000000000000;
	sram_mem[71445] = 16'b0000000000000000;
	sram_mem[71446] = 16'b0000000000000000;
	sram_mem[71447] = 16'b0000000000000000;
	sram_mem[71448] = 16'b0000000000000000;
	sram_mem[71449] = 16'b0000000000000000;
	sram_mem[71450] = 16'b0000000000000000;
	sram_mem[71451] = 16'b0000000000000000;
	sram_mem[71452] = 16'b0000000000000000;
	sram_mem[71453] = 16'b0000000000000000;
	sram_mem[71454] = 16'b0000000000000000;
	sram_mem[71455] = 16'b0000000000000000;
	sram_mem[71456] = 16'b0000000000000000;
	sram_mem[71457] = 16'b0000000000000000;
	sram_mem[71458] = 16'b0000000000000000;
	sram_mem[71459] = 16'b0000000000000000;
	sram_mem[71460] = 16'b0000000000000000;
	sram_mem[71461] = 16'b0000000000000000;
	sram_mem[71462] = 16'b0000000000000000;
	sram_mem[71463] = 16'b0000000000000000;
	sram_mem[71464] = 16'b0000000000000000;
	sram_mem[71465] = 16'b0000000000000000;
	sram_mem[71466] = 16'b0000000000000000;
	sram_mem[71467] = 16'b0000000000000000;
	sram_mem[71468] = 16'b0000000000000000;
	sram_mem[71469] = 16'b0000000000000000;
	sram_mem[71470] = 16'b0000000000000000;
	sram_mem[71471] = 16'b0000000000000000;
	sram_mem[71472] = 16'b0000000000000000;
	sram_mem[71473] = 16'b0000000000000000;
	sram_mem[71474] = 16'b0000000000000000;
	sram_mem[71475] = 16'b0000000000000000;
	sram_mem[71476] = 16'b0000000000000000;
	sram_mem[71477] = 16'b0000000000000000;
	sram_mem[71478] = 16'b0000000000000000;
	sram_mem[71479] = 16'b0000000000000000;
	sram_mem[71480] = 16'b0000000000000000;
	sram_mem[71481] = 16'b0000000000000000;
	sram_mem[71482] = 16'b0000000000000000;
	sram_mem[71483] = 16'b0000000000000000;
	sram_mem[71484] = 16'b0000000000000000;
	sram_mem[71485] = 16'b0000000000000000;
	sram_mem[71486] = 16'b0000000000000000;
	sram_mem[71487] = 16'b0000000000000000;
	sram_mem[71488] = 16'b0000000000000000;
	sram_mem[71489] = 16'b0000000000000000;
	sram_mem[71490] = 16'b0000000000000000;
	sram_mem[71491] = 16'b0000000000000000;
	sram_mem[71492] = 16'b0000000000000000;
	sram_mem[71493] = 16'b0000000000000000;
	sram_mem[71494] = 16'b0000000000000000;
	sram_mem[71495] = 16'b0000000000000000;
	sram_mem[71496] = 16'b0000000000000000;
	sram_mem[71497] = 16'b0000000000000000;
	sram_mem[71498] = 16'b0000000000000000;
	sram_mem[71499] = 16'b0000000000000000;
	sram_mem[71500] = 16'b0000000000000000;
	sram_mem[71501] = 16'b0000000000000000;
	sram_mem[71502] = 16'b0000000000000000;
	sram_mem[71503] = 16'b0000000000000000;
	sram_mem[71504] = 16'b0000000000000000;
	sram_mem[71505] = 16'b0000000000000000;
	sram_mem[71506] = 16'b0000000000000000;
	sram_mem[71507] = 16'b0000000000000000;
	sram_mem[71508] = 16'b0000000000000000;
	sram_mem[71509] = 16'b0000000000000000;
	sram_mem[71510] = 16'b0000000000000000;
	sram_mem[71511] = 16'b0000000000000000;
	sram_mem[71512] = 16'b0000000000000000;
	sram_mem[71513] = 16'b0000000000000000;
	sram_mem[71514] = 16'b0000000000000000;
	sram_mem[71515] = 16'b0000000000000000;
	sram_mem[71516] = 16'b0000000000000000;
	sram_mem[71517] = 16'b0000000000000000;
	sram_mem[71518] = 16'b0000000000000000;
	sram_mem[71519] = 16'b0000000000000000;
	sram_mem[71520] = 16'b0000000000000000;
	sram_mem[71521] = 16'b0000000000000000;
	sram_mem[71522] = 16'b0000000000000000;
	sram_mem[71523] = 16'b0000000000000000;
	sram_mem[71524] = 16'b0000000000000000;
	sram_mem[71525] = 16'b0000000000000000;
	sram_mem[71526] = 16'b0000000000000000;
	sram_mem[71527] = 16'b0000000000000000;
	sram_mem[71528] = 16'b0000000000000000;
	sram_mem[71529] = 16'b0000000000000000;
	sram_mem[71530] = 16'b0000000000000000;
	sram_mem[71531] = 16'b0000000000000000;
	sram_mem[71532] = 16'b0000000000000000;
	sram_mem[71533] = 16'b0000000000000000;
	sram_mem[71534] = 16'b0000000000000000;
	sram_mem[71535] = 16'b0000000000000000;
	sram_mem[71536] = 16'b0000000000000000;
	sram_mem[71537] = 16'b0000000000000000;
	sram_mem[71538] = 16'b0000000000000000;
	sram_mem[71539] = 16'b0000000000000000;
	sram_mem[71540] = 16'b0000000000000000;
	sram_mem[71541] = 16'b0000000000000000;
	sram_mem[71542] = 16'b0000000000000000;
	sram_mem[71543] = 16'b0000000000000000;
	sram_mem[71544] = 16'b0000000000000000;
	sram_mem[71545] = 16'b0000000000000000;
	sram_mem[71546] = 16'b0000000000000000;
	sram_mem[71547] = 16'b0000000000000000;
	sram_mem[71548] = 16'b0000000000000000;
	sram_mem[71549] = 16'b0000000000000000;
	sram_mem[71550] = 16'b0000000000000000;
	sram_mem[71551] = 16'b0000000000000000;
	sram_mem[71552] = 16'b0000000000000000;
	sram_mem[71553] = 16'b0000000000000000;
	sram_mem[71554] = 16'b0000000000000000;
	sram_mem[71555] = 16'b0000000000000000;
	sram_mem[71556] = 16'b0000000000000000;
	sram_mem[71557] = 16'b0000000000000000;
	sram_mem[71558] = 16'b0000000000000000;
	sram_mem[71559] = 16'b0000000000000000;
	sram_mem[71560] = 16'b0000000000000000;
	sram_mem[71561] = 16'b0000000000000000;
	sram_mem[71562] = 16'b0000000000000000;
	sram_mem[71563] = 16'b0000000000000000;
	sram_mem[71564] = 16'b0000000000000000;
	sram_mem[71565] = 16'b0000000000000000;
	sram_mem[71566] = 16'b0000000000000000;
	sram_mem[71567] = 16'b0000000000000000;
	sram_mem[71568] = 16'b0000000000000000;
	sram_mem[71569] = 16'b0000000000000000;
	sram_mem[71570] = 16'b0000000000000000;
	sram_mem[71571] = 16'b0000000000000000;
	sram_mem[71572] = 16'b0000000000000000;
	sram_mem[71573] = 16'b0000000000000000;
	sram_mem[71574] = 16'b0000000000000000;
	sram_mem[71575] = 16'b0000000000000000;
	sram_mem[71576] = 16'b0000000000000000;
	sram_mem[71577] = 16'b0000000000000000;
	sram_mem[71578] = 16'b0000000000000000;
	sram_mem[71579] = 16'b0000000000000000;
	sram_mem[71580] = 16'b0000000000000000;
	sram_mem[71581] = 16'b0000000000000000;
	sram_mem[71582] = 16'b0000000000000000;
	sram_mem[71583] = 16'b0000000000000000;
	sram_mem[71584] = 16'b0000000000000000;
	sram_mem[71585] = 16'b0000000000000000;
	sram_mem[71586] = 16'b0000000000000000;
	sram_mem[71587] = 16'b0000000000000000;
	sram_mem[71588] = 16'b0000000000000000;
	sram_mem[71589] = 16'b0000000000000000;
	sram_mem[71590] = 16'b0000000000000000;
	sram_mem[71591] = 16'b0000000000000000;
	sram_mem[71592] = 16'b0000000000000000;
	sram_mem[71593] = 16'b0000000000000000;
	sram_mem[71594] = 16'b0000000000000000;
	sram_mem[71595] = 16'b0000000000000000;
	sram_mem[71596] = 16'b0000000000000000;
	sram_mem[71597] = 16'b0000000000000000;
	sram_mem[71598] = 16'b0000000000000000;
	sram_mem[71599] = 16'b0000000000000000;
	sram_mem[71600] = 16'b0000000000000000;
	sram_mem[71601] = 16'b0000000000000000;
	sram_mem[71602] = 16'b0000000000000000;
	sram_mem[71603] = 16'b0000000000000000;
	sram_mem[71604] = 16'b0000000000000000;
	sram_mem[71605] = 16'b0000000000000000;
	sram_mem[71606] = 16'b0000000000000000;
	sram_mem[71607] = 16'b0000000000000000;
	sram_mem[71608] = 16'b0000000000000000;
	sram_mem[71609] = 16'b0000000000000000;
	sram_mem[71610] = 16'b0000000000000000;
	sram_mem[71611] = 16'b0000000000000000;
	sram_mem[71612] = 16'b0000000000000000;
	sram_mem[71613] = 16'b0000000000000000;
	sram_mem[71614] = 16'b0000000000000000;
	sram_mem[71615] = 16'b0000000000000000;
	sram_mem[71616] = 16'b0000000000000000;
	sram_mem[71617] = 16'b0000000000000000;
	sram_mem[71618] = 16'b0000000000000000;
	sram_mem[71619] = 16'b0000000000000000;
	sram_mem[71620] = 16'b0000000000000000;
	sram_mem[71621] = 16'b0000000000000000;
	sram_mem[71622] = 16'b0000000000000000;
	sram_mem[71623] = 16'b0000000000000000;
	sram_mem[71624] = 16'b0000000000000000;
	sram_mem[71625] = 16'b0000000000000000;
	sram_mem[71626] = 16'b0000000000000000;
	sram_mem[71627] = 16'b0000000000000000;
	sram_mem[71628] = 16'b0000000000000000;
	sram_mem[71629] = 16'b0000000000000000;
	sram_mem[71630] = 16'b0000000000000000;
	sram_mem[71631] = 16'b0000000000000000;
	sram_mem[71632] = 16'b0000000000000000;
	sram_mem[71633] = 16'b0000000000000000;
	sram_mem[71634] = 16'b0000000000000000;
	sram_mem[71635] = 16'b0000000000000000;
	sram_mem[71636] = 16'b0000000000000000;
	sram_mem[71637] = 16'b0000000000000000;
	sram_mem[71638] = 16'b0000000000000000;
	sram_mem[71639] = 16'b0000000000000000;
	sram_mem[71640] = 16'b0000000000000000;
	sram_mem[71641] = 16'b0000000000000000;
	sram_mem[71642] = 16'b0000000000000000;
	sram_mem[71643] = 16'b0000000000000000;
	sram_mem[71644] = 16'b0000000000000000;
	sram_mem[71645] = 16'b0000000000000000;
	sram_mem[71646] = 16'b0000000000000000;
	sram_mem[71647] = 16'b0000000000000000;
	sram_mem[71648] = 16'b0000000000000000;
	sram_mem[71649] = 16'b0000000000000000;
	sram_mem[71650] = 16'b0000000000000000;
	sram_mem[71651] = 16'b0000000000000000;
	sram_mem[71652] = 16'b0000000000000000;
	sram_mem[71653] = 16'b0000000000000000;
	sram_mem[71654] = 16'b0000000000000000;
	sram_mem[71655] = 16'b0000000000000000;
	sram_mem[71656] = 16'b0000000000000000;
	sram_mem[71657] = 16'b0000000000000000;
	sram_mem[71658] = 16'b0000000000000000;
	sram_mem[71659] = 16'b0000000000000000;
	sram_mem[71660] = 16'b0000000000000000;
	sram_mem[71661] = 16'b0000000000000000;
	sram_mem[71662] = 16'b0000000000000000;
	sram_mem[71663] = 16'b0000000000000000;
	sram_mem[71664] = 16'b0000000000000000;
	sram_mem[71665] = 16'b0000000000000000;
	sram_mem[71666] = 16'b0000000000000000;
	sram_mem[71667] = 16'b0000000000000000;
	sram_mem[71668] = 16'b0000000000000000;
	sram_mem[71669] = 16'b0000000000000000;
	sram_mem[71670] = 16'b0000000000000000;
	sram_mem[71671] = 16'b0000000000000000;
	sram_mem[71672] = 16'b0000000000000000;
	sram_mem[71673] = 16'b0000000000000000;
	sram_mem[71674] = 16'b0000000000000000;
	sram_mem[71675] = 16'b0000000000000000;
	sram_mem[71676] = 16'b0000000000000000;
	sram_mem[71677] = 16'b0000000000000000;
	sram_mem[71678] = 16'b0000000000000000;
	sram_mem[71679] = 16'b0000000000000000;
	sram_mem[71680] = 16'b0000000000000000;
	sram_mem[71681] = 16'b0000000000000000;
	sram_mem[71682] = 16'b0000000000000000;
	sram_mem[71683] = 16'b0000000000000000;
	sram_mem[71684] = 16'b0000000000000000;
	sram_mem[71685] = 16'b0000000000000000;
	sram_mem[71686] = 16'b0000000000000000;
	sram_mem[71687] = 16'b0000000000000000;
	sram_mem[71688] = 16'b0000000000000000;
	sram_mem[71689] = 16'b0000000000000000;
	sram_mem[71690] = 16'b0000000000000000;
	sram_mem[71691] = 16'b0000000000000000;
	sram_mem[71692] = 16'b0000000000000000;
	sram_mem[71693] = 16'b0000000000000000;
	sram_mem[71694] = 16'b0000000000000000;
	sram_mem[71695] = 16'b0000000000000000;
	sram_mem[71696] = 16'b0000000000000000;
	sram_mem[71697] = 16'b0000000000000000;
	sram_mem[71698] = 16'b0000000000000000;
	sram_mem[71699] = 16'b0000000000000000;
	sram_mem[71700] = 16'b0000000000000000;
	sram_mem[71701] = 16'b0000000000000000;
	sram_mem[71702] = 16'b0000000000000000;
	sram_mem[71703] = 16'b0000000000000000;
	sram_mem[71704] = 16'b0000000000000000;
	sram_mem[71705] = 16'b0000000000000000;
	sram_mem[71706] = 16'b0000000000000000;
	sram_mem[71707] = 16'b0000000000000000;
	sram_mem[71708] = 16'b0000000000000000;
	sram_mem[71709] = 16'b0000000000000000;
	sram_mem[71710] = 16'b0000000000000000;
	sram_mem[71711] = 16'b0000000000000000;
	sram_mem[71712] = 16'b0000000000000000;
	sram_mem[71713] = 16'b0000000000000000;
	sram_mem[71714] = 16'b0000000000000000;
	sram_mem[71715] = 16'b0000000000000000;
	sram_mem[71716] = 16'b0000000000000000;
	sram_mem[71717] = 16'b0000000000000000;
	sram_mem[71718] = 16'b0000000000000000;
	sram_mem[71719] = 16'b0000000000000000;
	sram_mem[71720] = 16'b0000000000000000;
	sram_mem[71721] = 16'b0000000000000000;
	sram_mem[71722] = 16'b0000000000000000;
	sram_mem[71723] = 16'b0000000000000000;
	sram_mem[71724] = 16'b0000000000000000;
	sram_mem[71725] = 16'b0000000000000000;
	sram_mem[71726] = 16'b0000000000000000;
	sram_mem[71727] = 16'b0000000000000000;
	sram_mem[71728] = 16'b0000000000000000;
	sram_mem[71729] = 16'b0000000000000000;
	sram_mem[71730] = 16'b0000000000000000;
	sram_mem[71731] = 16'b0000000000000000;
	sram_mem[71732] = 16'b0000000000000000;
	sram_mem[71733] = 16'b0000000000000000;
	sram_mem[71734] = 16'b0000000000000000;
	sram_mem[71735] = 16'b0000000000000000;
	sram_mem[71736] = 16'b0000000000000000;
	sram_mem[71737] = 16'b0000000000000000;
	sram_mem[71738] = 16'b0000000000000000;
	sram_mem[71739] = 16'b0000000000000000;
	sram_mem[71740] = 16'b0000000000000000;
	sram_mem[71741] = 16'b0000000000000000;
	sram_mem[71742] = 16'b0000000000000000;
	sram_mem[71743] = 16'b0000000000000000;
	sram_mem[71744] = 16'b0000000000000000;
	sram_mem[71745] = 16'b0000000000000000;
	sram_mem[71746] = 16'b0000000000000000;
	sram_mem[71747] = 16'b0000000000000000;
	sram_mem[71748] = 16'b0000000000000000;
	sram_mem[71749] = 16'b0000000000000000;
	sram_mem[71750] = 16'b0000000000000000;
	sram_mem[71751] = 16'b0000000000000000;
	sram_mem[71752] = 16'b0000000000000000;
	sram_mem[71753] = 16'b0000000000000000;
	sram_mem[71754] = 16'b0000000000000000;
	sram_mem[71755] = 16'b0000000000000000;
	sram_mem[71756] = 16'b0000000000000000;
	sram_mem[71757] = 16'b0000000000000000;
	sram_mem[71758] = 16'b0000000000000000;
	sram_mem[71759] = 16'b0000000000000000;
	sram_mem[71760] = 16'b0000000000000000;
	sram_mem[71761] = 16'b0000000000000000;
	sram_mem[71762] = 16'b0000000000000000;
	sram_mem[71763] = 16'b0000000000000000;
	sram_mem[71764] = 16'b0000000000000000;
	sram_mem[71765] = 16'b0000000000000000;
	sram_mem[71766] = 16'b0000000000000000;
	sram_mem[71767] = 16'b0000000000000000;
	sram_mem[71768] = 16'b0000000000000000;
	sram_mem[71769] = 16'b0000000000000000;
	sram_mem[71770] = 16'b0000000000000000;
	sram_mem[71771] = 16'b0000000000000000;
	sram_mem[71772] = 16'b0000000000000000;
	sram_mem[71773] = 16'b0000000000000000;
	sram_mem[71774] = 16'b0000000000000000;
	sram_mem[71775] = 16'b0000000000000000;
	sram_mem[71776] = 16'b0000000000000000;
	sram_mem[71777] = 16'b0000000000000000;
	sram_mem[71778] = 16'b0000000000000000;
	sram_mem[71779] = 16'b0000000000000000;
	sram_mem[71780] = 16'b0000000000000000;
	sram_mem[71781] = 16'b0000000000000000;
	sram_mem[71782] = 16'b0000000000000000;
	sram_mem[71783] = 16'b0000000000000000;
	sram_mem[71784] = 16'b0000000000000000;
	sram_mem[71785] = 16'b0000000000000000;
	sram_mem[71786] = 16'b0000000000000000;
	sram_mem[71787] = 16'b0000000000000000;
	sram_mem[71788] = 16'b0000000000000000;
	sram_mem[71789] = 16'b0000000000000000;
	sram_mem[71790] = 16'b0000000000000000;
	sram_mem[71791] = 16'b0000000000000000;
	sram_mem[71792] = 16'b0000000000000000;
	sram_mem[71793] = 16'b0000000000000000;
	sram_mem[71794] = 16'b0000000000000000;
	sram_mem[71795] = 16'b0000000000000000;
	sram_mem[71796] = 16'b0000000000000000;
	sram_mem[71797] = 16'b0000000000000000;
	sram_mem[71798] = 16'b0000000000000000;
	sram_mem[71799] = 16'b0000000000000000;
	sram_mem[71800] = 16'b0000000000000000;
	sram_mem[71801] = 16'b0000000000000000;
	sram_mem[71802] = 16'b0000000000000000;
	sram_mem[71803] = 16'b0000000000000000;
	sram_mem[71804] = 16'b0000000000000000;
	sram_mem[71805] = 16'b0000000000000000;
	sram_mem[71806] = 16'b0000000000000000;
	sram_mem[71807] = 16'b0000000000000000;
	sram_mem[71808] = 16'b0000000000000000;
	sram_mem[71809] = 16'b0000000000000000;
	sram_mem[71810] = 16'b0000000000000000;
	sram_mem[71811] = 16'b0000000000000000;
	sram_mem[71812] = 16'b0000000000000000;
	sram_mem[71813] = 16'b0000000000000000;
	sram_mem[71814] = 16'b0000000000000000;
	sram_mem[71815] = 16'b0000000000000000;
	sram_mem[71816] = 16'b0000000000000000;
	sram_mem[71817] = 16'b0000000000000000;
	sram_mem[71818] = 16'b0000000000000000;
	sram_mem[71819] = 16'b0000000000000000;
	sram_mem[71820] = 16'b0000000000000000;
	sram_mem[71821] = 16'b0000000000000000;
	sram_mem[71822] = 16'b0000000000000000;
	sram_mem[71823] = 16'b0000000000000000;
	sram_mem[71824] = 16'b0000000000000000;
	sram_mem[71825] = 16'b0000000000000000;
	sram_mem[71826] = 16'b0000000000000000;
	sram_mem[71827] = 16'b0000000000000000;
	sram_mem[71828] = 16'b0000000000000000;
	sram_mem[71829] = 16'b0000000000000000;
	sram_mem[71830] = 16'b0000000000000000;
	sram_mem[71831] = 16'b0000000000000000;
	sram_mem[71832] = 16'b0000000000000000;
	sram_mem[71833] = 16'b0000000000000000;
	sram_mem[71834] = 16'b0000000000000000;
	sram_mem[71835] = 16'b0000000000000000;
	sram_mem[71836] = 16'b0000000000000000;
	sram_mem[71837] = 16'b0000000000000000;
	sram_mem[71838] = 16'b0000000000000000;
	sram_mem[71839] = 16'b0000000000000000;
	sram_mem[71840] = 16'b0000000000000000;
	sram_mem[71841] = 16'b0000000000000000;
	sram_mem[71842] = 16'b0000000000000000;
	sram_mem[71843] = 16'b0000000000000000;
	sram_mem[71844] = 16'b0000000000000000;
	sram_mem[71845] = 16'b0000000000000000;
	sram_mem[71846] = 16'b0000000000000000;
	sram_mem[71847] = 16'b0000000000000000;
	sram_mem[71848] = 16'b0000000000000000;
	sram_mem[71849] = 16'b0000000000000000;
	sram_mem[71850] = 16'b0000000000000000;
	sram_mem[71851] = 16'b0000000000000000;
	sram_mem[71852] = 16'b0000000000000000;
	sram_mem[71853] = 16'b0000000000000000;
	sram_mem[71854] = 16'b0000000000000000;
	sram_mem[71855] = 16'b0000000000000000;
	sram_mem[71856] = 16'b0000000000000000;
	sram_mem[71857] = 16'b0000000000000000;
	sram_mem[71858] = 16'b0000000000000000;
	sram_mem[71859] = 16'b0000000000000000;
	sram_mem[71860] = 16'b0000000000000000;
	sram_mem[71861] = 16'b0000000000000000;
	sram_mem[71862] = 16'b0000000000000000;
	sram_mem[71863] = 16'b0000000000000000;
	sram_mem[71864] = 16'b0000000000000000;
	sram_mem[71865] = 16'b0000000000000000;
	sram_mem[71866] = 16'b0000000000000000;
	sram_mem[71867] = 16'b0000000000000000;
	sram_mem[71868] = 16'b0000000000000000;
	sram_mem[71869] = 16'b0000000000000000;
	sram_mem[71870] = 16'b0000000000000000;
	sram_mem[71871] = 16'b0000000000000000;
	sram_mem[71872] = 16'b0000000000000000;
	sram_mem[71873] = 16'b0000000000000000;
	sram_mem[71874] = 16'b0000000000000000;
	sram_mem[71875] = 16'b0000000000000000;
	sram_mem[71876] = 16'b0000000000000000;
	sram_mem[71877] = 16'b0000000000000000;
	sram_mem[71878] = 16'b0000000000000000;
	sram_mem[71879] = 16'b0000000000000000;
	sram_mem[71880] = 16'b0000000000000000;
	sram_mem[71881] = 16'b0000000000000000;
	sram_mem[71882] = 16'b0000000000000000;
	sram_mem[71883] = 16'b0000000000000000;
	sram_mem[71884] = 16'b0000000000000000;
	sram_mem[71885] = 16'b0000000000000000;
	sram_mem[71886] = 16'b0000000000000000;
	sram_mem[71887] = 16'b0000000000000000;
	sram_mem[71888] = 16'b0000000000000000;
	sram_mem[71889] = 16'b0000000000000000;
	sram_mem[71890] = 16'b0000000000000000;
	sram_mem[71891] = 16'b0000000000000000;
	sram_mem[71892] = 16'b0000000000000000;
	sram_mem[71893] = 16'b0000000000000000;
	sram_mem[71894] = 16'b0000000000000000;
	sram_mem[71895] = 16'b0000000000000000;
	sram_mem[71896] = 16'b0000000000000000;
	sram_mem[71897] = 16'b0000000000000000;
	sram_mem[71898] = 16'b0000000000000000;
	sram_mem[71899] = 16'b0000000000000000;
	sram_mem[71900] = 16'b0000000000000000;
	sram_mem[71901] = 16'b0000000000000000;
	sram_mem[71902] = 16'b0000000000000000;
	sram_mem[71903] = 16'b0000000000000000;
	sram_mem[71904] = 16'b0000000000000000;
	sram_mem[71905] = 16'b0000000000000000;
	sram_mem[71906] = 16'b0000000000000000;
	sram_mem[71907] = 16'b0000000000000000;
	sram_mem[71908] = 16'b0000000000000000;
	sram_mem[71909] = 16'b0000000000000000;
	sram_mem[71910] = 16'b0000000000000000;
	sram_mem[71911] = 16'b0000000000000000;
	sram_mem[71912] = 16'b0000000000000000;
	sram_mem[71913] = 16'b0000000000000000;
	sram_mem[71914] = 16'b0000000000000000;
	sram_mem[71915] = 16'b0000000000000000;
	sram_mem[71916] = 16'b0000000000000000;
	sram_mem[71917] = 16'b0000000000000000;
	sram_mem[71918] = 16'b0000000000000000;
	sram_mem[71919] = 16'b0000000000000000;
	sram_mem[71920] = 16'b0000000000000000;
	sram_mem[71921] = 16'b0000000000000000;
	sram_mem[71922] = 16'b0000000000000000;
	sram_mem[71923] = 16'b0000000000000000;
	sram_mem[71924] = 16'b0000000000000000;
	sram_mem[71925] = 16'b0000000000000000;
	sram_mem[71926] = 16'b0000000000000000;
	sram_mem[71927] = 16'b0000000000000000;
	sram_mem[71928] = 16'b0000000000000000;
	sram_mem[71929] = 16'b0000000000000000;
	sram_mem[71930] = 16'b0000000000000000;
	sram_mem[71931] = 16'b0000000000000000;
	sram_mem[71932] = 16'b0000000000000000;
	sram_mem[71933] = 16'b0000000000000000;
	sram_mem[71934] = 16'b0000000000000000;
	sram_mem[71935] = 16'b0000000000000000;
	sram_mem[71936] = 16'b0000000000000000;
	sram_mem[71937] = 16'b0000000000000000;
	sram_mem[71938] = 16'b0000000000000000;
	sram_mem[71939] = 16'b0000000000000000;
	sram_mem[71940] = 16'b0000000000000000;
	sram_mem[71941] = 16'b0000000000000000;
	sram_mem[71942] = 16'b0000000000000000;
	sram_mem[71943] = 16'b0000000000000000;
	sram_mem[71944] = 16'b0000000000000000;
	sram_mem[71945] = 16'b0000000000000000;
	sram_mem[71946] = 16'b0000000000000000;
	sram_mem[71947] = 16'b0000000000000000;
	sram_mem[71948] = 16'b0000000000000000;
	sram_mem[71949] = 16'b0000000000000000;
	sram_mem[71950] = 16'b0000000000000000;
	sram_mem[71951] = 16'b0000000000000000;
	sram_mem[71952] = 16'b0000000000000000;
	sram_mem[71953] = 16'b0000000000000000;
	sram_mem[71954] = 16'b0000000000000000;
	sram_mem[71955] = 16'b0000000000000000;
	sram_mem[71956] = 16'b0000000000000000;
	sram_mem[71957] = 16'b0000000000000000;
	sram_mem[71958] = 16'b0000000000000000;
	sram_mem[71959] = 16'b0000000000000000;
	sram_mem[71960] = 16'b0000000000000000;
	sram_mem[71961] = 16'b0000000000000000;
	sram_mem[71962] = 16'b0000000000000000;
	sram_mem[71963] = 16'b0000000000000000;
	sram_mem[71964] = 16'b0000000000000000;
	sram_mem[71965] = 16'b0000000000000000;
	sram_mem[71966] = 16'b0000000000000000;
	sram_mem[71967] = 16'b0000000000000000;
	sram_mem[71968] = 16'b0000000000000000;
	sram_mem[71969] = 16'b0000000000000000;
	sram_mem[71970] = 16'b0000000000000000;
	sram_mem[71971] = 16'b0000000000000000;
	sram_mem[71972] = 16'b0000000000000000;
	sram_mem[71973] = 16'b0000000000000000;
	sram_mem[71974] = 16'b0000000000000000;
	sram_mem[71975] = 16'b0000000000000000;
	sram_mem[71976] = 16'b0000000000000000;
	sram_mem[71977] = 16'b0000000000000000;
	sram_mem[71978] = 16'b0000000000000000;
	sram_mem[71979] = 16'b0000000000000000;
	sram_mem[71980] = 16'b0000000000000000;
	sram_mem[71981] = 16'b0000000000000000;
	sram_mem[71982] = 16'b0000000000000000;
	sram_mem[71983] = 16'b0000000000000000;
	sram_mem[71984] = 16'b0000000000000000;
	sram_mem[71985] = 16'b0000000000000000;
	sram_mem[71986] = 16'b0000000000000000;
	sram_mem[71987] = 16'b0000000000000000;
	sram_mem[71988] = 16'b0000000000000000;
	sram_mem[71989] = 16'b0000000000000000;
	sram_mem[71990] = 16'b0000000000000000;
	sram_mem[71991] = 16'b0000000000000000;
	sram_mem[71992] = 16'b0000000000000000;
	sram_mem[71993] = 16'b0000000000000000;
	sram_mem[71994] = 16'b0000000000000000;
	sram_mem[71995] = 16'b0000000000000000;
	sram_mem[71996] = 16'b0000000000000000;
	sram_mem[71997] = 16'b0000000000000000;
	sram_mem[71998] = 16'b0000000000000000;
	sram_mem[71999] = 16'b0000000000000000;
	sram_mem[72000] = 16'b0000000000000000;
	sram_mem[72001] = 16'b0000000000000000;
	sram_mem[72002] = 16'b0000000000000000;
	sram_mem[72003] = 16'b0000000000000000;
	sram_mem[72004] = 16'b0000000000000000;
	sram_mem[72005] = 16'b0000000000000000;
	sram_mem[72006] = 16'b0000000000000000;
	sram_mem[72007] = 16'b0000000000000000;
	sram_mem[72008] = 16'b0000000000000000;
	sram_mem[72009] = 16'b0000000000000000;
	sram_mem[72010] = 16'b0000000000000000;
	sram_mem[72011] = 16'b0000000000000000;
	sram_mem[72012] = 16'b0000000000000000;
	sram_mem[72013] = 16'b0000000000000000;
	sram_mem[72014] = 16'b0000000000000000;
	sram_mem[72015] = 16'b0000000000000000;
	sram_mem[72016] = 16'b0000000000000000;
	sram_mem[72017] = 16'b0000000000000000;
	sram_mem[72018] = 16'b0000000000000000;
	sram_mem[72019] = 16'b0000000000000000;
	sram_mem[72020] = 16'b0000000000000000;
	sram_mem[72021] = 16'b0000000000000000;
	sram_mem[72022] = 16'b0000000000000000;
	sram_mem[72023] = 16'b0000000000000000;
	sram_mem[72024] = 16'b0000000000000000;
	sram_mem[72025] = 16'b0000000000000000;
	sram_mem[72026] = 16'b0000000000000000;
	sram_mem[72027] = 16'b0000000000000000;
	sram_mem[72028] = 16'b0000000000000000;
	sram_mem[72029] = 16'b0000000000000000;
	sram_mem[72030] = 16'b0000000000000000;
	sram_mem[72031] = 16'b0000000000000000;
	sram_mem[72032] = 16'b0000000000000000;
	sram_mem[72033] = 16'b0000000000000000;
	sram_mem[72034] = 16'b0000000000000000;
	sram_mem[72035] = 16'b0000000000000000;
	sram_mem[72036] = 16'b0000000000000000;
	sram_mem[72037] = 16'b0000000000000000;
	sram_mem[72038] = 16'b0000000000000000;
	sram_mem[72039] = 16'b0000000000000000;
	sram_mem[72040] = 16'b0000000000000000;
	sram_mem[72041] = 16'b0000000000000000;
	sram_mem[72042] = 16'b0000000000000000;
	sram_mem[72043] = 16'b0000000000000000;
	sram_mem[72044] = 16'b0000000000000000;
	sram_mem[72045] = 16'b0000000000000000;
	sram_mem[72046] = 16'b0000000000000000;
	sram_mem[72047] = 16'b0000000000000000;
	sram_mem[72048] = 16'b0000000000000000;
	sram_mem[72049] = 16'b0000000000000000;
	sram_mem[72050] = 16'b0000000000000000;
	sram_mem[72051] = 16'b0000000000000000;
	sram_mem[72052] = 16'b0000000000000000;
	sram_mem[72053] = 16'b0000000000000000;
	sram_mem[72054] = 16'b0000000000000000;
	sram_mem[72055] = 16'b0000000000000000;
	sram_mem[72056] = 16'b0000000000000000;
	sram_mem[72057] = 16'b0000000000000000;
	sram_mem[72058] = 16'b0000000000000000;
	sram_mem[72059] = 16'b0000000000000000;
	sram_mem[72060] = 16'b0000000000000000;
	sram_mem[72061] = 16'b0000000000000000;
	sram_mem[72062] = 16'b0000000000000000;
	sram_mem[72063] = 16'b0000000000000000;
	sram_mem[72064] = 16'b0000000000000000;
	sram_mem[72065] = 16'b0000000000000000;
	sram_mem[72066] = 16'b0000000000000000;
	sram_mem[72067] = 16'b0000000000000000;
	sram_mem[72068] = 16'b0000000000000000;
	sram_mem[72069] = 16'b0000000000000000;
	sram_mem[72070] = 16'b0000000000000000;
	sram_mem[72071] = 16'b0000000000000000;
	sram_mem[72072] = 16'b0000000000000000;
	sram_mem[72073] = 16'b0000000000000000;
	sram_mem[72074] = 16'b0000000000000000;
	sram_mem[72075] = 16'b0000000000000000;
	sram_mem[72076] = 16'b0000000000000000;
	sram_mem[72077] = 16'b0000000000000000;
	sram_mem[72078] = 16'b0000000000000000;
	sram_mem[72079] = 16'b0000000000000000;
	sram_mem[72080] = 16'b0000000000000000;
	sram_mem[72081] = 16'b0000000000000000;
	sram_mem[72082] = 16'b0000000000000000;
	sram_mem[72083] = 16'b0000000000000000;
	sram_mem[72084] = 16'b0000000000000000;
	sram_mem[72085] = 16'b0000000000000000;
	sram_mem[72086] = 16'b0000000000000000;
	sram_mem[72087] = 16'b0000000000000000;
	sram_mem[72088] = 16'b0000000000000000;
	sram_mem[72089] = 16'b0000000000000000;
	sram_mem[72090] = 16'b0000000000000000;
	sram_mem[72091] = 16'b0000000000000000;
	sram_mem[72092] = 16'b0000000000000000;
	sram_mem[72093] = 16'b0000000000000000;
	sram_mem[72094] = 16'b0000000000000000;
	sram_mem[72095] = 16'b0000000000000000;
	sram_mem[72096] = 16'b0000000000000000;
	sram_mem[72097] = 16'b0000000000000000;
	sram_mem[72098] = 16'b0000000000000000;
	sram_mem[72099] = 16'b0000000000000000;
	sram_mem[72100] = 16'b0000000000000000;
	sram_mem[72101] = 16'b0000000000000000;
	sram_mem[72102] = 16'b0000000000000000;
	sram_mem[72103] = 16'b0000000000000000;
	sram_mem[72104] = 16'b0000000000000000;
	sram_mem[72105] = 16'b0000000000000000;
	sram_mem[72106] = 16'b0000000000000000;
	sram_mem[72107] = 16'b0000000000000000;
	sram_mem[72108] = 16'b0000000000000000;
	sram_mem[72109] = 16'b0000000000000000;
	sram_mem[72110] = 16'b0000000000000000;
	sram_mem[72111] = 16'b0000000000000000;
	sram_mem[72112] = 16'b0000000000000000;
	sram_mem[72113] = 16'b0000000000000000;
	sram_mem[72114] = 16'b0000000000000000;
	sram_mem[72115] = 16'b0000000000000000;
	sram_mem[72116] = 16'b0000000000000000;
	sram_mem[72117] = 16'b0000000000000000;
	sram_mem[72118] = 16'b0000000000000000;
	sram_mem[72119] = 16'b0000000000000000;
	sram_mem[72120] = 16'b0000000000000000;
	sram_mem[72121] = 16'b0000000000000000;
	sram_mem[72122] = 16'b0000000000000000;
	sram_mem[72123] = 16'b0000000000000000;
	sram_mem[72124] = 16'b0000000000000000;
	sram_mem[72125] = 16'b0000000000000000;
	sram_mem[72126] = 16'b0000000000000000;
	sram_mem[72127] = 16'b0000000000000000;
	sram_mem[72128] = 16'b0000000000000000;
	sram_mem[72129] = 16'b0000000000000000;
	sram_mem[72130] = 16'b0000000000000000;
	sram_mem[72131] = 16'b0000000000000000;
	sram_mem[72132] = 16'b0000000000000000;
	sram_mem[72133] = 16'b0000000000000000;
	sram_mem[72134] = 16'b0000000000000000;
	sram_mem[72135] = 16'b0000000000000000;
	sram_mem[72136] = 16'b0000000000000000;
	sram_mem[72137] = 16'b0000000000000000;
	sram_mem[72138] = 16'b0000000000000000;
	sram_mem[72139] = 16'b0000000000000000;
	sram_mem[72140] = 16'b0000000000000000;
	sram_mem[72141] = 16'b0000000000000000;
	sram_mem[72142] = 16'b0000000000000000;
	sram_mem[72143] = 16'b0000000000000000;
	sram_mem[72144] = 16'b0000000000000000;
	sram_mem[72145] = 16'b0000000000000000;
	sram_mem[72146] = 16'b0000000000000000;
	sram_mem[72147] = 16'b0000000000000000;
	sram_mem[72148] = 16'b0000000000000000;
	sram_mem[72149] = 16'b0000000000000000;
	sram_mem[72150] = 16'b0000000000000000;
	sram_mem[72151] = 16'b0000000000000000;
	sram_mem[72152] = 16'b0000000000000000;
	sram_mem[72153] = 16'b0000000000000000;
	sram_mem[72154] = 16'b0000000000000000;
	sram_mem[72155] = 16'b0000000000000000;
	sram_mem[72156] = 16'b0000000000000000;
	sram_mem[72157] = 16'b0000000000000000;
	sram_mem[72158] = 16'b0000000000000000;
	sram_mem[72159] = 16'b0000000000000000;
	sram_mem[72160] = 16'b0000000000000000;
	sram_mem[72161] = 16'b0000000000000000;
	sram_mem[72162] = 16'b0000000000000000;
	sram_mem[72163] = 16'b0000000000000000;
	sram_mem[72164] = 16'b0000000000000000;
	sram_mem[72165] = 16'b0000000000000000;
	sram_mem[72166] = 16'b0000000000000000;
	sram_mem[72167] = 16'b0000000000000000;
	sram_mem[72168] = 16'b0000000000000000;
	sram_mem[72169] = 16'b0000000000000000;
	sram_mem[72170] = 16'b0000000000000000;
	sram_mem[72171] = 16'b0000000000000000;
	sram_mem[72172] = 16'b0000000000000000;
	sram_mem[72173] = 16'b0000000000000000;
	sram_mem[72174] = 16'b0000000000000000;
	sram_mem[72175] = 16'b0000000000000000;
	sram_mem[72176] = 16'b0000000000000000;
	sram_mem[72177] = 16'b0000000000000000;
	sram_mem[72178] = 16'b0000000000000000;
	sram_mem[72179] = 16'b0000000000000000;
	sram_mem[72180] = 16'b0000000000000000;
	sram_mem[72181] = 16'b0000000000000000;
	sram_mem[72182] = 16'b0000000000000000;
	sram_mem[72183] = 16'b0000000000000000;
	sram_mem[72184] = 16'b0000000000000000;
	sram_mem[72185] = 16'b0000000000000000;
	sram_mem[72186] = 16'b0000000000000000;
	sram_mem[72187] = 16'b0000000000000000;
	sram_mem[72188] = 16'b0000000000000000;
	sram_mem[72189] = 16'b0000000000000000;
	sram_mem[72190] = 16'b0000000000000000;
	sram_mem[72191] = 16'b0000000000000000;
	sram_mem[72192] = 16'b0000000000000000;
	sram_mem[72193] = 16'b0000000000000000;
	sram_mem[72194] = 16'b0000000000000000;
	sram_mem[72195] = 16'b0000000000000000;
	sram_mem[72196] = 16'b0000000000000000;
	sram_mem[72197] = 16'b0000000000000000;
	sram_mem[72198] = 16'b0000000000000000;
	sram_mem[72199] = 16'b0000000000000000;
	sram_mem[72200] = 16'b0000000000000000;
	sram_mem[72201] = 16'b0000000000000000;
	sram_mem[72202] = 16'b0000000000000000;
	sram_mem[72203] = 16'b0000000000000000;
	sram_mem[72204] = 16'b0000000000000000;
	sram_mem[72205] = 16'b0000000000000000;
	sram_mem[72206] = 16'b0000000000000000;
	sram_mem[72207] = 16'b0000000000000000;
	sram_mem[72208] = 16'b0000000000000000;
	sram_mem[72209] = 16'b0000000000000000;
	sram_mem[72210] = 16'b0000000000000000;
	sram_mem[72211] = 16'b0000000000000000;
	sram_mem[72212] = 16'b0000000000000000;
	sram_mem[72213] = 16'b0000000000000000;
	sram_mem[72214] = 16'b0000000000000000;
	sram_mem[72215] = 16'b0000000000000000;
	sram_mem[72216] = 16'b0000000000000000;
	sram_mem[72217] = 16'b0000000000000000;
	sram_mem[72218] = 16'b0000000000000000;
	sram_mem[72219] = 16'b0000000000000000;
	sram_mem[72220] = 16'b0000000000000000;
	sram_mem[72221] = 16'b0000000000000000;
	sram_mem[72222] = 16'b0000000000000000;
	sram_mem[72223] = 16'b0000000000000000;
	sram_mem[72224] = 16'b0000000000000000;
	sram_mem[72225] = 16'b0000000000000000;
	sram_mem[72226] = 16'b0000000000000000;
	sram_mem[72227] = 16'b0000000000000000;
	sram_mem[72228] = 16'b0000000000000000;
	sram_mem[72229] = 16'b0000000000000000;
	sram_mem[72230] = 16'b0000000000000000;
	sram_mem[72231] = 16'b0000000000000000;
	sram_mem[72232] = 16'b0000000000000000;
	sram_mem[72233] = 16'b0000000000000000;
	sram_mem[72234] = 16'b0000000000000000;
	sram_mem[72235] = 16'b0000000000000000;
	sram_mem[72236] = 16'b0000000000000000;
	sram_mem[72237] = 16'b0000000000000000;
	sram_mem[72238] = 16'b0000000000000000;
	sram_mem[72239] = 16'b0000000000000000;
	sram_mem[72240] = 16'b0000000000000000;
	sram_mem[72241] = 16'b0000000000000000;
	sram_mem[72242] = 16'b0000000000000000;
	sram_mem[72243] = 16'b0000000000000000;
	sram_mem[72244] = 16'b0000000000000000;
	sram_mem[72245] = 16'b0000000000000000;
	sram_mem[72246] = 16'b0000000000000000;
	sram_mem[72247] = 16'b0000000000000000;
	sram_mem[72248] = 16'b0000000000000000;
	sram_mem[72249] = 16'b0000000000000000;
	sram_mem[72250] = 16'b0000000000000000;
	sram_mem[72251] = 16'b0000000000000000;
	sram_mem[72252] = 16'b0000000000000000;
	sram_mem[72253] = 16'b0000000000000000;
	sram_mem[72254] = 16'b0000000000000000;
	sram_mem[72255] = 16'b0000000000000000;
	sram_mem[72256] = 16'b0000000000000000;
	sram_mem[72257] = 16'b0000000000000000;
	sram_mem[72258] = 16'b0000000000000000;
	sram_mem[72259] = 16'b0000000000000000;
	sram_mem[72260] = 16'b0000000000000000;
	sram_mem[72261] = 16'b0000000000000000;
	sram_mem[72262] = 16'b0000000000000000;
	sram_mem[72263] = 16'b0000000000000000;
	sram_mem[72264] = 16'b0000000000000000;
	sram_mem[72265] = 16'b0000000000000000;
	sram_mem[72266] = 16'b0000000000000000;
	sram_mem[72267] = 16'b0000000000000000;
	sram_mem[72268] = 16'b0000000000000000;
	sram_mem[72269] = 16'b0000000000000000;
	sram_mem[72270] = 16'b0000000000000000;
	sram_mem[72271] = 16'b0000000000000000;
	sram_mem[72272] = 16'b0000000000000000;
	sram_mem[72273] = 16'b0000000000000000;
	sram_mem[72274] = 16'b0000000000000000;
	sram_mem[72275] = 16'b0000000000000000;
	sram_mem[72276] = 16'b0000000000000000;
	sram_mem[72277] = 16'b0000000000000000;
	sram_mem[72278] = 16'b0000000000000000;
	sram_mem[72279] = 16'b0000000000000000;
	sram_mem[72280] = 16'b0000000000000000;
	sram_mem[72281] = 16'b0000000000000000;
	sram_mem[72282] = 16'b0000000000000000;
	sram_mem[72283] = 16'b0000000000000000;
	sram_mem[72284] = 16'b0000000000000000;
	sram_mem[72285] = 16'b0000000000000000;
	sram_mem[72286] = 16'b0000000000000000;
	sram_mem[72287] = 16'b0000000000000000;
	sram_mem[72288] = 16'b0000000000000000;
	sram_mem[72289] = 16'b0000000000000000;
	sram_mem[72290] = 16'b0000000000000000;
	sram_mem[72291] = 16'b0000000000000000;
	sram_mem[72292] = 16'b0000000000000000;
	sram_mem[72293] = 16'b0000000000000000;
	sram_mem[72294] = 16'b0000000000000000;
	sram_mem[72295] = 16'b0000000000000000;
	sram_mem[72296] = 16'b0000000000000000;
	sram_mem[72297] = 16'b0000000000000000;
	sram_mem[72298] = 16'b0000000000000000;
	sram_mem[72299] = 16'b0000000000000000;
	sram_mem[72300] = 16'b0000000000000000;
	sram_mem[72301] = 16'b0000000000000000;
	sram_mem[72302] = 16'b0000000000000000;
	sram_mem[72303] = 16'b0000000000000000;
	sram_mem[72304] = 16'b0000000000000000;
	sram_mem[72305] = 16'b0000000000000000;
	sram_mem[72306] = 16'b0000000000000000;
	sram_mem[72307] = 16'b0000000000000000;
	sram_mem[72308] = 16'b0000000000000000;
	sram_mem[72309] = 16'b0000000000000000;
	sram_mem[72310] = 16'b0000000000000000;
	sram_mem[72311] = 16'b0000000000000000;
	sram_mem[72312] = 16'b0000000000000000;
	sram_mem[72313] = 16'b0000000000000000;
	sram_mem[72314] = 16'b0000000000000000;
	sram_mem[72315] = 16'b0000000000000000;
	sram_mem[72316] = 16'b0000000000000000;
	sram_mem[72317] = 16'b0000000000000000;
	sram_mem[72318] = 16'b0000000000000000;
	sram_mem[72319] = 16'b0000000000000000;
	sram_mem[72320] = 16'b0000000000000000;
	sram_mem[72321] = 16'b0000000000000000;
	sram_mem[72322] = 16'b0000000000000000;
	sram_mem[72323] = 16'b0000000000000000;
	sram_mem[72324] = 16'b0000000000000000;
	sram_mem[72325] = 16'b0000000000000000;
	sram_mem[72326] = 16'b0000000000000000;
	sram_mem[72327] = 16'b0000000000000000;
	sram_mem[72328] = 16'b0000000000000000;
	sram_mem[72329] = 16'b0000000000000000;
	sram_mem[72330] = 16'b0000000000000000;
	sram_mem[72331] = 16'b0000000000000000;
	sram_mem[72332] = 16'b0000000000000000;
	sram_mem[72333] = 16'b0000000000000000;
	sram_mem[72334] = 16'b0000000000000000;
	sram_mem[72335] = 16'b0000000000000000;
	sram_mem[72336] = 16'b0000000000000000;
	sram_mem[72337] = 16'b0000000000000000;
	sram_mem[72338] = 16'b0000000000000000;
	sram_mem[72339] = 16'b0000000000000000;
	sram_mem[72340] = 16'b0000000000000000;
	sram_mem[72341] = 16'b0000000000000000;
	sram_mem[72342] = 16'b0000000000000000;
	sram_mem[72343] = 16'b0000000000000000;
	sram_mem[72344] = 16'b0000000000000000;
	sram_mem[72345] = 16'b0000000000000000;
	sram_mem[72346] = 16'b0000000000000000;
	sram_mem[72347] = 16'b0000000000000000;
	sram_mem[72348] = 16'b0000000000000000;
	sram_mem[72349] = 16'b0000000000000000;
	sram_mem[72350] = 16'b0000000000000000;
	sram_mem[72351] = 16'b0000000000000000;
	sram_mem[72352] = 16'b0000000000000000;
	sram_mem[72353] = 16'b0000000000000000;
	sram_mem[72354] = 16'b0000000000000000;
	sram_mem[72355] = 16'b0000000000000000;
	sram_mem[72356] = 16'b0000000000000000;
	sram_mem[72357] = 16'b0000000000000000;
	sram_mem[72358] = 16'b0000000000000000;
	sram_mem[72359] = 16'b0000000000000000;
	sram_mem[72360] = 16'b0000000000000000;
	sram_mem[72361] = 16'b0000000000000000;
	sram_mem[72362] = 16'b0000000000000000;
	sram_mem[72363] = 16'b0000000000000000;
	sram_mem[72364] = 16'b0000000000000000;
	sram_mem[72365] = 16'b0000000000000000;
	sram_mem[72366] = 16'b0000000000000000;
	sram_mem[72367] = 16'b0000000000000000;
	sram_mem[72368] = 16'b0000000000000000;
	sram_mem[72369] = 16'b0000000000000000;
	sram_mem[72370] = 16'b0000000000000000;
	sram_mem[72371] = 16'b0000000000000000;
	sram_mem[72372] = 16'b0000000000000000;
	sram_mem[72373] = 16'b0000000000000000;
	sram_mem[72374] = 16'b0000000000000000;
	sram_mem[72375] = 16'b0000000000000000;
	sram_mem[72376] = 16'b0000000000000000;
	sram_mem[72377] = 16'b0000000000000000;
	sram_mem[72378] = 16'b0000000000000000;
	sram_mem[72379] = 16'b0000000000000000;
	sram_mem[72380] = 16'b0000000000000000;
	sram_mem[72381] = 16'b0000000000000000;
	sram_mem[72382] = 16'b0000000000000000;
	sram_mem[72383] = 16'b0000000000000000;
	sram_mem[72384] = 16'b0000000000000000;
	sram_mem[72385] = 16'b0000000000000000;
	sram_mem[72386] = 16'b0000000000000000;
	sram_mem[72387] = 16'b0000000000000000;
	sram_mem[72388] = 16'b0000000000000000;
	sram_mem[72389] = 16'b0000000000000000;
	sram_mem[72390] = 16'b0000000000000000;
	sram_mem[72391] = 16'b0000000000000000;
	sram_mem[72392] = 16'b0000000000000000;
	sram_mem[72393] = 16'b0000000000000000;
	sram_mem[72394] = 16'b0000000000000000;
	sram_mem[72395] = 16'b0000000000000000;
	sram_mem[72396] = 16'b0000000000000000;
	sram_mem[72397] = 16'b0000000000000000;
	sram_mem[72398] = 16'b0000000000000000;
	sram_mem[72399] = 16'b0000000000000000;
	sram_mem[72400] = 16'b0000000000000000;
	sram_mem[72401] = 16'b0000000000000000;
	sram_mem[72402] = 16'b0000000000000000;
	sram_mem[72403] = 16'b0000000000000000;
	sram_mem[72404] = 16'b0000000000000000;
	sram_mem[72405] = 16'b0000000000000000;
	sram_mem[72406] = 16'b0000000000000000;
	sram_mem[72407] = 16'b0000000000000000;
	sram_mem[72408] = 16'b0000000000000000;
	sram_mem[72409] = 16'b0000000000000000;
	sram_mem[72410] = 16'b0000000000000000;
	sram_mem[72411] = 16'b0000000000000000;
	sram_mem[72412] = 16'b0000000000000000;
	sram_mem[72413] = 16'b0000000000000000;
	sram_mem[72414] = 16'b0000000000000000;
	sram_mem[72415] = 16'b0000000000000000;
	sram_mem[72416] = 16'b0000000000000000;
	sram_mem[72417] = 16'b0000000000000000;
	sram_mem[72418] = 16'b0000000000000000;
	sram_mem[72419] = 16'b0000000000000000;
	sram_mem[72420] = 16'b0000000000000000;
	sram_mem[72421] = 16'b0000000000000000;
	sram_mem[72422] = 16'b0000000000000000;
	sram_mem[72423] = 16'b0000000000000000;
	sram_mem[72424] = 16'b0000000000000000;
	sram_mem[72425] = 16'b0000000000000000;
	sram_mem[72426] = 16'b0000000000000000;
	sram_mem[72427] = 16'b0000000000000000;
	sram_mem[72428] = 16'b0000000000000000;
	sram_mem[72429] = 16'b0000000000000000;
	sram_mem[72430] = 16'b0000000000000000;
	sram_mem[72431] = 16'b0000000000000000;
	sram_mem[72432] = 16'b0000000000000000;
	sram_mem[72433] = 16'b0000000000000000;
	sram_mem[72434] = 16'b0000000000000000;
	sram_mem[72435] = 16'b0000000000000000;
	sram_mem[72436] = 16'b0000000000000000;
	sram_mem[72437] = 16'b0000000000000000;
	sram_mem[72438] = 16'b0000000000000000;
	sram_mem[72439] = 16'b0000000000000000;
	sram_mem[72440] = 16'b0000000000000000;
	sram_mem[72441] = 16'b0000000000000000;
	sram_mem[72442] = 16'b0000000000000000;
	sram_mem[72443] = 16'b0000000000000000;
	sram_mem[72444] = 16'b0000000000000000;
	sram_mem[72445] = 16'b0000000000000000;
	sram_mem[72446] = 16'b0000000000000000;
	sram_mem[72447] = 16'b0000000000000000;
	sram_mem[72448] = 16'b0000000000000000;
	sram_mem[72449] = 16'b0000000000000000;
	sram_mem[72450] = 16'b0000000000000000;
	sram_mem[72451] = 16'b0000000000000000;
	sram_mem[72452] = 16'b0000000000000000;
	sram_mem[72453] = 16'b0000000000000000;
	sram_mem[72454] = 16'b0000000000000000;
	sram_mem[72455] = 16'b0000000000000000;
	sram_mem[72456] = 16'b0000000000000000;
	sram_mem[72457] = 16'b0000000000000000;
	sram_mem[72458] = 16'b0000000000000000;
	sram_mem[72459] = 16'b0000000000000000;
	sram_mem[72460] = 16'b0000000000000000;
	sram_mem[72461] = 16'b0000000000000000;
	sram_mem[72462] = 16'b0000000000000000;
	sram_mem[72463] = 16'b0000000000000000;
	sram_mem[72464] = 16'b0000000000000000;
	sram_mem[72465] = 16'b0000000000000000;
	sram_mem[72466] = 16'b0000000000000000;
	sram_mem[72467] = 16'b0000000000000000;
	sram_mem[72468] = 16'b0000000000000000;
	sram_mem[72469] = 16'b0000000000000000;
	sram_mem[72470] = 16'b0000000000000000;
	sram_mem[72471] = 16'b0000000000000000;
	sram_mem[72472] = 16'b0000000000000000;
	sram_mem[72473] = 16'b0000000000000000;
	sram_mem[72474] = 16'b0000000000000000;
	sram_mem[72475] = 16'b0000000000000000;
	sram_mem[72476] = 16'b0000000000000000;
	sram_mem[72477] = 16'b0000000000000000;
	sram_mem[72478] = 16'b0000000000000000;
	sram_mem[72479] = 16'b0000000000000000;
	sram_mem[72480] = 16'b0000000000000000;
	sram_mem[72481] = 16'b0000000000000000;
	sram_mem[72482] = 16'b0000000000000000;
	sram_mem[72483] = 16'b0000000000000000;
	sram_mem[72484] = 16'b0000000000000000;
	sram_mem[72485] = 16'b0000000000000000;
	sram_mem[72486] = 16'b0000000000000000;
	sram_mem[72487] = 16'b0000000000000000;
	sram_mem[72488] = 16'b0000000000000000;
	sram_mem[72489] = 16'b0000000000000000;
	sram_mem[72490] = 16'b0000000000000000;
	sram_mem[72491] = 16'b0000000000000000;
	sram_mem[72492] = 16'b0000000000000000;
	sram_mem[72493] = 16'b0000000000000000;
	sram_mem[72494] = 16'b0000000000000000;
	sram_mem[72495] = 16'b0000000000000000;
	sram_mem[72496] = 16'b0000000000000000;
	sram_mem[72497] = 16'b0000000000000000;
	sram_mem[72498] = 16'b0000000000000000;
	sram_mem[72499] = 16'b0000000000000000;
	sram_mem[72500] = 16'b0000000000000000;
	sram_mem[72501] = 16'b0000000000000000;
	sram_mem[72502] = 16'b0000000000000000;
	sram_mem[72503] = 16'b0000000000000000;
	sram_mem[72504] = 16'b0000000000000000;
	sram_mem[72505] = 16'b0000000000000000;
	sram_mem[72506] = 16'b0000000000000000;
	sram_mem[72507] = 16'b0000000000000000;
	sram_mem[72508] = 16'b0000000000000000;
	sram_mem[72509] = 16'b0000000000000000;
	sram_mem[72510] = 16'b0000000000000000;
	sram_mem[72511] = 16'b0000000000000000;
	sram_mem[72512] = 16'b0000000000000000;
	sram_mem[72513] = 16'b0000000000000000;
	sram_mem[72514] = 16'b0000000000000000;
	sram_mem[72515] = 16'b0000000000000000;
	sram_mem[72516] = 16'b0000000000000000;
	sram_mem[72517] = 16'b0000000000000000;
	sram_mem[72518] = 16'b0000000000000000;
	sram_mem[72519] = 16'b0000000000000000;
	sram_mem[72520] = 16'b0000000000000000;
	sram_mem[72521] = 16'b0000000000000000;
	sram_mem[72522] = 16'b0000000000000000;
	sram_mem[72523] = 16'b0000000000000000;
	sram_mem[72524] = 16'b0000000000000000;
	sram_mem[72525] = 16'b0000000000000000;
	sram_mem[72526] = 16'b0000000000000000;
	sram_mem[72527] = 16'b0000000000000000;
	sram_mem[72528] = 16'b0000000000000000;
	sram_mem[72529] = 16'b0000000000000000;
	sram_mem[72530] = 16'b0000000000000000;
	sram_mem[72531] = 16'b0000000000000000;
	sram_mem[72532] = 16'b0000000000000000;
	sram_mem[72533] = 16'b0000000000000000;
	sram_mem[72534] = 16'b0000000000000000;
	sram_mem[72535] = 16'b0000000000000000;
	sram_mem[72536] = 16'b0000000000000000;
	sram_mem[72537] = 16'b0000000000000000;
	sram_mem[72538] = 16'b0000000000000000;
	sram_mem[72539] = 16'b0000000000000000;
	sram_mem[72540] = 16'b0000000000000000;
	sram_mem[72541] = 16'b0000000000000000;
	sram_mem[72542] = 16'b0000000000000000;
	sram_mem[72543] = 16'b0000000000000000;
	sram_mem[72544] = 16'b0000000000000000;
	sram_mem[72545] = 16'b0000000000000000;
	sram_mem[72546] = 16'b0000000000000000;
	sram_mem[72547] = 16'b0000000000000000;
	sram_mem[72548] = 16'b0000000000000000;
	sram_mem[72549] = 16'b0000000000000000;
	sram_mem[72550] = 16'b0000000000000000;
	sram_mem[72551] = 16'b0000000000000000;
	sram_mem[72552] = 16'b0000000000000000;
	sram_mem[72553] = 16'b0000000000000000;
	sram_mem[72554] = 16'b0000000000000000;
	sram_mem[72555] = 16'b0000000000000000;
	sram_mem[72556] = 16'b0000000000000000;
	sram_mem[72557] = 16'b0000000000000000;
	sram_mem[72558] = 16'b0000000000000000;
	sram_mem[72559] = 16'b0000000000000000;
	sram_mem[72560] = 16'b0000000000000000;
	sram_mem[72561] = 16'b0000000000000000;
	sram_mem[72562] = 16'b0000000000000000;
	sram_mem[72563] = 16'b0000000000000000;
	sram_mem[72564] = 16'b0000000000000000;
	sram_mem[72565] = 16'b0000000000000000;
	sram_mem[72566] = 16'b0000000000000000;
	sram_mem[72567] = 16'b0000000000000000;
	sram_mem[72568] = 16'b0000000000000000;
	sram_mem[72569] = 16'b0000000000000000;
	sram_mem[72570] = 16'b0000000000000000;
	sram_mem[72571] = 16'b0000000000000000;
	sram_mem[72572] = 16'b0000000000000000;
	sram_mem[72573] = 16'b0000000000000000;
	sram_mem[72574] = 16'b0000000000000000;
	sram_mem[72575] = 16'b0000000000000000;
	sram_mem[72576] = 16'b0000000000000000;
	sram_mem[72577] = 16'b0000000000000000;
	sram_mem[72578] = 16'b0000000000000000;
	sram_mem[72579] = 16'b0000000000000000;
	sram_mem[72580] = 16'b0000000000000000;
	sram_mem[72581] = 16'b0000000000000000;
	sram_mem[72582] = 16'b0000000000000000;
	sram_mem[72583] = 16'b0000000000000000;
	sram_mem[72584] = 16'b0000000000000000;
	sram_mem[72585] = 16'b0000000000000000;
	sram_mem[72586] = 16'b0000000000000000;
	sram_mem[72587] = 16'b0000000000000000;
	sram_mem[72588] = 16'b0000000000000000;
	sram_mem[72589] = 16'b0000000000000000;
	sram_mem[72590] = 16'b0000000000000000;
	sram_mem[72591] = 16'b0000000000000000;
	sram_mem[72592] = 16'b0000000000000000;
	sram_mem[72593] = 16'b0000000000000000;
	sram_mem[72594] = 16'b0000000000000000;
	sram_mem[72595] = 16'b0000000000000000;
	sram_mem[72596] = 16'b0000000000000000;
	sram_mem[72597] = 16'b0000000000000000;
	sram_mem[72598] = 16'b0000000000000000;
	sram_mem[72599] = 16'b0000000000000000;
	sram_mem[72600] = 16'b0000000000000000;
	sram_mem[72601] = 16'b0000000000000000;
	sram_mem[72602] = 16'b0000000000000000;
	sram_mem[72603] = 16'b0000000000000000;
	sram_mem[72604] = 16'b0000000000000000;
	sram_mem[72605] = 16'b0000000000000000;
	sram_mem[72606] = 16'b0000000000000000;
	sram_mem[72607] = 16'b0000000000000000;
	sram_mem[72608] = 16'b0000000000000000;
	sram_mem[72609] = 16'b0000000000000000;
	sram_mem[72610] = 16'b0000000000000000;
	sram_mem[72611] = 16'b0000000000000000;
	sram_mem[72612] = 16'b0000000000000000;
	sram_mem[72613] = 16'b0000000000000000;
	sram_mem[72614] = 16'b0000000000000000;
	sram_mem[72615] = 16'b0000000000000000;
	sram_mem[72616] = 16'b0000000000000000;
	sram_mem[72617] = 16'b0000000000000000;
	sram_mem[72618] = 16'b0000000000000000;
	sram_mem[72619] = 16'b0000000000000000;
	sram_mem[72620] = 16'b0000000000000000;
	sram_mem[72621] = 16'b0000000000000000;
	sram_mem[72622] = 16'b0000000000000000;
	sram_mem[72623] = 16'b0000000000000000;
	sram_mem[72624] = 16'b0000000000000000;
	sram_mem[72625] = 16'b0000000000000000;
	sram_mem[72626] = 16'b0000000000000000;
	sram_mem[72627] = 16'b0000000000000000;
	sram_mem[72628] = 16'b0000000000000000;
	sram_mem[72629] = 16'b0000000000000000;
	sram_mem[72630] = 16'b0000000000000000;
	sram_mem[72631] = 16'b0000000000000000;
	sram_mem[72632] = 16'b0000000000000000;
	sram_mem[72633] = 16'b0000000000000000;
	sram_mem[72634] = 16'b0000000000000000;
	sram_mem[72635] = 16'b0000000000000000;
	sram_mem[72636] = 16'b0000000000000000;
	sram_mem[72637] = 16'b0000000000000000;
	sram_mem[72638] = 16'b0000000000000000;
	sram_mem[72639] = 16'b0000000000000000;
	sram_mem[72640] = 16'b0000000000000000;
	sram_mem[72641] = 16'b0000000000000000;
	sram_mem[72642] = 16'b0000000000000000;
	sram_mem[72643] = 16'b0000000000000000;
	sram_mem[72644] = 16'b0000000000000000;
	sram_mem[72645] = 16'b0000000000000000;
	sram_mem[72646] = 16'b0000000000000000;
	sram_mem[72647] = 16'b0000000000000000;
	sram_mem[72648] = 16'b0000000000000000;
	sram_mem[72649] = 16'b0000000000000000;
	sram_mem[72650] = 16'b0000000000000000;
	sram_mem[72651] = 16'b0000000000000000;
	sram_mem[72652] = 16'b0000000000000000;
	sram_mem[72653] = 16'b0000000000000000;
	sram_mem[72654] = 16'b0000000000000000;
	sram_mem[72655] = 16'b0000000000000000;
	sram_mem[72656] = 16'b0000000000000000;
	sram_mem[72657] = 16'b0000000000000000;
	sram_mem[72658] = 16'b0000000000000000;
	sram_mem[72659] = 16'b0000000000000000;
	sram_mem[72660] = 16'b0000000000000000;
	sram_mem[72661] = 16'b0000000000000000;
	sram_mem[72662] = 16'b0000000000000000;
	sram_mem[72663] = 16'b0000000000000000;
	sram_mem[72664] = 16'b0000000000000000;
	sram_mem[72665] = 16'b0000000000000000;
	sram_mem[72666] = 16'b0000000000000000;
	sram_mem[72667] = 16'b0000000000000000;
	sram_mem[72668] = 16'b0000000000000000;
	sram_mem[72669] = 16'b0000000000000000;
	sram_mem[72670] = 16'b0000000000000000;
	sram_mem[72671] = 16'b0000000000000000;
	sram_mem[72672] = 16'b0000000000000000;
	sram_mem[72673] = 16'b0000000000000000;
	sram_mem[72674] = 16'b0000000000000000;
	sram_mem[72675] = 16'b0000000000000000;
	sram_mem[72676] = 16'b0000000000000000;
	sram_mem[72677] = 16'b0000000000000000;
	sram_mem[72678] = 16'b0000000000000000;
	sram_mem[72679] = 16'b0000000000000000;
	sram_mem[72680] = 16'b0000000000000000;
	sram_mem[72681] = 16'b0000000000000000;
	sram_mem[72682] = 16'b0000000000000000;
	sram_mem[72683] = 16'b0000000000000000;
	sram_mem[72684] = 16'b0000000000000000;
	sram_mem[72685] = 16'b0000000000000000;
	sram_mem[72686] = 16'b0000000000000000;
	sram_mem[72687] = 16'b0000000000000000;
	sram_mem[72688] = 16'b0000000000000000;
	sram_mem[72689] = 16'b0000000000000000;
	sram_mem[72690] = 16'b0000000000000000;
	sram_mem[72691] = 16'b0000000000000000;
	sram_mem[72692] = 16'b0000000000000000;
	sram_mem[72693] = 16'b0000000000000000;
	sram_mem[72694] = 16'b0000000000000000;
	sram_mem[72695] = 16'b0000000000000000;
	sram_mem[72696] = 16'b0000000000000000;
	sram_mem[72697] = 16'b0000000000000000;
	sram_mem[72698] = 16'b0000000000000000;
	sram_mem[72699] = 16'b0000000000000000;
	sram_mem[72700] = 16'b0000000000000000;
	sram_mem[72701] = 16'b0000000000000000;
	sram_mem[72702] = 16'b0000000000000000;
	sram_mem[72703] = 16'b0000000000000000;
	sram_mem[72704] = 16'b0000000000000000;
	sram_mem[72705] = 16'b0000000000000000;
	sram_mem[72706] = 16'b0000000000000000;
	sram_mem[72707] = 16'b0000000000000000;
	sram_mem[72708] = 16'b0000000000000000;
	sram_mem[72709] = 16'b0000000000000000;
	sram_mem[72710] = 16'b0000000000000000;
	sram_mem[72711] = 16'b0000000000000000;
	sram_mem[72712] = 16'b0000000000000000;
	sram_mem[72713] = 16'b0000000000000000;
	sram_mem[72714] = 16'b0000000000000000;
	sram_mem[72715] = 16'b0000000000000000;
	sram_mem[72716] = 16'b0000000000000000;
	sram_mem[72717] = 16'b0000000000000000;
	sram_mem[72718] = 16'b0000000000000000;
	sram_mem[72719] = 16'b0000000000000000;
	sram_mem[72720] = 16'b0000000000000000;
	sram_mem[72721] = 16'b0000000000000000;
	sram_mem[72722] = 16'b0000000000000000;
	sram_mem[72723] = 16'b0000000000000000;
	sram_mem[72724] = 16'b0000000000000000;
	sram_mem[72725] = 16'b0000000000000000;
	sram_mem[72726] = 16'b0000000000000000;
	sram_mem[72727] = 16'b0000000000000000;
	sram_mem[72728] = 16'b0000000000000000;
	sram_mem[72729] = 16'b0000000000000000;
	sram_mem[72730] = 16'b0000000000000000;
	sram_mem[72731] = 16'b0000000000000000;
	sram_mem[72732] = 16'b0000000000000000;
	sram_mem[72733] = 16'b0000000000000000;
	sram_mem[72734] = 16'b0000000000000000;
	sram_mem[72735] = 16'b0000000000000000;
	sram_mem[72736] = 16'b0000000000000000;
	sram_mem[72737] = 16'b0000000000000000;
	sram_mem[72738] = 16'b0000000000000000;
	sram_mem[72739] = 16'b0000000000000000;
	sram_mem[72740] = 16'b0000000000000000;
	sram_mem[72741] = 16'b0000000000000000;
	sram_mem[72742] = 16'b0000000000000000;
	sram_mem[72743] = 16'b0000000000000000;
	sram_mem[72744] = 16'b0000000000000000;
	sram_mem[72745] = 16'b0000000000000000;
	sram_mem[72746] = 16'b0000000000000000;
	sram_mem[72747] = 16'b0000000000000000;
	sram_mem[72748] = 16'b0000000000000000;
	sram_mem[72749] = 16'b0000000000000000;
	sram_mem[72750] = 16'b0000000000000000;
	sram_mem[72751] = 16'b0000000000000000;
	sram_mem[72752] = 16'b0000000000000000;
	sram_mem[72753] = 16'b0000000000000000;
	sram_mem[72754] = 16'b0000000000000000;
	sram_mem[72755] = 16'b0000000000000000;
	sram_mem[72756] = 16'b0000000000000000;
	sram_mem[72757] = 16'b0000000000000000;
	sram_mem[72758] = 16'b0000000000000000;
	sram_mem[72759] = 16'b0000000000000000;
	sram_mem[72760] = 16'b0000000000000000;
	sram_mem[72761] = 16'b0000000000000000;
	sram_mem[72762] = 16'b0000000000000000;
	sram_mem[72763] = 16'b0000000000000000;
	sram_mem[72764] = 16'b0000000000000000;
	sram_mem[72765] = 16'b0000000000000000;
	sram_mem[72766] = 16'b0000000000000000;
	sram_mem[72767] = 16'b0000000000000000;
	sram_mem[72768] = 16'b0000000000000000;
	sram_mem[72769] = 16'b0000000000000000;
	sram_mem[72770] = 16'b0000000000000000;
	sram_mem[72771] = 16'b0000000000000000;
	sram_mem[72772] = 16'b0000000000000000;
	sram_mem[72773] = 16'b0000000000000000;
	sram_mem[72774] = 16'b0000000000000000;
	sram_mem[72775] = 16'b0000000000000000;
	sram_mem[72776] = 16'b0000000000000000;
	sram_mem[72777] = 16'b0000000000000000;
	sram_mem[72778] = 16'b0000000000000000;
	sram_mem[72779] = 16'b0000000000000000;
	sram_mem[72780] = 16'b0000000000000000;
	sram_mem[72781] = 16'b0000000000000000;
	sram_mem[72782] = 16'b0000000000000000;
	sram_mem[72783] = 16'b0000000000000000;
	sram_mem[72784] = 16'b0000000000000000;
	sram_mem[72785] = 16'b0000000000000000;
	sram_mem[72786] = 16'b0000000000000000;
	sram_mem[72787] = 16'b0000000000000000;
	sram_mem[72788] = 16'b0000000000000000;
	sram_mem[72789] = 16'b0000000000000000;
	sram_mem[72790] = 16'b0000000000000000;
	sram_mem[72791] = 16'b0000000000000000;
	sram_mem[72792] = 16'b0000000000000000;
	sram_mem[72793] = 16'b0000000000000000;
	sram_mem[72794] = 16'b0000000000000000;
	sram_mem[72795] = 16'b0000000000000000;
	sram_mem[72796] = 16'b0000000000000000;
	sram_mem[72797] = 16'b0000000000000000;
	sram_mem[72798] = 16'b0000000000000000;
	sram_mem[72799] = 16'b0000000000000000;
	sram_mem[72800] = 16'b0000000000000000;
	sram_mem[72801] = 16'b0000000000000000;
	sram_mem[72802] = 16'b0000000000000000;
	sram_mem[72803] = 16'b0000000000000000;
	sram_mem[72804] = 16'b0000000000000000;
	sram_mem[72805] = 16'b0000000000000000;
	sram_mem[72806] = 16'b0000000000000000;
	sram_mem[72807] = 16'b0000000000000000;
	sram_mem[72808] = 16'b0000000000000000;
	sram_mem[72809] = 16'b0000000000000000;
	sram_mem[72810] = 16'b0000000000000000;
	sram_mem[72811] = 16'b0000000000000000;
	sram_mem[72812] = 16'b0000000000000000;
	sram_mem[72813] = 16'b0000000000000000;
	sram_mem[72814] = 16'b0000000000000000;
	sram_mem[72815] = 16'b0000000000000000;
	sram_mem[72816] = 16'b0000000000000000;
	sram_mem[72817] = 16'b0000000000000000;
	sram_mem[72818] = 16'b0000000000000000;
	sram_mem[72819] = 16'b0000000000000000;
	sram_mem[72820] = 16'b0000000000000000;
	sram_mem[72821] = 16'b0000000000000000;
	sram_mem[72822] = 16'b0000000000000000;
	sram_mem[72823] = 16'b0000000000000000;
	sram_mem[72824] = 16'b0000000000000000;
	sram_mem[72825] = 16'b0000000000000000;
	sram_mem[72826] = 16'b0000000000000000;
	sram_mem[72827] = 16'b0000000000000000;
	sram_mem[72828] = 16'b0000000000000000;
	sram_mem[72829] = 16'b0000000000000000;
	sram_mem[72830] = 16'b0000000000000000;
	sram_mem[72831] = 16'b0000000000000000;
	sram_mem[72832] = 16'b0000000000000000;
	sram_mem[72833] = 16'b0000000000000000;
	sram_mem[72834] = 16'b0000000000000000;
	sram_mem[72835] = 16'b0000000000000000;
	sram_mem[72836] = 16'b0000000000000000;
	sram_mem[72837] = 16'b0000000000000000;
	sram_mem[72838] = 16'b0000000000000000;
	sram_mem[72839] = 16'b0000000000000000;
	sram_mem[72840] = 16'b0000000000000000;
	sram_mem[72841] = 16'b0000000000000000;
	sram_mem[72842] = 16'b0000000000000000;
	sram_mem[72843] = 16'b0000000000000000;
	sram_mem[72844] = 16'b0000000000000000;
	sram_mem[72845] = 16'b0000000000000000;
	sram_mem[72846] = 16'b0000000000000000;
	sram_mem[72847] = 16'b0000000000000000;
	sram_mem[72848] = 16'b0000000000000000;
	sram_mem[72849] = 16'b0000000000000000;
	sram_mem[72850] = 16'b0000000000000000;
	sram_mem[72851] = 16'b0000000000000000;
	sram_mem[72852] = 16'b0000000000000000;
	sram_mem[72853] = 16'b0000000000000000;
	sram_mem[72854] = 16'b0000000000000000;
	sram_mem[72855] = 16'b0000000000000000;
	sram_mem[72856] = 16'b0000000000000000;
	sram_mem[72857] = 16'b0000000000000000;
	sram_mem[72858] = 16'b0000000000000000;
	sram_mem[72859] = 16'b0000000000000000;
	sram_mem[72860] = 16'b0000000000000000;
	sram_mem[72861] = 16'b0000000000000000;
	sram_mem[72862] = 16'b0000000000000000;
	sram_mem[72863] = 16'b0000000000000000;
	sram_mem[72864] = 16'b0000000000000000;
	sram_mem[72865] = 16'b0000000000000000;
	sram_mem[72866] = 16'b0000000000000000;
	sram_mem[72867] = 16'b0000000000000000;
	sram_mem[72868] = 16'b0000000000000000;
	sram_mem[72869] = 16'b0000000000000000;
	sram_mem[72870] = 16'b0000000000000000;
	sram_mem[72871] = 16'b0000000000000000;
	sram_mem[72872] = 16'b0000000000000000;
	sram_mem[72873] = 16'b0000000000000000;
	sram_mem[72874] = 16'b0000000000000000;
	sram_mem[72875] = 16'b0000000000000000;
	sram_mem[72876] = 16'b0000000000000000;
	sram_mem[72877] = 16'b0000000000000000;
	sram_mem[72878] = 16'b0000000000000000;
	sram_mem[72879] = 16'b0000000000000000;
	sram_mem[72880] = 16'b0000000000000000;
	sram_mem[72881] = 16'b0000000000000000;
	sram_mem[72882] = 16'b0000000000000000;
	sram_mem[72883] = 16'b0000000000000000;
	sram_mem[72884] = 16'b0000000000000000;
	sram_mem[72885] = 16'b0000000000000000;
	sram_mem[72886] = 16'b0000000000000000;
	sram_mem[72887] = 16'b0000000000000000;
	sram_mem[72888] = 16'b0000000000000000;
	sram_mem[72889] = 16'b0000000000000000;
	sram_mem[72890] = 16'b0000000000000000;
	sram_mem[72891] = 16'b0000000000000000;
	sram_mem[72892] = 16'b0000000000000000;
	sram_mem[72893] = 16'b0000000000000000;
	sram_mem[72894] = 16'b0000000000000000;
	sram_mem[72895] = 16'b0000000000000000;
	sram_mem[72896] = 16'b0000000000000000;
	sram_mem[72897] = 16'b0000000000000000;
	sram_mem[72898] = 16'b0000000000000000;
	sram_mem[72899] = 16'b0000000000000000;
	sram_mem[72900] = 16'b0000000000000000;
	sram_mem[72901] = 16'b0000000000000000;
	sram_mem[72902] = 16'b0000000000000000;
	sram_mem[72903] = 16'b0000000000000000;
	sram_mem[72904] = 16'b0000000000000000;
	sram_mem[72905] = 16'b0000000000000000;
	sram_mem[72906] = 16'b0000000000000000;
	sram_mem[72907] = 16'b0000000000000000;
	sram_mem[72908] = 16'b0000000000000000;
	sram_mem[72909] = 16'b0000000000000000;
	sram_mem[72910] = 16'b0000000000000000;
	sram_mem[72911] = 16'b0000000000000000;
	sram_mem[72912] = 16'b0000000000000000;
	sram_mem[72913] = 16'b0000000000000000;
	sram_mem[72914] = 16'b0000000000000000;
	sram_mem[72915] = 16'b0000000000000000;
	sram_mem[72916] = 16'b0000000000000000;
	sram_mem[72917] = 16'b0000000000000000;
	sram_mem[72918] = 16'b0000000000000000;
	sram_mem[72919] = 16'b0000000000000000;
	sram_mem[72920] = 16'b0000000000000000;
	sram_mem[72921] = 16'b0000000000000000;
	sram_mem[72922] = 16'b0000000000000000;
	sram_mem[72923] = 16'b0000000000000000;
	sram_mem[72924] = 16'b0000000000000000;
	sram_mem[72925] = 16'b0000000000000000;
	sram_mem[72926] = 16'b0000000000000000;
	sram_mem[72927] = 16'b0000000000000000;
	sram_mem[72928] = 16'b0000000000000000;
	sram_mem[72929] = 16'b0000000000000000;
	sram_mem[72930] = 16'b0000000000000000;
	sram_mem[72931] = 16'b0000000000000000;
	sram_mem[72932] = 16'b0000000000000000;
	sram_mem[72933] = 16'b0000000000000000;
	sram_mem[72934] = 16'b0000000000000000;
	sram_mem[72935] = 16'b0000000000000000;
	sram_mem[72936] = 16'b0000000000000000;
	sram_mem[72937] = 16'b0000000000000000;
	sram_mem[72938] = 16'b0000000000000000;
	sram_mem[72939] = 16'b0000000000000000;
	sram_mem[72940] = 16'b0000000000000000;
	sram_mem[72941] = 16'b0000000000000000;
	sram_mem[72942] = 16'b0000000000000000;
	sram_mem[72943] = 16'b0000000000000000;
	sram_mem[72944] = 16'b0000000000000000;
	sram_mem[72945] = 16'b0000000000000000;
	sram_mem[72946] = 16'b0000000000000000;
	sram_mem[72947] = 16'b0000000000000000;
	sram_mem[72948] = 16'b0000000000000000;
	sram_mem[72949] = 16'b0000000000000000;
	sram_mem[72950] = 16'b0000000000000000;
	sram_mem[72951] = 16'b0000000000000000;
	sram_mem[72952] = 16'b0000000000000000;
	sram_mem[72953] = 16'b0000000000000000;
	sram_mem[72954] = 16'b0000000000000000;
	sram_mem[72955] = 16'b0000000000000000;
	sram_mem[72956] = 16'b0000000000000000;
	sram_mem[72957] = 16'b0000000000000000;
	sram_mem[72958] = 16'b0000000000000000;
	sram_mem[72959] = 16'b0000000000000000;
	sram_mem[72960] = 16'b0000000000000000;
	sram_mem[72961] = 16'b0000000000000000;
	sram_mem[72962] = 16'b0000000000000000;
	sram_mem[72963] = 16'b0000000000000000;
	sram_mem[72964] = 16'b0000000000000000;
	sram_mem[72965] = 16'b0000000000000000;
	sram_mem[72966] = 16'b0000000000000000;
	sram_mem[72967] = 16'b0000000000000000;
	sram_mem[72968] = 16'b0000000000000000;
	sram_mem[72969] = 16'b0000000000000000;
	sram_mem[72970] = 16'b0000000000000000;
	sram_mem[72971] = 16'b0000000000000000;
	sram_mem[72972] = 16'b0000000000000000;
	sram_mem[72973] = 16'b0000000000000000;
	sram_mem[72974] = 16'b0000000000000000;
	sram_mem[72975] = 16'b0000000000000000;
	sram_mem[72976] = 16'b0000000000000000;
	sram_mem[72977] = 16'b0000000000000000;
	sram_mem[72978] = 16'b0000000000000000;
	sram_mem[72979] = 16'b0000000000000000;
	sram_mem[72980] = 16'b0000000000000000;
	sram_mem[72981] = 16'b0000000000000000;
	sram_mem[72982] = 16'b0000000000000000;
	sram_mem[72983] = 16'b0000000000000000;
	sram_mem[72984] = 16'b0000000000000000;
	sram_mem[72985] = 16'b0000000000000000;
	sram_mem[72986] = 16'b0000000000000000;
	sram_mem[72987] = 16'b0000000000000000;
	sram_mem[72988] = 16'b0000000000000000;
	sram_mem[72989] = 16'b0000000000000000;
	sram_mem[72990] = 16'b0000000000000000;
	sram_mem[72991] = 16'b0000000000000000;
	sram_mem[72992] = 16'b0000000000000000;
	sram_mem[72993] = 16'b0000000000000000;
	sram_mem[72994] = 16'b0000000000000000;
	sram_mem[72995] = 16'b0000000000000000;
	sram_mem[72996] = 16'b0000000000000000;
	sram_mem[72997] = 16'b0000000000000000;
	sram_mem[72998] = 16'b0000000000000000;
	sram_mem[72999] = 16'b0000000000000000;
	sram_mem[73000] = 16'b0000000000000000;
	sram_mem[73001] = 16'b0000000000000000;
	sram_mem[73002] = 16'b0000000000000000;
	sram_mem[73003] = 16'b0000000000000000;
	sram_mem[73004] = 16'b0000000000000000;
	sram_mem[73005] = 16'b0000000000000000;
	sram_mem[73006] = 16'b0000000000000000;
	sram_mem[73007] = 16'b0000000000000000;
	sram_mem[73008] = 16'b0000000000000000;
	sram_mem[73009] = 16'b0000000000000000;
	sram_mem[73010] = 16'b0000000000000000;
	sram_mem[73011] = 16'b0000000000000000;
	sram_mem[73012] = 16'b0000000000000000;
	sram_mem[73013] = 16'b0000000000000000;
	sram_mem[73014] = 16'b0000000000000000;
	sram_mem[73015] = 16'b0000000000000000;
	sram_mem[73016] = 16'b0000000000000000;
	sram_mem[73017] = 16'b0000000000000000;
	sram_mem[73018] = 16'b0000000000000000;
	sram_mem[73019] = 16'b0000000000000000;
	sram_mem[73020] = 16'b0000000000000000;
	sram_mem[73021] = 16'b0000000000000000;
	sram_mem[73022] = 16'b0000000000000000;
	sram_mem[73023] = 16'b0000000000000000;
	sram_mem[73024] = 16'b0000000000000000;
	sram_mem[73025] = 16'b0000000000000000;
	sram_mem[73026] = 16'b0000000000000000;
	sram_mem[73027] = 16'b0000000000000000;
	sram_mem[73028] = 16'b0000000000000000;
	sram_mem[73029] = 16'b0000000000000000;
	sram_mem[73030] = 16'b0000000000000000;
	sram_mem[73031] = 16'b0000000000000000;
	sram_mem[73032] = 16'b0000000000000000;
	sram_mem[73033] = 16'b0000000000000000;
	sram_mem[73034] = 16'b0000000000000000;
	sram_mem[73035] = 16'b0000000000000000;
	sram_mem[73036] = 16'b0000000000000000;
	sram_mem[73037] = 16'b0000000000000000;
	sram_mem[73038] = 16'b0000000000000000;
	sram_mem[73039] = 16'b0000000000000000;
	sram_mem[73040] = 16'b0000000000000000;
	sram_mem[73041] = 16'b0000000000000000;
	sram_mem[73042] = 16'b0000000000000000;
	sram_mem[73043] = 16'b0000000000000000;
	sram_mem[73044] = 16'b0000000000000000;
	sram_mem[73045] = 16'b0000000000000000;
	sram_mem[73046] = 16'b0000000000000000;
	sram_mem[73047] = 16'b0000000000000000;
	sram_mem[73048] = 16'b0000000000000000;
	sram_mem[73049] = 16'b0000000000000000;
	sram_mem[73050] = 16'b0000000000000000;
	sram_mem[73051] = 16'b0000000000000000;
	sram_mem[73052] = 16'b0000000000000000;
	sram_mem[73053] = 16'b0000000000000000;
	sram_mem[73054] = 16'b0000000000000000;
	sram_mem[73055] = 16'b0000000000000000;
	sram_mem[73056] = 16'b0000000000000000;
	sram_mem[73057] = 16'b0000000000000000;
	sram_mem[73058] = 16'b0000000000000000;
	sram_mem[73059] = 16'b0000000000000000;
	sram_mem[73060] = 16'b0000000000000000;
	sram_mem[73061] = 16'b0000000000000000;
	sram_mem[73062] = 16'b0000000000000000;
	sram_mem[73063] = 16'b0000000000000000;
	sram_mem[73064] = 16'b0000000000000000;
	sram_mem[73065] = 16'b0000000000000000;
	sram_mem[73066] = 16'b0000000000000000;
	sram_mem[73067] = 16'b0000000000000000;
	sram_mem[73068] = 16'b0000000000000000;
	sram_mem[73069] = 16'b0000000000000000;
	sram_mem[73070] = 16'b0000000000000000;
	sram_mem[73071] = 16'b0000000000000000;
	sram_mem[73072] = 16'b0000000000000000;
	sram_mem[73073] = 16'b0000000000000000;
	sram_mem[73074] = 16'b0000000000000000;
	sram_mem[73075] = 16'b0000000000000000;
	sram_mem[73076] = 16'b0000000000000000;
	sram_mem[73077] = 16'b0000000000000000;
	sram_mem[73078] = 16'b0000000000000000;
	sram_mem[73079] = 16'b0000000000000000;
	sram_mem[73080] = 16'b0000000000000000;
	sram_mem[73081] = 16'b0000000000000000;
	sram_mem[73082] = 16'b0000000000000000;
	sram_mem[73083] = 16'b0000000000000000;
	sram_mem[73084] = 16'b0000000000000000;
	sram_mem[73085] = 16'b0000000000000000;
	sram_mem[73086] = 16'b0000000000000000;
	sram_mem[73087] = 16'b0000000000000000;
	sram_mem[73088] = 16'b0000000000000000;
	sram_mem[73089] = 16'b0000000000000000;
	sram_mem[73090] = 16'b0000000000000000;
	sram_mem[73091] = 16'b0000000000000000;
	sram_mem[73092] = 16'b0000000000000000;
	sram_mem[73093] = 16'b0000000000000000;
	sram_mem[73094] = 16'b0000000000000000;
	sram_mem[73095] = 16'b0000000000000000;
	sram_mem[73096] = 16'b0000000000000000;
	sram_mem[73097] = 16'b0000000000000000;
	sram_mem[73098] = 16'b0000000000000000;
	sram_mem[73099] = 16'b0000000000000000;
	sram_mem[73100] = 16'b0000000000000000;
	sram_mem[73101] = 16'b0000000000000000;
	sram_mem[73102] = 16'b0000000000000000;
	sram_mem[73103] = 16'b0000000000000000;
	sram_mem[73104] = 16'b0000000000000000;
	sram_mem[73105] = 16'b0000000000000000;
	sram_mem[73106] = 16'b0000000000000000;
	sram_mem[73107] = 16'b0000000000000000;
	sram_mem[73108] = 16'b0000000000000000;
	sram_mem[73109] = 16'b0000000000000000;
	sram_mem[73110] = 16'b0000000000000000;
	sram_mem[73111] = 16'b0000000000000000;
	sram_mem[73112] = 16'b0000000000000000;
	sram_mem[73113] = 16'b0000000000000000;
	sram_mem[73114] = 16'b0000000000000000;
	sram_mem[73115] = 16'b0000000000000000;
	sram_mem[73116] = 16'b0000000000000000;
	sram_mem[73117] = 16'b0000000000000000;
	sram_mem[73118] = 16'b0000000000000000;
	sram_mem[73119] = 16'b0000000000000000;
	sram_mem[73120] = 16'b0000000000000000;
	sram_mem[73121] = 16'b0000000000000000;
	sram_mem[73122] = 16'b0000000000000000;
	sram_mem[73123] = 16'b0000000000000000;
	sram_mem[73124] = 16'b0000000000000000;
	sram_mem[73125] = 16'b0000000000000000;
	sram_mem[73126] = 16'b0000000000000000;
	sram_mem[73127] = 16'b0000000000000000;
	sram_mem[73128] = 16'b0000000000000000;
	sram_mem[73129] = 16'b0000000000000000;
	sram_mem[73130] = 16'b0000000000000000;
	sram_mem[73131] = 16'b0000000000000000;
	sram_mem[73132] = 16'b0000000000000000;
	sram_mem[73133] = 16'b0000000000000000;
	sram_mem[73134] = 16'b0000000000000000;
	sram_mem[73135] = 16'b0000000000000000;
	sram_mem[73136] = 16'b0000000000000000;
	sram_mem[73137] = 16'b0000000000000000;
	sram_mem[73138] = 16'b0000000000000000;
	sram_mem[73139] = 16'b0000000000000000;
	sram_mem[73140] = 16'b0000000000000000;
	sram_mem[73141] = 16'b0000000000000000;
	sram_mem[73142] = 16'b0000000000000000;
	sram_mem[73143] = 16'b0000000000000000;
	sram_mem[73144] = 16'b0000000000000000;
	sram_mem[73145] = 16'b0000000000000000;
	sram_mem[73146] = 16'b0000000000000000;
	sram_mem[73147] = 16'b0000000000000000;
	sram_mem[73148] = 16'b0000000000000000;
	sram_mem[73149] = 16'b0000000000000000;
	sram_mem[73150] = 16'b0000000000000000;
	sram_mem[73151] = 16'b0000000000000000;
	sram_mem[73152] = 16'b0000000000000000;
	sram_mem[73153] = 16'b0000000000000000;
	sram_mem[73154] = 16'b0000000000000000;
	sram_mem[73155] = 16'b0000000000000000;
	sram_mem[73156] = 16'b0000000000000000;
	sram_mem[73157] = 16'b0000000000000000;
	sram_mem[73158] = 16'b0000000000000000;
	sram_mem[73159] = 16'b0000000000000000;
	sram_mem[73160] = 16'b0000000000000000;
	sram_mem[73161] = 16'b0000000000000000;
	sram_mem[73162] = 16'b0000000000000000;
	sram_mem[73163] = 16'b0000000000000000;
	sram_mem[73164] = 16'b0000000000000000;
	sram_mem[73165] = 16'b0000000000000000;
	sram_mem[73166] = 16'b0000000000000000;
	sram_mem[73167] = 16'b0000000000000000;
	sram_mem[73168] = 16'b0000000000000000;
	sram_mem[73169] = 16'b0000000000000000;
	sram_mem[73170] = 16'b0000000000000000;
	sram_mem[73171] = 16'b0000000000000000;
	sram_mem[73172] = 16'b0000000000000000;
	sram_mem[73173] = 16'b0000000000000000;
	sram_mem[73174] = 16'b0000000000000000;
	sram_mem[73175] = 16'b0000000000000000;
	sram_mem[73176] = 16'b0000000000000000;
	sram_mem[73177] = 16'b0000000000000000;
	sram_mem[73178] = 16'b0000000000000000;
	sram_mem[73179] = 16'b0000000000000000;
	sram_mem[73180] = 16'b0000000000000000;
	sram_mem[73181] = 16'b0000000000000000;
	sram_mem[73182] = 16'b0000000000000000;
	sram_mem[73183] = 16'b0000000000000000;
	sram_mem[73184] = 16'b0000000000000000;
	sram_mem[73185] = 16'b0000000000000000;
	sram_mem[73186] = 16'b0000000000000000;
	sram_mem[73187] = 16'b0000000000000000;
	sram_mem[73188] = 16'b0000000000000000;
	sram_mem[73189] = 16'b0000000000000000;
	sram_mem[73190] = 16'b0000000000000000;
	sram_mem[73191] = 16'b0000000000000000;
	sram_mem[73192] = 16'b0000000000000000;
	sram_mem[73193] = 16'b0000000000000000;
	sram_mem[73194] = 16'b0000000000000000;
	sram_mem[73195] = 16'b0000000000000000;
	sram_mem[73196] = 16'b0000000000000000;
	sram_mem[73197] = 16'b0000000000000000;
	sram_mem[73198] = 16'b0000000000000000;
	sram_mem[73199] = 16'b0000000000000000;
	sram_mem[73200] = 16'b0000000000000000;
	sram_mem[73201] = 16'b0000000000000000;
	sram_mem[73202] = 16'b0000000000000000;
	sram_mem[73203] = 16'b0000000000000000;
	sram_mem[73204] = 16'b0000000000000000;
	sram_mem[73205] = 16'b0000000000000000;
	sram_mem[73206] = 16'b0000000000000000;
	sram_mem[73207] = 16'b0000000000000000;
	sram_mem[73208] = 16'b0000000000000000;
	sram_mem[73209] = 16'b0000000000000000;
	sram_mem[73210] = 16'b0000000000000000;
	sram_mem[73211] = 16'b0000000000000000;
	sram_mem[73212] = 16'b0000000000000000;
	sram_mem[73213] = 16'b0000000000000000;
	sram_mem[73214] = 16'b0000000000000000;
	sram_mem[73215] = 16'b0000000000000000;
	sram_mem[73216] = 16'b0000000000000000;
	sram_mem[73217] = 16'b0000000000000000;
	sram_mem[73218] = 16'b0000000000000000;
	sram_mem[73219] = 16'b0000000000000000;
	sram_mem[73220] = 16'b0000000000000000;
	sram_mem[73221] = 16'b0000000000000000;
	sram_mem[73222] = 16'b0000000000000000;
	sram_mem[73223] = 16'b0000000000000000;
	sram_mem[73224] = 16'b0000000000000000;
	sram_mem[73225] = 16'b0000000000000000;
	sram_mem[73226] = 16'b0000000000000000;
	sram_mem[73227] = 16'b0000000000000000;
	sram_mem[73228] = 16'b0000000000000000;
	sram_mem[73229] = 16'b0000000000000000;
	sram_mem[73230] = 16'b0000000000000000;
	sram_mem[73231] = 16'b0000000000000000;
	sram_mem[73232] = 16'b0000000000000000;
	sram_mem[73233] = 16'b0000000000000000;
	sram_mem[73234] = 16'b0000000000000000;
	sram_mem[73235] = 16'b0000000000000000;
	sram_mem[73236] = 16'b0000000000000000;
	sram_mem[73237] = 16'b0000000000000000;
	sram_mem[73238] = 16'b0000000000000000;
	sram_mem[73239] = 16'b0000000000000000;
	sram_mem[73240] = 16'b0000000000000000;
	sram_mem[73241] = 16'b0000000000000000;
	sram_mem[73242] = 16'b0000000000000000;
	sram_mem[73243] = 16'b0000000000000000;
	sram_mem[73244] = 16'b0000000000000000;
	sram_mem[73245] = 16'b0000000000000000;
	sram_mem[73246] = 16'b0000000000000000;
	sram_mem[73247] = 16'b0000000000000000;
	sram_mem[73248] = 16'b0000000000000000;
	sram_mem[73249] = 16'b0000000000000000;
	sram_mem[73250] = 16'b0000000000000000;
	sram_mem[73251] = 16'b0000000000000000;
	sram_mem[73252] = 16'b0000000000000000;
	sram_mem[73253] = 16'b0000000000000000;
	sram_mem[73254] = 16'b0000000000000000;
	sram_mem[73255] = 16'b0000000000000000;
	sram_mem[73256] = 16'b0000000000000000;
	sram_mem[73257] = 16'b0000000000000000;
	sram_mem[73258] = 16'b0000000000000000;
	sram_mem[73259] = 16'b0000000000000000;
	sram_mem[73260] = 16'b0000000000000000;
	sram_mem[73261] = 16'b0000000000000000;
	sram_mem[73262] = 16'b0000000000000000;
	sram_mem[73263] = 16'b0000000000000000;
	sram_mem[73264] = 16'b0000000000000000;
	sram_mem[73265] = 16'b0000000000000000;
	sram_mem[73266] = 16'b0000000000000000;
	sram_mem[73267] = 16'b0000000000000000;
	sram_mem[73268] = 16'b0000000000000000;
	sram_mem[73269] = 16'b0000000000000000;
	sram_mem[73270] = 16'b0000000000000000;
	sram_mem[73271] = 16'b0000000000000000;
	sram_mem[73272] = 16'b0000000000000000;
	sram_mem[73273] = 16'b0000000000000000;
	sram_mem[73274] = 16'b0000000000000000;
	sram_mem[73275] = 16'b0000000000000000;
	sram_mem[73276] = 16'b0000000000000000;
	sram_mem[73277] = 16'b0000000000000000;
	sram_mem[73278] = 16'b0000000000000000;
	sram_mem[73279] = 16'b0000000000000000;
	sram_mem[73280] = 16'b0000000000000000;
	sram_mem[73281] = 16'b0000000000000000;
	sram_mem[73282] = 16'b0000000000000000;
	sram_mem[73283] = 16'b0000000000000000;
	sram_mem[73284] = 16'b0000000000000000;
	sram_mem[73285] = 16'b0000000000000000;
	sram_mem[73286] = 16'b0000000000000000;
	sram_mem[73287] = 16'b0000000000000000;
	sram_mem[73288] = 16'b0000000000000000;
	sram_mem[73289] = 16'b0000000000000000;
	sram_mem[73290] = 16'b0000000000000000;
	sram_mem[73291] = 16'b0000000000000000;
	sram_mem[73292] = 16'b0000000000000000;
	sram_mem[73293] = 16'b0000000000000000;
	sram_mem[73294] = 16'b0000000000000000;
	sram_mem[73295] = 16'b0000000000000000;
	sram_mem[73296] = 16'b0000000000000000;
	sram_mem[73297] = 16'b0000000000000000;
	sram_mem[73298] = 16'b0000000000000000;
	sram_mem[73299] = 16'b0000000000000000;
	sram_mem[73300] = 16'b0000000000000000;
	sram_mem[73301] = 16'b0000000000000000;
	sram_mem[73302] = 16'b0000000000000000;
	sram_mem[73303] = 16'b0000000000000000;
	sram_mem[73304] = 16'b0000000000000000;
	sram_mem[73305] = 16'b0000000000000000;
	sram_mem[73306] = 16'b0000000000000000;
	sram_mem[73307] = 16'b0000000000000000;
	sram_mem[73308] = 16'b0000000000000000;
	sram_mem[73309] = 16'b0000000000000000;
	sram_mem[73310] = 16'b0000000000000000;
	sram_mem[73311] = 16'b0000000000000000;
	sram_mem[73312] = 16'b0000000000000000;
	sram_mem[73313] = 16'b0000000000000000;
	sram_mem[73314] = 16'b0000000000000000;
	sram_mem[73315] = 16'b0000000000000000;
	sram_mem[73316] = 16'b0000000000000000;
	sram_mem[73317] = 16'b0000000000000000;
	sram_mem[73318] = 16'b0000000000000000;
	sram_mem[73319] = 16'b0000000000000000;
	sram_mem[73320] = 16'b0000000000000000;
	sram_mem[73321] = 16'b0000000000000000;
	sram_mem[73322] = 16'b0000000000000000;
	sram_mem[73323] = 16'b0000000000000000;
	sram_mem[73324] = 16'b0000000000000000;
	sram_mem[73325] = 16'b0000000000000000;
	sram_mem[73326] = 16'b0000000000000000;
	sram_mem[73327] = 16'b0000000000000000;
	sram_mem[73328] = 16'b0000000000000000;
	sram_mem[73329] = 16'b0000000000000000;
	sram_mem[73330] = 16'b0000000000000000;
	sram_mem[73331] = 16'b0000000000000000;
	sram_mem[73332] = 16'b0000000000000000;
	sram_mem[73333] = 16'b0000000000000000;
	sram_mem[73334] = 16'b0000000000000000;
	sram_mem[73335] = 16'b0000000000000000;
	sram_mem[73336] = 16'b0000000000000000;
	sram_mem[73337] = 16'b0000000000000000;
	sram_mem[73338] = 16'b0000000000000000;
	sram_mem[73339] = 16'b0000000000000000;
	sram_mem[73340] = 16'b0000000000000000;
	sram_mem[73341] = 16'b0000000000000000;
	sram_mem[73342] = 16'b0000000000000000;
	sram_mem[73343] = 16'b0000000000000000;
	sram_mem[73344] = 16'b0000000000000000;
	sram_mem[73345] = 16'b0000000000000000;
	sram_mem[73346] = 16'b0000000000000000;
	sram_mem[73347] = 16'b0000000000000000;
	sram_mem[73348] = 16'b0000000000000000;
	sram_mem[73349] = 16'b0000000000000000;
	sram_mem[73350] = 16'b0000000000000000;
	sram_mem[73351] = 16'b0000000000000000;
	sram_mem[73352] = 16'b0000000000000000;
	sram_mem[73353] = 16'b0000000000000000;
	sram_mem[73354] = 16'b0000000000000000;
	sram_mem[73355] = 16'b0000000000000000;
	sram_mem[73356] = 16'b0000000000000000;
	sram_mem[73357] = 16'b0000000000000000;
	sram_mem[73358] = 16'b0000000000000000;
	sram_mem[73359] = 16'b0000000000000000;
	sram_mem[73360] = 16'b0000000000000000;
	sram_mem[73361] = 16'b0000000000000000;
	sram_mem[73362] = 16'b0000000000000000;
	sram_mem[73363] = 16'b0000000000000000;
	sram_mem[73364] = 16'b0000000000000000;
	sram_mem[73365] = 16'b0000000000000000;
	sram_mem[73366] = 16'b0000000000000000;
	sram_mem[73367] = 16'b0000000000000000;
	sram_mem[73368] = 16'b0000000000000000;
	sram_mem[73369] = 16'b0000000000000000;
	sram_mem[73370] = 16'b0000000000000000;
	sram_mem[73371] = 16'b0000000000000000;
	sram_mem[73372] = 16'b0000000000000000;
	sram_mem[73373] = 16'b0000000000000000;
	sram_mem[73374] = 16'b0000000000000000;
	sram_mem[73375] = 16'b0000000000000000;
	sram_mem[73376] = 16'b0000000000000000;
	sram_mem[73377] = 16'b0000000000000000;
	sram_mem[73378] = 16'b0000000000000000;
	sram_mem[73379] = 16'b0000000000000000;
	sram_mem[73380] = 16'b0000000000000000;
	sram_mem[73381] = 16'b0000000000000000;
	sram_mem[73382] = 16'b0000000000000000;
	sram_mem[73383] = 16'b0000000000000000;
	sram_mem[73384] = 16'b0000000000000000;
	sram_mem[73385] = 16'b0000000000000000;
	sram_mem[73386] = 16'b0000000000000000;
	sram_mem[73387] = 16'b0000000000000000;
	sram_mem[73388] = 16'b0000000000000000;
	sram_mem[73389] = 16'b0000000000000000;
	sram_mem[73390] = 16'b0000000000000000;
	sram_mem[73391] = 16'b0000000000000000;
	sram_mem[73392] = 16'b0000000000000000;
	sram_mem[73393] = 16'b0000000000000000;
	sram_mem[73394] = 16'b0000000000000000;
	sram_mem[73395] = 16'b0000000000000000;
	sram_mem[73396] = 16'b0000000000000000;
	sram_mem[73397] = 16'b0000000000000000;
	sram_mem[73398] = 16'b0000000000000000;
	sram_mem[73399] = 16'b0000000000000000;
	sram_mem[73400] = 16'b0000000000000000;
	sram_mem[73401] = 16'b0000000000000000;
	sram_mem[73402] = 16'b0000000000000000;
	sram_mem[73403] = 16'b0000000000000000;
	sram_mem[73404] = 16'b0000000000000000;
	sram_mem[73405] = 16'b0000000000000000;
	sram_mem[73406] = 16'b0000000000000000;
	sram_mem[73407] = 16'b0000000000000000;
	sram_mem[73408] = 16'b0000000000000000;
	sram_mem[73409] = 16'b0000000000000000;
	sram_mem[73410] = 16'b0000000000000000;
	sram_mem[73411] = 16'b0000000000000000;
	sram_mem[73412] = 16'b0000000000000000;
	sram_mem[73413] = 16'b0000000000000000;
	sram_mem[73414] = 16'b0000000000000000;
	sram_mem[73415] = 16'b0000000000000000;
	sram_mem[73416] = 16'b0000000000000000;
	sram_mem[73417] = 16'b0000000000000000;
	sram_mem[73418] = 16'b0000000000000000;
	sram_mem[73419] = 16'b0000000000000000;
	sram_mem[73420] = 16'b0000000000000000;
	sram_mem[73421] = 16'b0000000000000000;
	sram_mem[73422] = 16'b0000000000000000;
	sram_mem[73423] = 16'b0000000000000000;
	sram_mem[73424] = 16'b0000000000000000;
	sram_mem[73425] = 16'b0000000000000000;
	sram_mem[73426] = 16'b0000000000000000;
	sram_mem[73427] = 16'b0000000000000000;
	sram_mem[73428] = 16'b0000000000000000;
	sram_mem[73429] = 16'b0000000000000000;
	sram_mem[73430] = 16'b0000000000000000;
	sram_mem[73431] = 16'b0000000000000000;
	sram_mem[73432] = 16'b0000000000000000;
	sram_mem[73433] = 16'b0000000000000000;
	sram_mem[73434] = 16'b0000000000000000;
	sram_mem[73435] = 16'b0000000000000000;
	sram_mem[73436] = 16'b0000000000000000;
	sram_mem[73437] = 16'b0000000000000000;
	sram_mem[73438] = 16'b0000000000000000;
	sram_mem[73439] = 16'b0000000000000000;
	sram_mem[73440] = 16'b0000000000000000;
	sram_mem[73441] = 16'b0000000000000000;
	sram_mem[73442] = 16'b0000000000000000;
	sram_mem[73443] = 16'b0000000000000000;
	sram_mem[73444] = 16'b0000000000000000;
	sram_mem[73445] = 16'b0000000000000000;
	sram_mem[73446] = 16'b0000000000000000;
	sram_mem[73447] = 16'b0000000000000000;
	sram_mem[73448] = 16'b0000000000000000;
	sram_mem[73449] = 16'b0000000000000000;
	sram_mem[73450] = 16'b0000000000000000;
	sram_mem[73451] = 16'b0000000000000000;
	sram_mem[73452] = 16'b0000000000000000;
	sram_mem[73453] = 16'b0000000000000000;
	sram_mem[73454] = 16'b0000000000000000;
	sram_mem[73455] = 16'b0000000000000000;
	sram_mem[73456] = 16'b0000000000000000;
	sram_mem[73457] = 16'b0000000000000000;
	sram_mem[73458] = 16'b0000000000000000;
	sram_mem[73459] = 16'b0000000000000000;
	sram_mem[73460] = 16'b0000000000000000;
	sram_mem[73461] = 16'b0000000000000000;
	sram_mem[73462] = 16'b0000000000000000;
	sram_mem[73463] = 16'b0000000000000000;
	sram_mem[73464] = 16'b0000000000000000;
	sram_mem[73465] = 16'b0000000000000000;
	sram_mem[73466] = 16'b0000000000000000;
	sram_mem[73467] = 16'b0000000000000000;
	sram_mem[73468] = 16'b0000000000000000;
	sram_mem[73469] = 16'b0000000000000000;
	sram_mem[73470] = 16'b0000000000000000;
	sram_mem[73471] = 16'b0000000000000000;
	sram_mem[73472] = 16'b0000000000000000;
	sram_mem[73473] = 16'b0000000000000000;
	sram_mem[73474] = 16'b0000000000000000;
	sram_mem[73475] = 16'b0000000000000000;
	sram_mem[73476] = 16'b0000000000000000;
	sram_mem[73477] = 16'b0000000000000000;
	sram_mem[73478] = 16'b0000000000000000;
	sram_mem[73479] = 16'b0000000000000000;
	sram_mem[73480] = 16'b0000000000000000;
	sram_mem[73481] = 16'b0000000000000000;
	sram_mem[73482] = 16'b0000000000000000;
	sram_mem[73483] = 16'b0000000000000000;
	sram_mem[73484] = 16'b0000000000000000;
	sram_mem[73485] = 16'b0000000000000000;
	sram_mem[73486] = 16'b0000000000000000;
	sram_mem[73487] = 16'b0000000000000000;
	sram_mem[73488] = 16'b0000000000000000;
	sram_mem[73489] = 16'b0000000000000000;
	sram_mem[73490] = 16'b0000000000000000;
	sram_mem[73491] = 16'b0000000000000000;
	sram_mem[73492] = 16'b0000000000000000;
	sram_mem[73493] = 16'b0000000000000000;
	sram_mem[73494] = 16'b0000000000000000;
	sram_mem[73495] = 16'b0000000000000000;
	sram_mem[73496] = 16'b0000000000000000;
	sram_mem[73497] = 16'b0000000000000000;
	sram_mem[73498] = 16'b0000000000000000;
	sram_mem[73499] = 16'b0000000000000000;
	sram_mem[73500] = 16'b0000000000000000;
	sram_mem[73501] = 16'b0000000000000000;
	sram_mem[73502] = 16'b0000000000000000;
	sram_mem[73503] = 16'b0000000000000000;
	sram_mem[73504] = 16'b0000000000000000;
	sram_mem[73505] = 16'b0000000000000000;
	sram_mem[73506] = 16'b0000000000000000;
	sram_mem[73507] = 16'b0000000000000000;
	sram_mem[73508] = 16'b0000000000000000;
	sram_mem[73509] = 16'b0000000000000000;
	sram_mem[73510] = 16'b0000000000000000;
	sram_mem[73511] = 16'b0000000000000000;
	sram_mem[73512] = 16'b0000000000000000;
	sram_mem[73513] = 16'b0000000000000000;
	sram_mem[73514] = 16'b0000000000000000;
	sram_mem[73515] = 16'b0000000000000000;
	sram_mem[73516] = 16'b0000000000000000;
	sram_mem[73517] = 16'b0000000000000000;
	sram_mem[73518] = 16'b0000000000000000;
	sram_mem[73519] = 16'b0000000000000000;
	sram_mem[73520] = 16'b0000000000000000;
	sram_mem[73521] = 16'b0000000000000000;
	sram_mem[73522] = 16'b0000000000000000;
	sram_mem[73523] = 16'b0000000000000000;
	sram_mem[73524] = 16'b0000000000000000;
	sram_mem[73525] = 16'b0000000000000000;
	sram_mem[73526] = 16'b0000000000000000;
	sram_mem[73527] = 16'b0000000000000000;
	sram_mem[73528] = 16'b0000000000000000;
	sram_mem[73529] = 16'b0000000000000000;
	sram_mem[73530] = 16'b0000000000000000;
	sram_mem[73531] = 16'b0000000000000000;
	sram_mem[73532] = 16'b0000000000000000;
	sram_mem[73533] = 16'b0000000000000000;
	sram_mem[73534] = 16'b0000000000000000;
	sram_mem[73535] = 16'b0000000000000000;
	sram_mem[73536] = 16'b0000000000000000;
	sram_mem[73537] = 16'b0000000000000000;
	sram_mem[73538] = 16'b0000000000000000;
	sram_mem[73539] = 16'b0000000000000000;
	sram_mem[73540] = 16'b0000000000000000;
	sram_mem[73541] = 16'b0000000000000000;
	sram_mem[73542] = 16'b0000000000000000;
	sram_mem[73543] = 16'b0000000000000000;
	sram_mem[73544] = 16'b0000000000000000;
	sram_mem[73545] = 16'b0000000000000000;
	sram_mem[73546] = 16'b0000000000000000;
	sram_mem[73547] = 16'b0000000000000000;
	sram_mem[73548] = 16'b0000000000000000;
	sram_mem[73549] = 16'b0000000000000000;
	sram_mem[73550] = 16'b0000000000000000;
	sram_mem[73551] = 16'b0000000000000000;
	sram_mem[73552] = 16'b0000000000000000;
	sram_mem[73553] = 16'b0000000000000000;
	sram_mem[73554] = 16'b0000000000000000;
	sram_mem[73555] = 16'b0000000000000000;
	sram_mem[73556] = 16'b0000000000000000;
	sram_mem[73557] = 16'b0000000000000000;
	sram_mem[73558] = 16'b0000000000000000;
	sram_mem[73559] = 16'b0000000000000000;
	sram_mem[73560] = 16'b0000000000000000;
	sram_mem[73561] = 16'b0000000000000000;
	sram_mem[73562] = 16'b0000000000000000;
	sram_mem[73563] = 16'b0000000000000000;
	sram_mem[73564] = 16'b0000000000000000;
	sram_mem[73565] = 16'b0000000000000000;
	sram_mem[73566] = 16'b0000000000000000;
	sram_mem[73567] = 16'b0000000000000000;
	sram_mem[73568] = 16'b0000000000000000;
	sram_mem[73569] = 16'b0000000000000000;
	sram_mem[73570] = 16'b0000000000000000;
	sram_mem[73571] = 16'b0000000000000000;
	sram_mem[73572] = 16'b0000000000000000;
	sram_mem[73573] = 16'b0000000000000000;
	sram_mem[73574] = 16'b0000000000000000;
	sram_mem[73575] = 16'b0000000000000000;
	sram_mem[73576] = 16'b0000000000000000;
	sram_mem[73577] = 16'b0000000000000000;
	sram_mem[73578] = 16'b0000000000000000;
	sram_mem[73579] = 16'b0000000000000000;
	sram_mem[73580] = 16'b0000000000000000;
	sram_mem[73581] = 16'b0000000000000000;
	sram_mem[73582] = 16'b0000000000000000;
	sram_mem[73583] = 16'b0000000000000000;
	sram_mem[73584] = 16'b0000000000000000;
	sram_mem[73585] = 16'b0000000000000000;
	sram_mem[73586] = 16'b0000000000000000;
	sram_mem[73587] = 16'b0000000000000000;
	sram_mem[73588] = 16'b0000000000000000;
	sram_mem[73589] = 16'b0000000000000000;
	sram_mem[73590] = 16'b0000000000000000;
	sram_mem[73591] = 16'b0000000000000000;
	sram_mem[73592] = 16'b0000000000000000;
	sram_mem[73593] = 16'b0000000000000000;
	sram_mem[73594] = 16'b0000000000000000;
	sram_mem[73595] = 16'b0000000000000000;
	sram_mem[73596] = 16'b0000000000000000;
	sram_mem[73597] = 16'b0000000000000000;
	sram_mem[73598] = 16'b0000000000000000;
	sram_mem[73599] = 16'b0000000000000000;
	sram_mem[73600] = 16'b0000000000000000;
	sram_mem[73601] = 16'b0000000000000000;
	sram_mem[73602] = 16'b0000000000000000;
	sram_mem[73603] = 16'b0000000000000000;
	sram_mem[73604] = 16'b0000000000000000;
	sram_mem[73605] = 16'b0000000000000000;
	sram_mem[73606] = 16'b0000000000000000;
	sram_mem[73607] = 16'b0000000000000000;
	sram_mem[73608] = 16'b0000000000000000;
	sram_mem[73609] = 16'b0000000000000000;
	sram_mem[73610] = 16'b0000000000000000;
	sram_mem[73611] = 16'b0000000000000000;
	sram_mem[73612] = 16'b0000000000000000;
	sram_mem[73613] = 16'b0000000000000000;
	sram_mem[73614] = 16'b0000000000000000;
	sram_mem[73615] = 16'b0000000000000000;
	sram_mem[73616] = 16'b0000000000000000;
	sram_mem[73617] = 16'b0000000000000000;
	sram_mem[73618] = 16'b0000000000000000;
	sram_mem[73619] = 16'b0000000000000000;
	sram_mem[73620] = 16'b0000000000000000;
	sram_mem[73621] = 16'b0000000000000000;
	sram_mem[73622] = 16'b0000000000000000;
	sram_mem[73623] = 16'b0000000000000000;
	sram_mem[73624] = 16'b0000000000000000;
	sram_mem[73625] = 16'b0000000000000000;
	sram_mem[73626] = 16'b0000000000000000;
	sram_mem[73627] = 16'b0000000000000000;
	sram_mem[73628] = 16'b0000000000000000;
	sram_mem[73629] = 16'b0000000000000000;
	sram_mem[73630] = 16'b0000000000000000;
	sram_mem[73631] = 16'b0000000000000000;
	sram_mem[73632] = 16'b0000000000000000;
	sram_mem[73633] = 16'b0000000000000000;
	sram_mem[73634] = 16'b0000000000000000;
	sram_mem[73635] = 16'b0000000000000000;
	sram_mem[73636] = 16'b0000000000000000;
	sram_mem[73637] = 16'b0000000000000000;
	sram_mem[73638] = 16'b0000000000000000;
	sram_mem[73639] = 16'b0000000000000000;
	sram_mem[73640] = 16'b0000000000000000;
	sram_mem[73641] = 16'b0000000000000000;
	sram_mem[73642] = 16'b0000000000000000;
	sram_mem[73643] = 16'b0000000000000000;
	sram_mem[73644] = 16'b0000000000000000;
	sram_mem[73645] = 16'b0000000000000000;
	sram_mem[73646] = 16'b0000000000000000;
	sram_mem[73647] = 16'b0000000000000000;
	sram_mem[73648] = 16'b0000000000000000;
	sram_mem[73649] = 16'b0000000000000000;
	sram_mem[73650] = 16'b0000000000000000;
	sram_mem[73651] = 16'b0000000000000000;
	sram_mem[73652] = 16'b0000000000000000;
	sram_mem[73653] = 16'b0000000000000000;
	sram_mem[73654] = 16'b0000000000000000;
	sram_mem[73655] = 16'b0000000000000000;
	sram_mem[73656] = 16'b0000000000000000;
	sram_mem[73657] = 16'b0000000000000000;
	sram_mem[73658] = 16'b0000000000000000;
	sram_mem[73659] = 16'b0000000000000000;
	sram_mem[73660] = 16'b0000000000000000;
	sram_mem[73661] = 16'b0000000000000000;
	sram_mem[73662] = 16'b0000000000000000;
	sram_mem[73663] = 16'b0000000000000000;
	sram_mem[73664] = 16'b0000000000000000;
	sram_mem[73665] = 16'b0000000000000000;
	sram_mem[73666] = 16'b0000000000000000;
	sram_mem[73667] = 16'b0000000000000000;
	sram_mem[73668] = 16'b0000000000000000;
	sram_mem[73669] = 16'b0000000000000000;
	sram_mem[73670] = 16'b0000000000000000;
	sram_mem[73671] = 16'b0000000000000000;
	sram_mem[73672] = 16'b0000000000000000;
	sram_mem[73673] = 16'b0000000000000000;
	sram_mem[73674] = 16'b0000000000000000;
	sram_mem[73675] = 16'b0000000000000000;
	sram_mem[73676] = 16'b0000000000000000;
	sram_mem[73677] = 16'b0000000000000000;
	sram_mem[73678] = 16'b0000000000000000;
	sram_mem[73679] = 16'b0000000000000000;
	sram_mem[73680] = 16'b0000000000000000;
	sram_mem[73681] = 16'b0000000000000000;
	sram_mem[73682] = 16'b0000000000000000;
	sram_mem[73683] = 16'b0000000000000000;
	sram_mem[73684] = 16'b0000000000000000;
	sram_mem[73685] = 16'b0000000000000000;
	sram_mem[73686] = 16'b0000000000000000;
	sram_mem[73687] = 16'b0000000000000000;
	sram_mem[73688] = 16'b0000000000000000;
	sram_mem[73689] = 16'b0000000000000000;
	sram_mem[73690] = 16'b0000000000000000;
	sram_mem[73691] = 16'b0000000000000000;
	sram_mem[73692] = 16'b0000000000000000;
	sram_mem[73693] = 16'b0000000000000000;
	sram_mem[73694] = 16'b0000000000000000;
	sram_mem[73695] = 16'b0000000000000000;
	sram_mem[73696] = 16'b0000000000000000;
	sram_mem[73697] = 16'b0000000000000000;
	sram_mem[73698] = 16'b0000000000000000;
	sram_mem[73699] = 16'b0000000000000000;
	sram_mem[73700] = 16'b0000000000000000;
	sram_mem[73701] = 16'b0000000000000000;
	sram_mem[73702] = 16'b0000000000000000;
	sram_mem[73703] = 16'b0000000000000000;
	sram_mem[73704] = 16'b0000000000000000;
	sram_mem[73705] = 16'b0000000000000000;
	sram_mem[73706] = 16'b0000000000000000;
	sram_mem[73707] = 16'b0000000000000000;
	sram_mem[73708] = 16'b0000000000000000;
	sram_mem[73709] = 16'b0000000000000000;
	sram_mem[73710] = 16'b0000000000000000;
	sram_mem[73711] = 16'b0000000000000000;
	sram_mem[73712] = 16'b0000000000000000;
	sram_mem[73713] = 16'b0000000000000000;
	sram_mem[73714] = 16'b0000000000000000;
	sram_mem[73715] = 16'b0000000000000000;
	sram_mem[73716] = 16'b0000000000000000;
	sram_mem[73717] = 16'b0000000000000000;
	sram_mem[73718] = 16'b0000000000000000;
	sram_mem[73719] = 16'b0000000000000000;
	sram_mem[73720] = 16'b0000000000000000;
	sram_mem[73721] = 16'b0000000000000000;
	sram_mem[73722] = 16'b0000000000000000;
	sram_mem[73723] = 16'b0000000000000000;
	sram_mem[73724] = 16'b0000000000000000;
	sram_mem[73725] = 16'b0000000000000000;
	sram_mem[73726] = 16'b0000000000000000;
	sram_mem[73727] = 16'b0000000000000000;
	sram_mem[73728] = 16'b0000000000000000;
	sram_mem[73729] = 16'b0000000000000000;
	sram_mem[73730] = 16'b0000000000000000;
	sram_mem[73731] = 16'b0000000000000000;
	sram_mem[73732] = 16'b0000000000000000;
	sram_mem[73733] = 16'b0000000000000000;
	sram_mem[73734] = 16'b0000000000000000;
	sram_mem[73735] = 16'b0000000000000000;
	sram_mem[73736] = 16'b0000000000000000;
	sram_mem[73737] = 16'b0000000000000000;
	sram_mem[73738] = 16'b0000000000000000;
	sram_mem[73739] = 16'b0000000000000000;
	sram_mem[73740] = 16'b0000000000000000;
	sram_mem[73741] = 16'b0000000000000000;
	sram_mem[73742] = 16'b0000000000000000;
	sram_mem[73743] = 16'b0000000000000000;
	sram_mem[73744] = 16'b0000000000000000;
	sram_mem[73745] = 16'b0000000000000000;
	sram_mem[73746] = 16'b0000000000000000;
	sram_mem[73747] = 16'b0000000000000000;
	sram_mem[73748] = 16'b0000000000000000;
	sram_mem[73749] = 16'b0000000000000000;
	sram_mem[73750] = 16'b0000000000000000;
	sram_mem[73751] = 16'b0000000000000000;
	sram_mem[73752] = 16'b0000000000000000;
	sram_mem[73753] = 16'b0000000000000000;
	sram_mem[73754] = 16'b0000000000000000;
	sram_mem[73755] = 16'b0000000000000000;
	sram_mem[73756] = 16'b0000000000000000;
	sram_mem[73757] = 16'b0000000000000000;
	sram_mem[73758] = 16'b0000000000000000;
	sram_mem[73759] = 16'b0000000000000000;
	sram_mem[73760] = 16'b0000000000000000;
	sram_mem[73761] = 16'b0000000000000000;
	sram_mem[73762] = 16'b0000000000000000;
	sram_mem[73763] = 16'b0000000000000000;
	sram_mem[73764] = 16'b0000000000000000;
	sram_mem[73765] = 16'b0000000000000000;
	sram_mem[73766] = 16'b0000000000000000;
	sram_mem[73767] = 16'b0000000000000000;
	sram_mem[73768] = 16'b0000000000000000;
	sram_mem[73769] = 16'b0000000000000000;
	sram_mem[73770] = 16'b0000000000000000;
	sram_mem[73771] = 16'b0000000000000000;
	sram_mem[73772] = 16'b0000000000000000;
	sram_mem[73773] = 16'b0000000000000000;
	sram_mem[73774] = 16'b0000000000000000;
	sram_mem[73775] = 16'b0000000000000000;
	sram_mem[73776] = 16'b0000000000000000;
	sram_mem[73777] = 16'b0000000000000000;
	sram_mem[73778] = 16'b0000000000000000;
	sram_mem[73779] = 16'b0000000000000000;
	sram_mem[73780] = 16'b0000000000000000;
	sram_mem[73781] = 16'b0000000000000000;
	sram_mem[73782] = 16'b0000000000000000;
	sram_mem[73783] = 16'b0000000000000000;
	sram_mem[73784] = 16'b0000000000000000;
	sram_mem[73785] = 16'b0000000000000000;
	sram_mem[73786] = 16'b0000000000000000;
	sram_mem[73787] = 16'b0000000000000000;
	sram_mem[73788] = 16'b0000000000000000;
	sram_mem[73789] = 16'b0000000000000000;
	sram_mem[73790] = 16'b0000000000000000;
	sram_mem[73791] = 16'b0000000000000000;
	sram_mem[73792] = 16'b0000000000000000;
	sram_mem[73793] = 16'b0000000000000000;
	sram_mem[73794] = 16'b0000000000000000;
	sram_mem[73795] = 16'b0000000000000000;
	sram_mem[73796] = 16'b0000000000000000;
	sram_mem[73797] = 16'b0000000000000000;
	sram_mem[73798] = 16'b0000000000000000;
	sram_mem[73799] = 16'b0000000000000000;
	sram_mem[73800] = 16'b0000000000000000;
	sram_mem[73801] = 16'b0000000000000000;
	sram_mem[73802] = 16'b0000000000000000;
	sram_mem[73803] = 16'b0000000000000000;
	sram_mem[73804] = 16'b0000000000000000;
	sram_mem[73805] = 16'b0000000000000000;
	sram_mem[73806] = 16'b0000000000000000;
	sram_mem[73807] = 16'b0000000000000000;
	sram_mem[73808] = 16'b0000000000000000;
	sram_mem[73809] = 16'b0000000000000000;
	sram_mem[73810] = 16'b0000000000000000;
	sram_mem[73811] = 16'b0000000000000000;
	sram_mem[73812] = 16'b0000000000000000;
	sram_mem[73813] = 16'b0000000000000000;
	sram_mem[73814] = 16'b0000000000000000;
	sram_mem[73815] = 16'b0000000000000000;
	sram_mem[73816] = 16'b0000000000000000;
	sram_mem[73817] = 16'b0000000000000000;
	sram_mem[73818] = 16'b0000000000000000;
	sram_mem[73819] = 16'b0000000000000000;
	sram_mem[73820] = 16'b0000000000000000;
	sram_mem[73821] = 16'b0000000000000000;
	sram_mem[73822] = 16'b0000000000000000;
	sram_mem[73823] = 16'b0000000000000000;
	sram_mem[73824] = 16'b0000000000000000;
	sram_mem[73825] = 16'b0000000000000000;
	sram_mem[73826] = 16'b0000000000000000;
	sram_mem[73827] = 16'b0000000000000000;
	sram_mem[73828] = 16'b0000000000000000;
	sram_mem[73829] = 16'b0000000000000000;
	sram_mem[73830] = 16'b0000000000000000;
	sram_mem[73831] = 16'b0000000000000000;
	sram_mem[73832] = 16'b0000000000000000;
	sram_mem[73833] = 16'b0000000000000000;
	sram_mem[73834] = 16'b0000000000000000;
	sram_mem[73835] = 16'b0000000000000000;
	sram_mem[73836] = 16'b0000000000000000;
	sram_mem[73837] = 16'b0000000000000000;
	sram_mem[73838] = 16'b0000000000000000;
	sram_mem[73839] = 16'b0000000000000000;
	sram_mem[73840] = 16'b0000000000000000;
	sram_mem[73841] = 16'b0000000000000000;
	sram_mem[73842] = 16'b0000000000000000;
	sram_mem[73843] = 16'b0000000000000000;
	sram_mem[73844] = 16'b0000000000000000;
	sram_mem[73845] = 16'b0000000000000000;
	sram_mem[73846] = 16'b0000000000000000;
	sram_mem[73847] = 16'b0000000000000000;
	sram_mem[73848] = 16'b0000000000000000;
	sram_mem[73849] = 16'b0000000000000000;
	sram_mem[73850] = 16'b0000000000000000;
	sram_mem[73851] = 16'b0000000000000000;
	sram_mem[73852] = 16'b0000000000000000;
	sram_mem[73853] = 16'b0000000000000000;
	sram_mem[73854] = 16'b0000000000000000;
	sram_mem[73855] = 16'b0000000000000000;
	sram_mem[73856] = 16'b0000000000000000;
	sram_mem[73857] = 16'b0000000000000000;
	sram_mem[73858] = 16'b0000000000000000;
	sram_mem[73859] = 16'b0000000000000000;
	sram_mem[73860] = 16'b0000000000000000;
	sram_mem[73861] = 16'b0000000000000000;
	sram_mem[73862] = 16'b0000000000000000;
	sram_mem[73863] = 16'b0000000000000000;
	sram_mem[73864] = 16'b0000000000000000;
	sram_mem[73865] = 16'b0000000000000000;
	sram_mem[73866] = 16'b0000000000000000;
	sram_mem[73867] = 16'b0000000000000000;
	sram_mem[73868] = 16'b0000000000000000;
	sram_mem[73869] = 16'b0000000000000000;
	sram_mem[73870] = 16'b0000000000000000;
	sram_mem[73871] = 16'b0000000000000000;
	sram_mem[73872] = 16'b0000000000000000;
	sram_mem[73873] = 16'b0000000000000000;
	sram_mem[73874] = 16'b0000000000000000;
	sram_mem[73875] = 16'b0000000000000000;
	sram_mem[73876] = 16'b0000000000000000;
	sram_mem[73877] = 16'b0000000000000000;
	sram_mem[73878] = 16'b0000000000000000;
	sram_mem[73879] = 16'b0000000000000000;
	sram_mem[73880] = 16'b0000000000000000;
	sram_mem[73881] = 16'b0000000000000000;
	sram_mem[73882] = 16'b0000000000000000;
	sram_mem[73883] = 16'b0000000000000000;
	sram_mem[73884] = 16'b0000000000000000;
	sram_mem[73885] = 16'b0000000000000000;
	sram_mem[73886] = 16'b0000000000000000;
	sram_mem[73887] = 16'b0000000000000000;
	sram_mem[73888] = 16'b0000000000000000;
	sram_mem[73889] = 16'b0000000000000000;
	sram_mem[73890] = 16'b0000000000000000;
	sram_mem[73891] = 16'b0000000000000000;
	sram_mem[73892] = 16'b0000000000000000;
	sram_mem[73893] = 16'b0000000000000000;
	sram_mem[73894] = 16'b0000000000000000;
	sram_mem[73895] = 16'b0000000000000000;
	sram_mem[73896] = 16'b0000000000000000;
	sram_mem[73897] = 16'b0000000000000000;
	sram_mem[73898] = 16'b0000000000000000;
	sram_mem[73899] = 16'b0000000000000000;
	sram_mem[73900] = 16'b0000000000000000;
	sram_mem[73901] = 16'b0000000000000000;
	sram_mem[73902] = 16'b0000000000000000;
	sram_mem[73903] = 16'b0000000000000000;
	sram_mem[73904] = 16'b0000000000000000;
	sram_mem[73905] = 16'b0000000000000000;
	sram_mem[73906] = 16'b0000000000000000;
	sram_mem[73907] = 16'b0000000000000000;
	sram_mem[73908] = 16'b0000000000000000;
	sram_mem[73909] = 16'b0000000000000000;
	sram_mem[73910] = 16'b0000000000000000;
	sram_mem[73911] = 16'b0000000000000000;
	sram_mem[73912] = 16'b0000000000000000;
	sram_mem[73913] = 16'b0000000000000000;
	sram_mem[73914] = 16'b0000000000000000;
	sram_mem[73915] = 16'b0000000000000000;
	sram_mem[73916] = 16'b0000000000000000;
	sram_mem[73917] = 16'b0000000000000000;
	sram_mem[73918] = 16'b0000000000000000;
	sram_mem[73919] = 16'b0000000000000000;
	sram_mem[73920] = 16'b0000000000000000;
	sram_mem[73921] = 16'b0000000000000000;
	sram_mem[73922] = 16'b0000000000000000;
	sram_mem[73923] = 16'b0000000000000000;
	sram_mem[73924] = 16'b0000000000000000;
	sram_mem[73925] = 16'b0000000000000000;
	sram_mem[73926] = 16'b0000000000000000;
	sram_mem[73927] = 16'b0000000000000000;
	sram_mem[73928] = 16'b0000000000000000;
	sram_mem[73929] = 16'b0000000000000000;
	sram_mem[73930] = 16'b0000000000000000;
	sram_mem[73931] = 16'b0000000000000000;
	sram_mem[73932] = 16'b0000000000000000;
	sram_mem[73933] = 16'b0000000000000000;
	sram_mem[73934] = 16'b0000000000000000;
	sram_mem[73935] = 16'b0000000000000000;
	sram_mem[73936] = 16'b0000000000000000;
	sram_mem[73937] = 16'b0000000000000000;
	sram_mem[73938] = 16'b0000000000000000;
	sram_mem[73939] = 16'b0000000000000000;
	sram_mem[73940] = 16'b0000000000000000;
	sram_mem[73941] = 16'b0000000000000000;
	sram_mem[73942] = 16'b0000000000000000;
	sram_mem[73943] = 16'b0000000000000000;
	sram_mem[73944] = 16'b0000000000000000;
	sram_mem[73945] = 16'b0000000000000000;
	sram_mem[73946] = 16'b0000000000000000;
	sram_mem[73947] = 16'b0000000000000000;
	sram_mem[73948] = 16'b0000000000000000;
	sram_mem[73949] = 16'b0000000000000000;
	sram_mem[73950] = 16'b0000000000000000;
	sram_mem[73951] = 16'b0000000000000000;
	sram_mem[73952] = 16'b0000000000000000;
	sram_mem[73953] = 16'b0000000000000000;
	sram_mem[73954] = 16'b0000000000000000;
	sram_mem[73955] = 16'b0000000000000000;
	sram_mem[73956] = 16'b0000000000000000;
	sram_mem[73957] = 16'b0000000000000000;
	sram_mem[73958] = 16'b0000000000000000;
	sram_mem[73959] = 16'b0000000000000000;
	sram_mem[73960] = 16'b0000000000000000;
	sram_mem[73961] = 16'b0000000000000000;
	sram_mem[73962] = 16'b0000000000000000;
	sram_mem[73963] = 16'b0000000000000000;
	sram_mem[73964] = 16'b0000000000000000;
	sram_mem[73965] = 16'b0000000000000000;
	sram_mem[73966] = 16'b0000000000000000;
	sram_mem[73967] = 16'b0000000000000000;
	sram_mem[73968] = 16'b0000000000000000;
	sram_mem[73969] = 16'b0000000000000000;
	sram_mem[73970] = 16'b0000000000000000;
	sram_mem[73971] = 16'b0000000000000000;
	sram_mem[73972] = 16'b0000000000000000;
	sram_mem[73973] = 16'b0000000000000000;
	sram_mem[73974] = 16'b0000000000000000;
	sram_mem[73975] = 16'b0000000000000000;
	sram_mem[73976] = 16'b0000000000000000;
	sram_mem[73977] = 16'b0000000000000000;
	sram_mem[73978] = 16'b0000000000000000;
	sram_mem[73979] = 16'b0000000000000000;
	sram_mem[73980] = 16'b0000000000000000;
	sram_mem[73981] = 16'b0000000000000000;
	sram_mem[73982] = 16'b0000000000000000;
	sram_mem[73983] = 16'b0000000000000000;
	sram_mem[73984] = 16'b0000000000000000;
	sram_mem[73985] = 16'b0000000000000000;
	sram_mem[73986] = 16'b0000000000000000;
	sram_mem[73987] = 16'b0000000000000000;
	sram_mem[73988] = 16'b0000000000000000;
	sram_mem[73989] = 16'b0000000000000000;
	sram_mem[73990] = 16'b0000000000000000;
	sram_mem[73991] = 16'b0000000000000000;
	sram_mem[73992] = 16'b0000000000000000;
	sram_mem[73993] = 16'b0000000000000000;
	sram_mem[73994] = 16'b0000000000000000;
	sram_mem[73995] = 16'b0000000000000000;
	sram_mem[73996] = 16'b0000000000000000;
	sram_mem[73997] = 16'b0000000000000000;
	sram_mem[73998] = 16'b0000000000000000;
	sram_mem[73999] = 16'b0000000000000000;
	sram_mem[74000] = 16'b0000000000000000;
	sram_mem[74001] = 16'b0000000000000000;
	sram_mem[74002] = 16'b0000000000000000;
	sram_mem[74003] = 16'b0000000000000000;
	sram_mem[74004] = 16'b0000000000000000;
	sram_mem[74005] = 16'b0000000000000000;
	sram_mem[74006] = 16'b0000000000000000;
	sram_mem[74007] = 16'b0000000000000000;
	sram_mem[74008] = 16'b0000000000000000;
	sram_mem[74009] = 16'b0000000000000000;
	sram_mem[74010] = 16'b0000000000000000;
	sram_mem[74011] = 16'b0000000000000000;
	sram_mem[74012] = 16'b0000000000000000;
	sram_mem[74013] = 16'b0000000000000000;
	sram_mem[74014] = 16'b0000000000000000;
	sram_mem[74015] = 16'b0000000000000000;
	sram_mem[74016] = 16'b0000000000000000;
	sram_mem[74017] = 16'b0000000000000000;
	sram_mem[74018] = 16'b0000000000000000;
	sram_mem[74019] = 16'b0000000000000000;
	sram_mem[74020] = 16'b0000000000000000;
	sram_mem[74021] = 16'b0000000000000000;
	sram_mem[74022] = 16'b0000000000000000;
	sram_mem[74023] = 16'b0000000000000000;
	sram_mem[74024] = 16'b0000000000000000;
	sram_mem[74025] = 16'b0000000000000000;
	sram_mem[74026] = 16'b0000000000000000;
	sram_mem[74027] = 16'b0000000000000000;
	sram_mem[74028] = 16'b0000000000000000;
	sram_mem[74029] = 16'b0000000000000000;
	sram_mem[74030] = 16'b0000000000000000;
	sram_mem[74031] = 16'b0000000000000000;
	sram_mem[74032] = 16'b0000000000000000;
	sram_mem[74033] = 16'b0000000000000000;
	sram_mem[74034] = 16'b0000000000000000;
	sram_mem[74035] = 16'b0000000000000000;
	sram_mem[74036] = 16'b0000000000000000;
	sram_mem[74037] = 16'b0000000000000000;
	sram_mem[74038] = 16'b0000000000000000;
	sram_mem[74039] = 16'b0000000000000000;
	sram_mem[74040] = 16'b0000000000000000;
	sram_mem[74041] = 16'b0000000000000000;
	sram_mem[74042] = 16'b0000000000000000;
	sram_mem[74043] = 16'b0000000000000000;
	sram_mem[74044] = 16'b0000000000000000;
	sram_mem[74045] = 16'b0000000000000000;
	sram_mem[74046] = 16'b0000000000000000;
	sram_mem[74047] = 16'b0000000000000000;
	sram_mem[74048] = 16'b0000000000000000;
	sram_mem[74049] = 16'b0000000000000000;
	sram_mem[74050] = 16'b0000000000000000;
	sram_mem[74051] = 16'b0000000000000000;
	sram_mem[74052] = 16'b0000000000000000;
	sram_mem[74053] = 16'b0000000000000000;
	sram_mem[74054] = 16'b0000000000000000;
	sram_mem[74055] = 16'b0000000000000000;
	sram_mem[74056] = 16'b0000000000000000;
	sram_mem[74057] = 16'b0000000000000000;
	sram_mem[74058] = 16'b0000000000000000;
	sram_mem[74059] = 16'b0000000000000000;
	sram_mem[74060] = 16'b0000000000000000;
	sram_mem[74061] = 16'b0000000000000000;
	sram_mem[74062] = 16'b0000000000000000;
	sram_mem[74063] = 16'b0000000000000000;
	sram_mem[74064] = 16'b0000000000000000;
	sram_mem[74065] = 16'b0000000000000000;
	sram_mem[74066] = 16'b0000000000000000;
	sram_mem[74067] = 16'b0000000000000000;
	sram_mem[74068] = 16'b0000000000000000;
	sram_mem[74069] = 16'b0000000000000000;
	sram_mem[74070] = 16'b0000000000000000;
	sram_mem[74071] = 16'b0000000000000000;
	sram_mem[74072] = 16'b0000000000000000;
	sram_mem[74073] = 16'b0000000000000000;
	sram_mem[74074] = 16'b0000000000000000;
	sram_mem[74075] = 16'b0000000000000000;
	sram_mem[74076] = 16'b0000000000000000;
	sram_mem[74077] = 16'b0000000000000000;
	sram_mem[74078] = 16'b0000000000000000;
	sram_mem[74079] = 16'b0000000000000000;
	sram_mem[74080] = 16'b0000000000000000;
	sram_mem[74081] = 16'b0000000000000000;
	sram_mem[74082] = 16'b0000000000000000;
	sram_mem[74083] = 16'b0000000000000000;
	sram_mem[74084] = 16'b0000000000000000;
	sram_mem[74085] = 16'b0000000000000000;
	sram_mem[74086] = 16'b0000000000000000;
	sram_mem[74087] = 16'b0000000000000000;
	sram_mem[74088] = 16'b0000000000000000;
	sram_mem[74089] = 16'b0000000000000000;
	sram_mem[74090] = 16'b0000000000000000;
	sram_mem[74091] = 16'b0000000000000000;
	sram_mem[74092] = 16'b0000000000000000;
	sram_mem[74093] = 16'b0000000000000000;
	sram_mem[74094] = 16'b0000000000000000;
	sram_mem[74095] = 16'b0000000000000000;
	sram_mem[74096] = 16'b0000000000000000;
	sram_mem[74097] = 16'b0000000000000000;
	sram_mem[74098] = 16'b0000000000000000;
	sram_mem[74099] = 16'b0000000000000000;
	sram_mem[74100] = 16'b0000000000000000;
	sram_mem[74101] = 16'b0000000000000000;
	sram_mem[74102] = 16'b0000000000000000;
	sram_mem[74103] = 16'b0000000000000000;
	sram_mem[74104] = 16'b0000000000000000;
	sram_mem[74105] = 16'b0000000000000000;
	sram_mem[74106] = 16'b0000000000000000;
	sram_mem[74107] = 16'b0000000000000000;
	sram_mem[74108] = 16'b0000000000000000;
	sram_mem[74109] = 16'b0000000000000000;
	sram_mem[74110] = 16'b0000000000000000;
	sram_mem[74111] = 16'b0000000000000000;
	sram_mem[74112] = 16'b0000000000000000;
	sram_mem[74113] = 16'b0000000000000000;
	sram_mem[74114] = 16'b0000000000000000;
	sram_mem[74115] = 16'b0000000000000000;
	sram_mem[74116] = 16'b0000000000000000;
	sram_mem[74117] = 16'b0000000000000000;
	sram_mem[74118] = 16'b0000000000000000;
	sram_mem[74119] = 16'b0000000000000000;
	sram_mem[74120] = 16'b0000000000000000;
	sram_mem[74121] = 16'b0000000000000000;
	sram_mem[74122] = 16'b0000000000000000;
	sram_mem[74123] = 16'b0000000000000000;
	sram_mem[74124] = 16'b0000000000000000;
	sram_mem[74125] = 16'b0000000000000000;
	sram_mem[74126] = 16'b0000000000000000;
	sram_mem[74127] = 16'b0000000000000000;
	sram_mem[74128] = 16'b0000000000000000;
	sram_mem[74129] = 16'b0000000000000000;
	sram_mem[74130] = 16'b0000000000000000;
	sram_mem[74131] = 16'b0000000000000000;
	sram_mem[74132] = 16'b0000000000000000;
	sram_mem[74133] = 16'b0000000000000000;
	sram_mem[74134] = 16'b0000000000000000;
	sram_mem[74135] = 16'b0000000000000000;
	sram_mem[74136] = 16'b0000000000000000;
	sram_mem[74137] = 16'b0000000000000000;
	sram_mem[74138] = 16'b0000000000000000;
	sram_mem[74139] = 16'b0000000000000000;
	sram_mem[74140] = 16'b0000000000000000;
	sram_mem[74141] = 16'b0000000000000000;
	sram_mem[74142] = 16'b0000000000000000;
	sram_mem[74143] = 16'b0000000000000000;
	sram_mem[74144] = 16'b0000000000000000;
	sram_mem[74145] = 16'b0000000000000000;
	sram_mem[74146] = 16'b0000000000000000;
	sram_mem[74147] = 16'b0000000000000000;
	sram_mem[74148] = 16'b0000000000000000;
	sram_mem[74149] = 16'b0000000000000000;
	sram_mem[74150] = 16'b0000000000000000;
	sram_mem[74151] = 16'b0000000000000000;
	sram_mem[74152] = 16'b0000000000000000;
	sram_mem[74153] = 16'b0000000000000000;
	sram_mem[74154] = 16'b0000000000000000;
	sram_mem[74155] = 16'b0000000000000000;
	sram_mem[74156] = 16'b0000000000000000;
	sram_mem[74157] = 16'b0000000000000000;
	sram_mem[74158] = 16'b0000000000000000;
	sram_mem[74159] = 16'b0000000000000000;
	sram_mem[74160] = 16'b0000000000000000;
	sram_mem[74161] = 16'b0000000000000000;
	sram_mem[74162] = 16'b0000000000000000;
	sram_mem[74163] = 16'b0000000000000000;
	sram_mem[74164] = 16'b0000000000000000;
	sram_mem[74165] = 16'b0000000000000000;
	sram_mem[74166] = 16'b0000000000000000;
	sram_mem[74167] = 16'b0000000000000000;
	sram_mem[74168] = 16'b0000000000000000;
	sram_mem[74169] = 16'b0000000000000000;
	sram_mem[74170] = 16'b0000000000000000;
	sram_mem[74171] = 16'b0000000000000000;
	sram_mem[74172] = 16'b0000000000000000;
	sram_mem[74173] = 16'b0000000000000000;
	sram_mem[74174] = 16'b0000000000000000;
	sram_mem[74175] = 16'b0000000000000000;
	sram_mem[74176] = 16'b0000000000000000;
	sram_mem[74177] = 16'b0000000000000000;
	sram_mem[74178] = 16'b0000000000000000;
	sram_mem[74179] = 16'b0000000000000000;
	sram_mem[74180] = 16'b0000000000000000;
	sram_mem[74181] = 16'b0000000000000000;
	sram_mem[74182] = 16'b0000000000000000;
	sram_mem[74183] = 16'b0000000000000000;
	sram_mem[74184] = 16'b0000000000000000;
	sram_mem[74185] = 16'b0000000000000000;
	sram_mem[74186] = 16'b0000000000000000;
	sram_mem[74187] = 16'b0000000000000000;
	sram_mem[74188] = 16'b0000000000000000;
	sram_mem[74189] = 16'b0000000000000000;
	sram_mem[74190] = 16'b0000000000000000;
	sram_mem[74191] = 16'b0000000000000000;
	sram_mem[74192] = 16'b0000000000000000;
	sram_mem[74193] = 16'b0000000000000000;
	sram_mem[74194] = 16'b0000000000000000;
	sram_mem[74195] = 16'b0000000000000000;
	sram_mem[74196] = 16'b0000000000000000;
	sram_mem[74197] = 16'b0000000000000000;
	sram_mem[74198] = 16'b0000000000000000;
	sram_mem[74199] = 16'b0000000000000000;
	sram_mem[74200] = 16'b0000000000000000;
	sram_mem[74201] = 16'b0000000000000000;
	sram_mem[74202] = 16'b0000000000000000;
	sram_mem[74203] = 16'b0000000000000000;
	sram_mem[74204] = 16'b0000000000000000;
	sram_mem[74205] = 16'b0000000000000000;
	sram_mem[74206] = 16'b0000000000000000;
	sram_mem[74207] = 16'b0000000000000000;
	sram_mem[74208] = 16'b0000000000000000;
	sram_mem[74209] = 16'b0000000000000000;
	sram_mem[74210] = 16'b0000000000000000;
	sram_mem[74211] = 16'b0000000000000000;
	sram_mem[74212] = 16'b0000000000000000;
	sram_mem[74213] = 16'b0000000000000000;
	sram_mem[74214] = 16'b0000000000000000;
	sram_mem[74215] = 16'b0000000000000000;
	sram_mem[74216] = 16'b0000000000000000;
	sram_mem[74217] = 16'b0000000000000000;
	sram_mem[74218] = 16'b0000000000000000;
	sram_mem[74219] = 16'b0000000000000000;
	sram_mem[74220] = 16'b0000000000000000;
	sram_mem[74221] = 16'b0000000000000000;
	sram_mem[74222] = 16'b0000000000000000;
	sram_mem[74223] = 16'b0000000000000000;
	sram_mem[74224] = 16'b0000000000000000;
	sram_mem[74225] = 16'b0000000000000000;
	sram_mem[74226] = 16'b0000000000000000;
	sram_mem[74227] = 16'b0000000000000000;
	sram_mem[74228] = 16'b0000000000000000;
	sram_mem[74229] = 16'b0000000000000000;
	sram_mem[74230] = 16'b0000000000000000;
	sram_mem[74231] = 16'b0000000000000000;
	sram_mem[74232] = 16'b0000000000000000;
	sram_mem[74233] = 16'b0000000000000000;
	sram_mem[74234] = 16'b0000000000000000;
	sram_mem[74235] = 16'b0000000000000000;
	sram_mem[74236] = 16'b0000000000000000;
	sram_mem[74237] = 16'b0000000000000000;
	sram_mem[74238] = 16'b0000000000000000;
	sram_mem[74239] = 16'b0000000000000000;
	sram_mem[74240] = 16'b0000000000000000;
	sram_mem[74241] = 16'b0000000000000000;
	sram_mem[74242] = 16'b0000000000000000;
	sram_mem[74243] = 16'b0000000000000000;
	sram_mem[74244] = 16'b0000000000000000;
	sram_mem[74245] = 16'b0000000000000000;
	sram_mem[74246] = 16'b0000000000000000;
	sram_mem[74247] = 16'b0000000000000000;
	sram_mem[74248] = 16'b0000000000000000;
	sram_mem[74249] = 16'b0000000000000000;
	sram_mem[74250] = 16'b0000000000000000;
	sram_mem[74251] = 16'b0000000000000000;
	sram_mem[74252] = 16'b0000000000000000;
	sram_mem[74253] = 16'b0000000000000000;
	sram_mem[74254] = 16'b0000000000000000;
	sram_mem[74255] = 16'b0000000000000000;
	sram_mem[74256] = 16'b0000000000000000;
	sram_mem[74257] = 16'b0000000000000000;
	sram_mem[74258] = 16'b0000000000000000;
	sram_mem[74259] = 16'b0000000000000000;
	sram_mem[74260] = 16'b0000000000000000;
	sram_mem[74261] = 16'b0000000000000000;
	sram_mem[74262] = 16'b0000000000000000;
	sram_mem[74263] = 16'b0000000000000000;
	sram_mem[74264] = 16'b0000000000000000;
	sram_mem[74265] = 16'b0000000000000000;
	sram_mem[74266] = 16'b0000000000000000;
	sram_mem[74267] = 16'b0000000000000000;
	sram_mem[74268] = 16'b0000000000000000;
	sram_mem[74269] = 16'b0000000000000000;
	sram_mem[74270] = 16'b0000000000000000;
	sram_mem[74271] = 16'b0000000000000000;
	sram_mem[74272] = 16'b0000000000000000;
	sram_mem[74273] = 16'b0000000000000000;
	sram_mem[74274] = 16'b0000000000000000;
	sram_mem[74275] = 16'b0000000000000000;
	sram_mem[74276] = 16'b0000000000000000;
	sram_mem[74277] = 16'b0000000000000000;
	sram_mem[74278] = 16'b0000000000000000;
	sram_mem[74279] = 16'b0000000000000000;
	sram_mem[74280] = 16'b0000000000000000;
	sram_mem[74281] = 16'b0000000000000000;
	sram_mem[74282] = 16'b0000000000000000;
	sram_mem[74283] = 16'b0000000000000000;
	sram_mem[74284] = 16'b0000000000000000;
	sram_mem[74285] = 16'b0000000000000000;
	sram_mem[74286] = 16'b0000000000000000;
	sram_mem[74287] = 16'b0000000000000000;
	sram_mem[74288] = 16'b0000000000000000;
	sram_mem[74289] = 16'b0000000000000000;
	sram_mem[74290] = 16'b0000000000000000;
	sram_mem[74291] = 16'b0000000000000000;
	sram_mem[74292] = 16'b0000000000000000;
	sram_mem[74293] = 16'b0000000000000000;
	sram_mem[74294] = 16'b0000000000000000;
	sram_mem[74295] = 16'b0000000000000000;
	sram_mem[74296] = 16'b0000000000000000;
	sram_mem[74297] = 16'b0000000000000000;
	sram_mem[74298] = 16'b0000000000000000;
	sram_mem[74299] = 16'b0000000000000000;
	sram_mem[74300] = 16'b0000000000000000;
	sram_mem[74301] = 16'b0000000000000000;
	sram_mem[74302] = 16'b0000000000000000;
	sram_mem[74303] = 16'b0000000000000000;
	sram_mem[74304] = 16'b0000000000000000;
	sram_mem[74305] = 16'b0000000000000000;
	sram_mem[74306] = 16'b0000000000000000;
	sram_mem[74307] = 16'b0000000000000000;
	sram_mem[74308] = 16'b0000000000000000;
	sram_mem[74309] = 16'b0000000000000000;
	sram_mem[74310] = 16'b0000000000000000;
	sram_mem[74311] = 16'b0000000000000000;
	sram_mem[74312] = 16'b0000000000000000;
	sram_mem[74313] = 16'b0000000000000000;
	sram_mem[74314] = 16'b0000000000000000;
	sram_mem[74315] = 16'b0000000000000000;
	sram_mem[74316] = 16'b0000000000000000;
	sram_mem[74317] = 16'b0000000000000000;
	sram_mem[74318] = 16'b0000000000000000;
	sram_mem[74319] = 16'b0000000000000000;
	sram_mem[74320] = 16'b0000000000000000;
	sram_mem[74321] = 16'b0000000000000000;
	sram_mem[74322] = 16'b0000000000000000;
	sram_mem[74323] = 16'b0000000000000000;
	sram_mem[74324] = 16'b0000000000000000;
	sram_mem[74325] = 16'b0000000000000000;
	sram_mem[74326] = 16'b0000000000000000;
	sram_mem[74327] = 16'b0000000000000000;
	sram_mem[74328] = 16'b0000000000000000;
	sram_mem[74329] = 16'b0000000000000000;
	sram_mem[74330] = 16'b0000000000000000;
	sram_mem[74331] = 16'b0000000000000000;
	sram_mem[74332] = 16'b0000000000000000;
	sram_mem[74333] = 16'b0000000000000000;
	sram_mem[74334] = 16'b0000000000000000;
	sram_mem[74335] = 16'b0000000000000000;
	sram_mem[74336] = 16'b0000000000000000;
	sram_mem[74337] = 16'b0000000000000000;
	sram_mem[74338] = 16'b0000000000000000;
	sram_mem[74339] = 16'b0000000000000000;
	sram_mem[74340] = 16'b0000000000000000;
	sram_mem[74341] = 16'b0000000000000000;
	sram_mem[74342] = 16'b0000000000000000;
	sram_mem[74343] = 16'b0000000000000000;
	sram_mem[74344] = 16'b0000000000000000;
	sram_mem[74345] = 16'b0000000000000000;
	sram_mem[74346] = 16'b0000000000000000;
	sram_mem[74347] = 16'b0000000000000000;
	sram_mem[74348] = 16'b0000000000000000;
	sram_mem[74349] = 16'b0000000000000000;
	sram_mem[74350] = 16'b0000000000000000;
	sram_mem[74351] = 16'b0000000000000000;
	sram_mem[74352] = 16'b0000000000000000;
	sram_mem[74353] = 16'b0000000000000000;
	sram_mem[74354] = 16'b0000000000000000;
	sram_mem[74355] = 16'b0000000000000000;
	sram_mem[74356] = 16'b0000000000000000;
	sram_mem[74357] = 16'b0000000000000000;
	sram_mem[74358] = 16'b0000000000000000;
	sram_mem[74359] = 16'b0000000000000000;
	sram_mem[74360] = 16'b0000000000000000;
	sram_mem[74361] = 16'b0000000000000000;
	sram_mem[74362] = 16'b0000000000000000;
	sram_mem[74363] = 16'b0000000000000000;
	sram_mem[74364] = 16'b0000000000000000;
	sram_mem[74365] = 16'b0000000000000000;
	sram_mem[74366] = 16'b0000000000000000;
	sram_mem[74367] = 16'b0000000000000000;
	sram_mem[74368] = 16'b0000000000000000;
	sram_mem[74369] = 16'b0000000000000000;
	sram_mem[74370] = 16'b0000000000000000;
	sram_mem[74371] = 16'b0000000000000000;
	sram_mem[74372] = 16'b0000000000000000;
	sram_mem[74373] = 16'b0000000000000000;
	sram_mem[74374] = 16'b0000000000000000;
	sram_mem[74375] = 16'b0000000000000000;
	sram_mem[74376] = 16'b0000000000000000;
	sram_mem[74377] = 16'b0000000000000000;
	sram_mem[74378] = 16'b0000000000000000;
	sram_mem[74379] = 16'b0000000000000000;
	sram_mem[74380] = 16'b0000000000000000;
	sram_mem[74381] = 16'b0000000000000000;
	sram_mem[74382] = 16'b0000000000000000;
	sram_mem[74383] = 16'b0000000000000000;
	sram_mem[74384] = 16'b0000000000000000;
	sram_mem[74385] = 16'b0000000000000000;
	sram_mem[74386] = 16'b0000000000000000;
	sram_mem[74387] = 16'b0000000000000000;
	sram_mem[74388] = 16'b0000000000000000;
	sram_mem[74389] = 16'b0000000000000000;
	sram_mem[74390] = 16'b0000000000000000;
	sram_mem[74391] = 16'b0000000000000000;
	sram_mem[74392] = 16'b0000000000000000;
	sram_mem[74393] = 16'b0000000000000000;
	sram_mem[74394] = 16'b0000000000000000;
	sram_mem[74395] = 16'b0000000000000000;
	sram_mem[74396] = 16'b0000000000000000;
	sram_mem[74397] = 16'b0000000000000000;
	sram_mem[74398] = 16'b0000000000000000;
	sram_mem[74399] = 16'b0000000000000000;
	sram_mem[74400] = 16'b0000000000000000;
	sram_mem[74401] = 16'b0000000000000000;
	sram_mem[74402] = 16'b0000000000000000;
	sram_mem[74403] = 16'b0000000000000000;
	sram_mem[74404] = 16'b0000000000000000;
	sram_mem[74405] = 16'b0000000000000000;
	sram_mem[74406] = 16'b0000000000000000;
	sram_mem[74407] = 16'b0000000000000000;
	sram_mem[74408] = 16'b0000000000000000;
	sram_mem[74409] = 16'b0000000000000000;
	sram_mem[74410] = 16'b0000000000000000;
	sram_mem[74411] = 16'b0000000000000000;
	sram_mem[74412] = 16'b0000000000000000;
	sram_mem[74413] = 16'b0000000000000000;
	sram_mem[74414] = 16'b0000000000000000;
	sram_mem[74415] = 16'b0000000000000000;
	sram_mem[74416] = 16'b0000000000000000;
	sram_mem[74417] = 16'b0000000000000000;
	sram_mem[74418] = 16'b0000000000000000;
	sram_mem[74419] = 16'b0000000000000000;
	sram_mem[74420] = 16'b0000000000000000;
	sram_mem[74421] = 16'b0000000000000000;
	sram_mem[74422] = 16'b0000000000000000;
	sram_mem[74423] = 16'b0000000000000000;
	sram_mem[74424] = 16'b0000000000000000;
	sram_mem[74425] = 16'b0000000000000000;
	sram_mem[74426] = 16'b0000000000000000;
	sram_mem[74427] = 16'b0000000000000000;
	sram_mem[74428] = 16'b0000000000000000;
	sram_mem[74429] = 16'b0000000000000000;
	sram_mem[74430] = 16'b0000000000000000;
	sram_mem[74431] = 16'b0000000000000000;
	sram_mem[74432] = 16'b0000000000000000;
	sram_mem[74433] = 16'b0000000000000000;
	sram_mem[74434] = 16'b0000000000000000;
	sram_mem[74435] = 16'b0000000000000000;
	sram_mem[74436] = 16'b0000000000000000;
	sram_mem[74437] = 16'b0000000000000000;
	sram_mem[74438] = 16'b0000000000000000;
	sram_mem[74439] = 16'b0000000000000000;
	sram_mem[74440] = 16'b0000000000000000;
	sram_mem[74441] = 16'b0000000000000000;
	sram_mem[74442] = 16'b0000000000000000;
	sram_mem[74443] = 16'b0000000000000000;
	sram_mem[74444] = 16'b0000000000000000;
	sram_mem[74445] = 16'b0000000000000000;
	sram_mem[74446] = 16'b0000000000000000;
	sram_mem[74447] = 16'b0000000000000000;
	sram_mem[74448] = 16'b0000000000000000;
	sram_mem[74449] = 16'b0000000000000000;
	sram_mem[74450] = 16'b0000000000000000;
	sram_mem[74451] = 16'b0000000000000000;
	sram_mem[74452] = 16'b0000000000000000;
	sram_mem[74453] = 16'b0000000000000000;
	sram_mem[74454] = 16'b0000000000000000;
	sram_mem[74455] = 16'b0000000000000000;
	sram_mem[74456] = 16'b0000000000000000;
	sram_mem[74457] = 16'b0000000000000000;
	sram_mem[74458] = 16'b0000000000000000;
	sram_mem[74459] = 16'b0000000000000000;
	sram_mem[74460] = 16'b0000000000000000;
	sram_mem[74461] = 16'b0000000000000000;
	sram_mem[74462] = 16'b0000000000000000;
	sram_mem[74463] = 16'b0000000000000000;
	sram_mem[74464] = 16'b0000000000000000;
	sram_mem[74465] = 16'b0000000000000000;
	sram_mem[74466] = 16'b0000000000000000;
	sram_mem[74467] = 16'b0000000000000000;
	sram_mem[74468] = 16'b0000000000000000;
	sram_mem[74469] = 16'b0000000000000000;
	sram_mem[74470] = 16'b0000000000000000;
	sram_mem[74471] = 16'b0000000000000000;
	sram_mem[74472] = 16'b0000000000000000;
	sram_mem[74473] = 16'b0000000000000000;
	sram_mem[74474] = 16'b0000000000000000;
	sram_mem[74475] = 16'b0000000000000000;
	sram_mem[74476] = 16'b0000000000000000;
	sram_mem[74477] = 16'b0000000000000000;
	sram_mem[74478] = 16'b0000000000000000;
	sram_mem[74479] = 16'b0000000000000000;
	sram_mem[74480] = 16'b0000000000000000;
	sram_mem[74481] = 16'b0000000000000000;
	sram_mem[74482] = 16'b0000000000000000;
	sram_mem[74483] = 16'b0000000000000000;
	sram_mem[74484] = 16'b0000000000000000;
	sram_mem[74485] = 16'b0000000000000000;
	sram_mem[74486] = 16'b0000000000000000;
	sram_mem[74487] = 16'b0000000000000000;
	sram_mem[74488] = 16'b0000000000000000;
	sram_mem[74489] = 16'b0000000000000000;
	sram_mem[74490] = 16'b0000000000000000;
	sram_mem[74491] = 16'b0000000000000000;
	sram_mem[74492] = 16'b0000000000000000;
	sram_mem[74493] = 16'b0000000000000000;
	sram_mem[74494] = 16'b0000000000000000;
	sram_mem[74495] = 16'b0000000000000000;
	sram_mem[74496] = 16'b0000000000000000;
	sram_mem[74497] = 16'b0000000000000000;
	sram_mem[74498] = 16'b0000000000000000;
	sram_mem[74499] = 16'b0000000000000000;
	sram_mem[74500] = 16'b0000000000000000;
	sram_mem[74501] = 16'b0000000000000000;
	sram_mem[74502] = 16'b0000000000000000;
	sram_mem[74503] = 16'b0000000000000000;
	sram_mem[74504] = 16'b0000000000000000;
	sram_mem[74505] = 16'b0000000000000000;
	sram_mem[74506] = 16'b0000000000000000;
	sram_mem[74507] = 16'b0000000000000000;
	sram_mem[74508] = 16'b0000000000000000;
	sram_mem[74509] = 16'b0000000000000000;
	sram_mem[74510] = 16'b0000000000000000;
	sram_mem[74511] = 16'b0000000000000000;
	sram_mem[74512] = 16'b0000000000000000;
	sram_mem[74513] = 16'b0000000000000000;
	sram_mem[74514] = 16'b0000000000000000;
	sram_mem[74515] = 16'b0000000000000000;
	sram_mem[74516] = 16'b0000000000000000;
	sram_mem[74517] = 16'b0000000000000000;
	sram_mem[74518] = 16'b0000000000000000;
	sram_mem[74519] = 16'b0000000000000000;
	sram_mem[74520] = 16'b0000000000000000;
	sram_mem[74521] = 16'b0000000000000000;
	sram_mem[74522] = 16'b0000000000000000;
	sram_mem[74523] = 16'b0000000000000000;
	sram_mem[74524] = 16'b0000000000000000;
	sram_mem[74525] = 16'b0000000000000000;
	sram_mem[74526] = 16'b0000000000000000;
	sram_mem[74527] = 16'b0000000000000000;
	sram_mem[74528] = 16'b0000000000000000;
	sram_mem[74529] = 16'b0000000000000000;
	sram_mem[74530] = 16'b0000000000000000;
	sram_mem[74531] = 16'b0000000000000000;
	sram_mem[74532] = 16'b0000000000000000;
	sram_mem[74533] = 16'b0000000000000000;
	sram_mem[74534] = 16'b0000000000000000;
	sram_mem[74535] = 16'b0000000000000000;
	sram_mem[74536] = 16'b0000000000000000;
	sram_mem[74537] = 16'b0000000000000000;
	sram_mem[74538] = 16'b0000000000000000;
	sram_mem[74539] = 16'b0000000000000000;
	sram_mem[74540] = 16'b0000000000000000;
	sram_mem[74541] = 16'b0000000000000000;
	sram_mem[74542] = 16'b0000000000000000;
	sram_mem[74543] = 16'b0000000000000000;
	sram_mem[74544] = 16'b0000000000000000;
	sram_mem[74545] = 16'b0000000000000000;
	sram_mem[74546] = 16'b0000000000000000;
	sram_mem[74547] = 16'b0000000000000000;
	sram_mem[74548] = 16'b0000000000000000;
	sram_mem[74549] = 16'b0000000000000000;
	sram_mem[74550] = 16'b0000000000000000;
	sram_mem[74551] = 16'b0000000000000000;
	sram_mem[74552] = 16'b0000000000000000;
	sram_mem[74553] = 16'b0000000000000000;
	sram_mem[74554] = 16'b0000000000000000;
	sram_mem[74555] = 16'b0000000000000000;
	sram_mem[74556] = 16'b0000000000000000;
	sram_mem[74557] = 16'b0000000000000000;
	sram_mem[74558] = 16'b0000000000000000;
	sram_mem[74559] = 16'b0000000000000000;
	sram_mem[74560] = 16'b0000000000000000;
	sram_mem[74561] = 16'b0000000000000000;
	sram_mem[74562] = 16'b0000000000000000;
	sram_mem[74563] = 16'b0000000000000000;
	sram_mem[74564] = 16'b0000000000000000;
	sram_mem[74565] = 16'b0000000000000000;
	sram_mem[74566] = 16'b0000000000000000;
	sram_mem[74567] = 16'b0000000000000000;
	sram_mem[74568] = 16'b0000000000000000;
	sram_mem[74569] = 16'b0000000000000000;
	sram_mem[74570] = 16'b0000000000000000;
	sram_mem[74571] = 16'b0000000000000000;
	sram_mem[74572] = 16'b0000000000000000;
	sram_mem[74573] = 16'b0000000000000000;
	sram_mem[74574] = 16'b0000000000000000;
	sram_mem[74575] = 16'b0000000000000000;
	sram_mem[74576] = 16'b0000000000000000;
	sram_mem[74577] = 16'b0000000000000000;
	sram_mem[74578] = 16'b0000000000000000;
	sram_mem[74579] = 16'b0000000000000000;
	sram_mem[74580] = 16'b0000000000000000;
	sram_mem[74581] = 16'b0000000000000000;
	sram_mem[74582] = 16'b0000000000000000;
	sram_mem[74583] = 16'b0000000000000000;
	sram_mem[74584] = 16'b0000000000000000;
	sram_mem[74585] = 16'b0000000000000000;
	sram_mem[74586] = 16'b0000000000000000;
	sram_mem[74587] = 16'b0000000000000000;
	sram_mem[74588] = 16'b0000000000000000;
	sram_mem[74589] = 16'b0000000000000000;
	sram_mem[74590] = 16'b0000000000000000;
	sram_mem[74591] = 16'b0000000000000000;
	sram_mem[74592] = 16'b0000000000000000;
	sram_mem[74593] = 16'b0000000000000000;
	sram_mem[74594] = 16'b0000000000000000;
	sram_mem[74595] = 16'b0000000000000000;
	sram_mem[74596] = 16'b0000000000000000;
	sram_mem[74597] = 16'b0000000000000000;
	sram_mem[74598] = 16'b0000000000000000;
	sram_mem[74599] = 16'b0000000000000000;
	sram_mem[74600] = 16'b0000000000000000;
	sram_mem[74601] = 16'b0000000000000000;
	sram_mem[74602] = 16'b0000000000000000;
	sram_mem[74603] = 16'b0000000000000000;
	sram_mem[74604] = 16'b0000000000000000;
	sram_mem[74605] = 16'b0000000000000000;
	sram_mem[74606] = 16'b0000000000000000;
	sram_mem[74607] = 16'b0000000000000000;
	sram_mem[74608] = 16'b0000000000000000;
	sram_mem[74609] = 16'b0000000000000000;
	sram_mem[74610] = 16'b0000000000000000;
	sram_mem[74611] = 16'b0000000000000000;
	sram_mem[74612] = 16'b0000000000000000;
	sram_mem[74613] = 16'b0000000000000000;
	sram_mem[74614] = 16'b0000000000000000;
	sram_mem[74615] = 16'b0000000000000000;
	sram_mem[74616] = 16'b0000000000000000;
	sram_mem[74617] = 16'b0000000000000000;
	sram_mem[74618] = 16'b0000000000000000;
	sram_mem[74619] = 16'b0000000000000000;
	sram_mem[74620] = 16'b0000000000000000;
	sram_mem[74621] = 16'b0000000000000000;
	sram_mem[74622] = 16'b0000000000000000;
	sram_mem[74623] = 16'b0000000000000000;
	sram_mem[74624] = 16'b0000000000000000;
	sram_mem[74625] = 16'b0000000000000000;
	sram_mem[74626] = 16'b0000000000000000;
	sram_mem[74627] = 16'b0000000000000000;
	sram_mem[74628] = 16'b0000000000000000;
	sram_mem[74629] = 16'b0000000000000000;
	sram_mem[74630] = 16'b0000000000000000;
	sram_mem[74631] = 16'b0000000000000000;
	sram_mem[74632] = 16'b0000000000000000;
	sram_mem[74633] = 16'b0000000000000000;
	sram_mem[74634] = 16'b0000000000000000;
	sram_mem[74635] = 16'b0000000000000000;
	sram_mem[74636] = 16'b0000000000000000;
	sram_mem[74637] = 16'b0000000000000000;
	sram_mem[74638] = 16'b0000000000000000;
	sram_mem[74639] = 16'b0000000000000000;
	sram_mem[74640] = 16'b0000000000000000;
	sram_mem[74641] = 16'b0000000000000000;
	sram_mem[74642] = 16'b0000000000000000;
	sram_mem[74643] = 16'b0000000000000000;
	sram_mem[74644] = 16'b0000000000000000;
	sram_mem[74645] = 16'b0000000000000000;
	sram_mem[74646] = 16'b0000000000000000;
	sram_mem[74647] = 16'b0000000000000000;
	sram_mem[74648] = 16'b0000000000000000;
	sram_mem[74649] = 16'b0000000000000000;
	sram_mem[74650] = 16'b0000000000000000;
	sram_mem[74651] = 16'b0000000000000000;
	sram_mem[74652] = 16'b0000000000000000;
	sram_mem[74653] = 16'b0000000000000000;
	sram_mem[74654] = 16'b0000000000000000;
	sram_mem[74655] = 16'b0000000000000000;
	sram_mem[74656] = 16'b0000000000000000;
	sram_mem[74657] = 16'b0000000000000000;
	sram_mem[74658] = 16'b0000000000000000;
	sram_mem[74659] = 16'b0000000000000000;
	sram_mem[74660] = 16'b0000000000000000;
	sram_mem[74661] = 16'b0000000000000000;
	sram_mem[74662] = 16'b0000000000000000;
	sram_mem[74663] = 16'b0000000000000000;
	sram_mem[74664] = 16'b0000000000000000;
	sram_mem[74665] = 16'b0000000000000000;
	sram_mem[74666] = 16'b0000000000000000;
	sram_mem[74667] = 16'b0000000000000000;
	sram_mem[74668] = 16'b0000000000000000;
	sram_mem[74669] = 16'b0000000000000000;
	sram_mem[74670] = 16'b0000000000000000;
	sram_mem[74671] = 16'b0000000000000000;
	sram_mem[74672] = 16'b0000000000000000;
	sram_mem[74673] = 16'b0000000000000000;
	sram_mem[74674] = 16'b0000000000000000;
	sram_mem[74675] = 16'b0000000000000000;
	sram_mem[74676] = 16'b0000000000000000;
	sram_mem[74677] = 16'b0000000000000000;
	sram_mem[74678] = 16'b0000000000000000;
	sram_mem[74679] = 16'b0000000000000000;
	sram_mem[74680] = 16'b0000000000000000;
	sram_mem[74681] = 16'b0000000000000000;
	sram_mem[74682] = 16'b0000000000000000;
	sram_mem[74683] = 16'b0000000000000000;
	sram_mem[74684] = 16'b0000000000000000;
	sram_mem[74685] = 16'b0000000000000000;
	sram_mem[74686] = 16'b0000000000000000;
	sram_mem[74687] = 16'b0000000000000000;
	sram_mem[74688] = 16'b0000000000000000;
	sram_mem[74689] = 16'b0000000000000000;
	sram_mem[74690] = 16'b0000000000000000;
	sram_mem[74691] = 16'b0000000000000000;
	sram_mem[74692] = 16'b0000000000000000;
	sram_mem[74693] = 16'b0000000000000000;
	sram_mem[74694] = 16'b0000000000000000;
	sram_mem[74695] = 16'b0000000000000000;
	sram_mem[74696] = 16'b0000000000000000;
	sram_mem[74697] = 16'b0000000000000000;
	sram_mem[74698] = 16'b0000000000000000;
	sram_mem[74699] = 16'b0000000000000000;
	sram_mem[74700] = 16'b0000000000000000;
	sram_mem[74701] = 16'b0000000000000000;
	sram_mem[74702] = 16'b0000000000000000;
	sram_mem[74703] = 16'b0000000000000000;
	sram_mem[74704] = 16'b0000000000000000;
	sram_mem[74705] = 16'b0000000000000000;
	sram_mem[74706] = 16'b0000000000000000;
	sram_mem[74707] = 16'b0000000000000000;
	sram_mem[74708] = 16'b0000000000000000;
	sram_mem[74709] = 16'b0000000000000000;
	sram_mem[74710] = 16'b0000000000000000;
	sram_mem[74711] = 16'b0000000000000000;
	sram_mem[74712] = 16'b0000000000000000;
	sram_mem[74713] = 16'b0000000000000000;
	sram_mem[74714] = 16'b0000000000000000;
	sram_mem[74715] = 16'b0000000000000000;
	sram_mem[74716] = 16'b0000000000000000;
	sram_mem[74717] = 16'b0000000000000000;
	sram_mem[74718] = 16'b0000000000000000;
	sram_mem[74719] = 16'b0000000000000000;
	sram_mem[74720] = 16'b0000000000000000;
	sram_mem[74721] = 16'b0000000000000000;
	sram_mem[74722] = 16'b0000000000000000;
	sram_mem[74723] = 16'b0000000000000000;
	sram_mem[74724] = 16'b0000000000000000;
	sram_mem[74725] = 16'b0000000000000000;
	sram_mem[74726] = 16'b0000000000000000;
	sram_mem[74727] = 16'b0000000000000000;
	sram_mem[74728] = 16'b0000000000000000;
	sram_mem[74729] = 16'b0000000000000000;
	sram_mem[74730] = 16'b0000000000000000;
	sram_mem[74731] = 16'b0000000000000000;
	sram_mem[74732] = 16'b0000000000000000;
	sram_mem[74733] = 16'b0000000000000000;
	sram_mem[74734] = 16'b0000000000000000;
	sram_mem[74735] = 16'b0000000000000000;
	sram_mem[74736] = 16'b0000000000000000;
	sram_mem[74737] = 16'b0000000000000000;
	sram_mem[74738] = 16'b0000000000000000;
	sram_mem[74739] = 16'b0000000000000000;
	sram_mem[74740] = 16'b0000000000000000;
	sram_mem[74741] = 16'b0000000000000000;
	sram_mem[74742] = 16'b0000000000000000;
	sram_mem[74743] = 16'b0000000000000000;
	sram_mem[74744] = 16'b0000000000000000;
	sram_mem[74745] = 16'b0000000000000000;
	sram_mem[74746] = 16'b0000000000000000;
	sram_mem[74747] = 16'b0000000000000000;
	sram_mem[74748] = 16'b0000000000000000;
	sram_mem[74749] = 16'b0000000000000000;
	sram_mem[74750] = 16'b0000000000000000;
	sram_mem[74751] = 16'b0000000000000000;
	sram_mem[74752] = 16'b0000000000000000;
	sram_mem[74753] = 16'b0000000000000000;
	sram_mem[74754] = 16'b0000000000000000;
	sram_mem[74755] = 16'b0000000000000000;
	sram_mem[74756] = 16'b0000000000000000;
	sram_mem[74757] = 16'b0000000000000000;
	sram_mem[74758] = 16'b0000000000000000;
	sram_mem[74759] = 16'b0000000000000000;
	sram_mem[74760] = 16'b0000000000000000;
	sram_mem[74761] = 16'b0000000000000000;
	sram_mem[74762] = 16'b0000000000000000;
	sram_mem[74763] = 16'b0000000000000000;
	sram_mem[74764] = 16'b0000000000000000;
	sram_mem[74765] = 16'b0000000000000000;
	sram_mem[74766] = 16'b0000000000000000;
	sram_mem[74767] = 16'b0000000000000000;
	sram_mem[74768] = 16'b0000000000000000;
	sram_mem[74769] = 16'b0000000000000000;
	sram_mem[74770] = 16'b0000000000000000;
	sram_mem[74771] = 16'b0000000000000000;
	sram_mem[74772] = 16'b0000000000000000;
	sram_mem[74773] = 16'b0000000000000000;
	sram_mem[74774] = 16'b0000000000000000;
	sram_mem[74775] = 16'b0000000000000000;
	sram_mem[74776] = 16'b0000000000000000;
	sram_mem[74777] = 16'b0000000000000000;
	sram_mem[74778] = 16'b0000000000000000;
	sram_mem[74779] = 16'b0000000000000000;
	sram_mem[74780] = 16'b0000000000000000;
	sram_mem[74781] = 16'b0000000000000000;
	sram_mem[74782] = 16'b0000000000000000;
	sram_mem[74783] = 16'b0000000000000000;
	sram_mem[74784] = 16'b0000000000000000;
	sram_mem[74785] = 16'b0000000000000000;
	sram_mem[74786] = 16'b0000000000000000;
	sram_mem[74787] = 16'b0000000000000000;
	sram_mem[74788] = 16'b0000000000000000;
	sram_mem[74789] = 16'b0000000000000000;
	sram_mem[74790] = 16'b0000000000000000;
	sram_mem[74791] = 16'b0000000000000000;
	sram_mem[74792] = 16'b0000000000000000;
	sram_mem[74793] = 16'b0000000000000000;
	sram_mem[74794] = 16'b0000000000000000;
	sram_mem[74795] = 16'b0000000000000000;
	sram_mem[74796] = 16'b0000000000000000;
	sram_mem[74797] = 16'b0000000000000000;
	sram_mem[74798] = 16'b0000000000000000;
	sram_mem[74799] = 16'b0000000000000000;
	sram_mem[74800] = 16'b0000000000000000;
	sram_mem[74801] = 16'b0000000000000000;
	sram_mem[74802] = 16'b0000000000000000;
	sram_mem[74803] = 16'b0000000000000000;
	sram_mem[74804] = 16'b0000000000000000;
	sram_mem[74805] = 16'b0000000000000000;
	sram_mem[74806] = 16'b0000000000000000;
	sram_mem[74807] = 16'b0000000000000000;
	sram_mem[74808] = 16'b0000000000000000;
	sram_mem[74809] = 16'b0000000000000000;
	sram_mem[74810] = 16'b0000000000000000;
	sram_mem[74811] = 16'b0000000000000000;
	sram_mem[74812] = 16'b0000000000000000;
	sram_mem[74813] = 16'b0000000000000000;
	sram_mem[74814] = 16'b0000000000000000;
	sram_mem[74815] = 16'b0000000000000000;
	sram_mem[74816] = 16'b0000000000000000;
	sram_mem[74817] = 16'b0000000000000000;
	sram_mem[74818] = 16'b0000000000000000;
	sram_mem[74819] = 16'b0000000000000000;
	sram_mem[74820] = 16'b0000000000000000;
	sram_mem[74821] = 16'b0000000000000000;
	sram_mem[74822] = 16'b0000000000000000;
	sram_mem[74823] = 16'b0000000000000000;
	sram_mem[74824] = 16'b0000000000000000;
	sram_mem[74825] = 16'b0000000000000000;
	sram_mem[74826] = 16'b0000000000000000;
	sram_mem[74827] = 16'b0000000000000000;
	sram_mem[74828] = 16'b0000000000000000;
	sram_mem[74829] = 16'b0000000000000000;
	sram_mem[74830] = 16'b0000000000000000;
	sram_mem[74831] = 16'b0000000000000000;
	sram_mem[74832] = 16'b0000000000000000;
	sram_mem[74833] = 16'b0000000000000000;
	sram_mem[74834] = 16'b0000000000000000;
	sram_mem[74835] = 16'b0000000000000000;
	sram_mem[74836] = 16'b0000000000000000;
	sram_mem[74837] = 16'b0000000000000000;
	sram_mem[74838] = 16'b0000000000000000;
	sram_mem[74839] = 16'b0000000000000000;
	sram_mem[74840] = 16'b0000000000000000;
	sram_mem[74841] = 16'b0000000000000000;
	sram_mem[74842] = 16'b0000000000000000;
	sram_mem[74843] = 16'b0000000000000000;
	sram_mem[74844] = 16'b0000000000000000;
	sram_mem[74845] = 16'b0000000000000000;
	sram_mem[74846] = 16'b0000000000000000;
	sram_mem[74847] = 16'b0000000000000000;
	sram_mem[74848] = 16'b0000000000000000;
	sram_mem[74849] = 16'b0000000000000000;
	sram_mem[74850] = 16'b0000000000000000;
	sram_mem[74851] = 16'b0000000000000000;
	sram_mem[74852] = 16'b0000000000000000;
	sram_mem[74853] = 16'b0000000000000000;
	sram_mem[74854] = 16'b0000000000000000;
	sram_mem[74855] = 16'b0000000000000000;
	sram_mem[74856] = 16'b0000000000000000;
	sram_mem[74857] = 16'b0000000000000000;
	sram_mem[74858] = 16'b0000000000000000;
	sram_mem[74859] = 16'b0000000000000000;
	sram_mem[74860] = 16'b0000000000000000;
	sram_mem[74861] = 16'b0000000000000000;
	sram_mem[74862] = 16'b0000000000000000;
	sram_mem[74863] = 16'b0000000000000000;
	sram_mem[74864] = 16'b0000000000000000;
	sram_mem[74865] = 16'b0000000000000000;
	sram_mem[74866] = 16'b0000000000000000;
	sram_mem[74867] = 16'b0000000000000000;
	sram_mem[74868] = 16'b0000000000000000;
	sram_mem[74869] = 16'b0000000000000000;
	sram_mem[74870] = 16'b0000000000000000;
	sram_mem[74871] = 16'b0000000000000000;
	sram_mem[74872] = 16'b0000000000000000;
	sram_mem[74873] = 16'b0000000000000000;
	sram_mem[74874] = 16'b0000000000000000;
	sram_mem[74875] = 16'b0000000000000000;
	sram_mem[74876] = 16'b0000000000000000;
	sram_mem[74877] = 16'b0000000000000000;
	sram_mem[74878] = 16'b0000000000000000;
	sram_mem[74879] = 16'b0000000000000000;
	sram_mem[74880] = 16'b0000000000000000;
	sram_mem[74881] = 16'b0000000000000000;
	sram_mem[74882] = 16'b0000000000000000;
	sram_mem[74883] = 16'b0000000000000000;
	sram_mem[74884] = 16'b0000000000000000;
	sram_mem[74885] = 16'b0000000000000000;
	sram_mem[74886] = 16'b0000000000000000;
	sram_mem[74887] = 16'b0000000000000000;
	sram_mem[74888] = 16'b0000000000000000;
	sram_mem[74889] = 16'b0000000000000000;
	sram_mem[74890] = 16'b0000000000000000;
	sram_mem[74891] = 16'b0000000000000000;
	sram_mem[74892] = 16'b0000000000000000;
	sram_mem[74893] = 16'b0000000000000000;
	sram_mem[74894] = 16'b0000000000000000;
	sram_mem[74895] = 16'b0000000000000000;
	sram_mem[74896] = 16'b0000000000000000;
	sram_mem[74897] = 16'b0000000000000000;
	sram_mem[74898] = 16'b0000000000000000;
	sram_mem[74899] = 16'b0000000000000000;
	sram_mem[74900] = 16'b0000000000000000;
	sram_mem[74901] = 16'b0000000000000000;
	sram_mem[74902] = 16'b0000000000000000;
	sram_mem[74903] = 16'b0000000000000000;
	sram_mem[74904] = 16'b0000000000000000;
	sram_mem[74905] = 16'b0000000000000000;
	sram_mem[74906] = 16'b0000000000000000;
	sram_mem[74907] = 16'b0000000000000000;
	sram_mem[74908] = 16'b0000000000000000;
	sram_mem[74909] = 16'b0000000000000000;
	sram_mem[74910] = 16'b0000000000000000;
	sram_mem[74911] = 16'b0000000000000000;
	sram_mem[74912] = 16'b0000000000000000;
	sram_mem[74913] = 16'b0000000000000000;
	sram_mem[74914] = 16'b0000000000000000;
	sram_mem[74915] = 16'b0000000000000000;
	sram_mem[74916] = 16'b0000000000000000;
	sram_mem[74917] = 16'b0000000000000000;
	sram_mem[74918] = 16'b0000000000000000;
	sram_mem[74919] = 16'b0000000000000000;
	sram_mem[74920] = 16'b0000000000000000;
	sram_mem[74921] = 16'b0000000000000000;
	sram_mem[74922] = 16'b0000000000000000;
	sram_mem[74923] = 16'b0000000000000000;
	sram_mem[74924] = 16'b0000000000000000;
	sram_mem[74925] = 16'b0000000000000000;
	sram_mem[74926] = 16'b0000000000000000;
	sram_mem[74927] = 16'b0000000000000000;
	sram_mem[74928] = 16'b0000000000000000;
	sram_mem[74929] = 16'b0000000000000000;
	sram_mem[74930] = 16'b0000000000000000;
	sram_mem[74931] = 16'b0000000000000000;
	sram_mem[74932] = 16'b0000000000000000;
	sram_mem[74933] = 16'b0000000000000000;
	sram_mem[74934] = 16'b0000000000000000;
	sram_mem[74935] = 16'b0000000000000000;
	sram_mem[74936] = 16'b0000000000000000;
	sram_mem[74937] = 16'b0000000000000000;
	sram_mem[74938] = 16'b0000000000000000;
	sram_mem[74939] = 16'b0000000000000000;
	sram_mem[74940] = 16'b0000000000000000;
	sram_mem[74941] = 16'b0000000000000000;
	sram_mem[74942] = 16'b0000000000000000;
	sram_mem[74943] = 16'b0000000000000000;
	sram_mem[74944] = 16'b0000000000000000;
	sram_mem[74945] = 16'b0000000000000000;
	sram_mem[74946] = 16'b0000000000000000;
	sram_mem[74947] = 16'b0000000000000000;
	sram_mem[74948] = 16'b0000000000000000;
	sram_mem[74949] = 16'b0000000000000000;
	sram_mem[74950] = 16'b0000000000000000;
	sram_mem[74951] = 16'b0000000000000000;
	sram_mem[74952] = 16'b0000000000000000;
	sram_mem[74953] = 16'b0000000000000000;
	sram_mem[74954] = 16'b0000000000000000;
	sram_mem[74955] = 16'b0000000000000000;
	sram_mem[74956] = 16'b0000000000000000;
	sram_mem[74957] = 16'b0000000000000000;
	sram_mem[74958] = 16'b0000000000000000;
	sram_mem[74959] = 16'b0000000000000000;
	sram_mem[74960] = 16'b0000000000000000;
	sram_mem[74961] = 16'b0000000000000000;
	sram_mem[74962] = 16'b0000000000000000;
	sram_mem[74963] = 16'b0000000000000000;
	sram_mem[74964] = 16'b0000000000000000;
	sram_mem[74965] = 16'b0000000000000000;
	sram_mem[74966] = 16'b0000000000000000;
	sram_mem[74967] = 16'b0000000000000000;
	sram_mem[74968] = 16'b0000000000000000;
	sram_mem[74969] = 16'b0000000000000000;
	sram_mem[74970] = 16'b0000000000000000;
	sram_mem[74971] = 16'b0000000000000000;
	sram_mem[74972] = 16'b0000000000000000;
	sram_mem[74973] = 16'b0000000000000000;
	sram_mem[74974] = 16'b0000000000000000;
	sram_mem[74975] = 16'b0000000000000000;
	sram_mem[74976] = 16'b0000000000000000;
	sram_mem[74977] = 16'b0000000000000000;
	sram_mem[74978] = 16'b0000000000000000;
	sram_mem[74979] = 16'b0000000000000000;
	sram_mem[74980] = 16'b0000000000000000;
	sram_mem[74981] = 16'b0000000000000000;
	sram_mem[74982] = 16'b0000000000000000;
	sram_mem[74983] = 16'b0000000000000000;
	sram_mem[74984] = 16'b0000000000000000;
	sram_mem[74985] = 16'b0000000000000000;
	sram_mem[74986] = 16'b0000000000000000;
	sram_mem[74987] = 16'b0000000000000000;
	sram_mem[74988] = 16'b0000000000000000;
	sram_mem[74989] = 16'b0000000000000000;
	sram_mem[74990] = 16'b0000000000000000;
	sram_mem[74991] = 16'b0000000000000000;
	sram_mem[74992] = 16'b0000000000000000;
	sram_mem[74993] = 16'b0000000000000000;
	sram_mem[74994] = 16'b0000000000000000;
	sram_mem[74995] = 16'b0000000000000000;
	sram_mem[74996] = 16'b0000000000000000;
	sram_mem[74997] = 16'b0000000000000000;
	sram_mem[74998] = 16'b0000000000000000;
	sram_mem[74999] = 16'b0000000000000000;
	sram_mem[75000] = 16'b0000000000000000;
	sram_mem[75001] = 16'b0000000000000000;
	sram_mem[75002] = 16'b0000000000000000;
	sram_mem[75003] = 16'b0000000000000000;
	sram_mem[75004] = 16'b0000000000000000;
	sram_mem[75005] = 16'b0000000000000000;
	sram_mem[75006] = 16'b0000000000000000;
	sram_mem[75007] = 16'b0000000000000000;
	sram_mem[75008] = 16'b0000000000000000;
	sram_mem[75009] = 16'b0000000000000000;
	sram_mem[75010] = 16'b0000000000000000;
	sram_mem[75011] = 16'b0000000000000000;
	sram_mem[75012] = 16'b0000000000000000;
	sram_mem[75013] = 16'b0000000000000000;
	sram_mem[75014] = 16'b0000000000000000;
	sram_mem[75015] = 16'b0000000000000000;
	sram_mem[75016] = 16'b0000000000000000;
	sram_mem[75017] = 16'b0000000000000000;
	sram_mem[75018] = 16'b0000000000000000;
	sram_mem[75019] = 16'b0000000000000000;
	sram_mem[75020] = 16'b0000000000000000;
	sram_mem[75021] = 16'b0000000000000000;
	sram_mem[75022] = 16'b0000000000000000;
	sram_mem[75023] = 16'b0000000000000000;
	sram_mem[75024] = 16'b0000000000000000;
	sram_mem[75025] = 16'b0000000000000000;
	sram_mem[75026] = 16'b0000000000000000;
	sram_mem[75027] = 16'b0000000000000000;
	sram_mem[75028] = 16'b0000000000000000;
	sram_mem[75029] = 16'b0000000000000000;
	sram_mem[75030] = 16'b0000000000000000;
	sram_mem[75031] = 16'b0000000000000000;
	sram_mem[75032] = 16'b0000000000000000;
	sram_mem[75033] = 16'b0000000000000000;
	sram_mem[75034] = 16'b0000000000000000;
	sram_mem[75035] = 16'b0000000000000000;
	sram_mem[75036] = 16'b0000000000000000;
	sram_mem[75037] = 16'b0000000000000000;
	sram_mem[75038] = 16'b0000000000000000;
	sram_mem[75039] = 16'b0000000000000000;
	sram_mem[75040] = 16'b0000000000000000;
	sram_mem[75041] = 16'b0000000000000000;
	sram_mem[75042] = 16'b0000000000000000;
	sram_mem[75043] = 16'b0000000000000000;
	sram_mem[75044] = 16'b0000000000000000;
	sram_mem[75045] = 16'b0000000000000000;
	sram_mem[75046] = 16'b0000000000000000;
	sram_mem[75047] = 16'b0000000000000000;
	sram_mem[75048] = 16'b0000000000000000;
	sram_mem[75049] = 16'b0000000000000000;
	sram_mem[75050] = 16'b0000000000000000;
	sram_mem[75051] = 16'b0000000000000000;
	sram_mem[75052] = 16'b0000000000000000;
	sram_mem[75053] = 16'b0000000000000000;
	sram_mem[75054] = 16'b0000000000000000;
	sram_mem[75055] = 16'b0000000000000000;
	sram_mem[75056] = 16'b0000000000000000;
	sram_mem[75057] = 16'b0000000000000000;
	sram_mem[75058] = 16'b0000000000000000;
	sram_mem[75059] = 16'b0000000000000000;
	sram_mem[75060] = 16'b0000000000000000;
	sram_mem[75061] = 16'b0000000000000000;
	sram_mem[75062] = 16'b0000000000000000;
	sram_mem[75063] = 16'b0000000000000000;
	sram_mem[75064] = 16'b0000000000000000;
	sram_mem[75065] = 16'b0000000000000000;
	sram_mem[75066] = 16'b0000000000000000;
	sram_mem[75067] = 16'b0000000000000000;
	sram_mem[75068] = 16'b0000000000000000;
	sram_mem[75069] = 16'b0000000000000000;
	sram_mem[75070] = 16'b0000000000000000;
	sram_mem[75071] = 16'b0000000000000000;
	sram_mem[75072] = 16'b0000000000000000;
	sram_mem[75073] = 16'b0000000000000000;
	sram_mem[75074] = 16'b0000000000000000;
	sram_mem[75075] = 16'b0000000000000000;
	sram_mem[75076] = 16'b0000000000000000;
	sram_mem[75077] = 16'b0000000000000000;
	sram_mem[75078] = 16'b0000000000000000;
	sram_mem[75079] = 16'b0000000000000000;
	sram_mem[75080] = 16'b0000000000000000;
	sram_mem[75081] = 16'b0000000000000000;
	sram_mem[75082] = 16'b0000000000000000;
	sram_mem[75083] = 16'b0000000000000000;
	sram_mem[75084] = 16'b0000000000000000;
	sram_mem[75085] = 16'b0000000000000000;
	sram_mem[75086] = 16'b0000000000000000;
	sram_mem[75087] = 16'b0000000000000000;
	sram_mem[75088] = 16'b0000000000000000;
	sram_mem[75089] = 16'b0000000000000000;
	sram_mem[75090] = 16'b0000000000000000;
	sram_mem[75091] = 16'b0000000000000000;
	sram_mem[75092] = 16'b0000000000000000;
	sram_mem[75093] = 16'b0000000000000000;
	sram_mem[75094] = 16'b0000000000000000;
	sram_mem[75095] = 16'b0000000000000000;
	sram_mem[75096] = 16'b0000000000000000;
	sram_mem[75097] = 16'b0000000000000000;
	sram_mem[75098] = 16'b0000000000000000;
	sram_mem[75099] = 16'b0000000000000000;
	sram_mem[75100] = 16'b0000000000000000;
	sram_mem[75101] = 16'b0000000000000000;
	sram_mem[75102] = 16'b0000000000000000;
	sram_mem[75103] = 16'b0000000000000000;
	sram_mem[75104] = 16'b0000000000000000;
	sram_mem[75105] = 16'b0000000000000000;
	sram_mem[75106] = 16'b0000000000000000;
	sram_mem[75107] = 16'b0000000000000000;
	sram_mem[75108] = 16'b0000000000000000;
	sram_mem[75109] = 16'b0000000000000000;
	sram_mem[75110] = 16'b0000000000000000;
	sram_mem[75111] = 16'b0000000000000000;
	sram_mem[75112] = 16'b0000000000000000;
	sram_mem[75113] = 16'b0000000000000000;
	sram_mem[75114] = 16'b0000000000000000;
	sram_mem[75115] = 16'b0000000000000000;
	sram_mem[75116] = 16'b0000000000000000;
	sram_mem[75117] = 16'b0000000000000000;
	sram_mem[75118] = 16'b0000000000000000;
	sram_mem[75119] = 16'b0000000000000000;
	sram_mem[75120] = 16'b0000000000000000;
	sram_mem[75121] = 16'b0000000000000000;
	sram_mem[75122] = 16'b0000000000000000;
	sram_mem[75123] = 16'b0000000000000000;
	sram_mem[75124] = 16'b0000000000000000;
	sram_mem[75125] = 16'b0000000000000000;
	sram_mem[75126] = 16'b0000000000000000;
	sram_mem[75127] = 16'b0000000000000000;
	sram_mem[75128] = 16'b0000000000000000;
	sram_mem[75129] = 16'b0000000000000000;
	sram_mem[75130] = 16'b0000000000000000;
	sram_mem[75131] = 16'b0000000000000000;
	sram_mem[75132] = 16'b0000000000000000;
	sram_mem[75133] = 16'b0000000000000000;
	sram_mem[75134] = 16'b0000000000000000;
	sram_mem[75135] = 16'b0000000000000000;
	sram_mem[75136] = 16'b0000000000000000;
	sram_mem[75137] = 16'b0000000000000000;
	sram_mem[75138] = 16'b0000000000000000;
	sram_mem[75139] = 16'b0000000000000000;
	sram_mem[75140] = 16'b0000000000000000;
	sram_mem[75141] = 16'b0000000000000000;
	sram_mem[75142] = 16'b0000000000000000;
	sram_mem[75143] = 16'b0000000000000000;
	sram_mem[75144] = 16'b0000000000000000;
	sram_mem[75145] = 16'b0000000000000000;
	sram_mem[75146] = 16'b0000000000000000;
	sram_mem[75147] = 16'b0000000000000000;
	sram_mem[75148] = 16'b0000000000000000;
	sram_mem[75149] = 16'b0000000000000000;
	sram_mem[75150] = 16'b0000000000000000;
	sram_mem[75151] = 16'b0000000000000000;
	sram_mem[75152] = 16'b0000000000000000;
	sram_mem[75153] = 16'b0000000000000000;
	sram_mem[75154] = 16'b0000000000000000;
	sram_mem[75155] = 16'b0000000000000000;
	sram_mem[75156] = 16'b0000000000000000;
	sram_mem[75157] = 16'b0000000000000000;
	sram_mem[75158] = 16'b0000000000000000;
	sram_mem[75159] = 16'b0000000000000000;
	sram_mem[75160] = 16'b0000000000000000;
	sram_mem[75161] = 16'b0000000000000000;
	sram_mem[75162] = 16'b0000000000000000;
	sram_mem[75163] = 16'b0000000000000000;
	sram_mem[75164] = 16'b0000000000000000;
	sram_mem[75165] = 16'b0000000000000000;
	sram_mem[75166] = 16'b0000000000000000;
	sram_mem[75167] = 16'b0000000000000000;
	sram_mem[75168] = 16'b0000000000000000;
	sram_mem[75169] = 16'b0000000000000000;
	sram_mem[75170] = 16'b0000000000000000;
	sram_mem[75171] = 16'b0000000000000000;
	sram_mem[75172] = 16'b0000000000000000;
	sram_mem[75173] = 16'b0000000000000000;
	sram_mem[75174] = 16'b0000000000000000;
	sram_mem[75175] = 16'b0000000000000000;
	sram_mem[75176] = 16'b0000000000000000;
	sram_mem[75177] = 16'b0000000000000000;
	sram_mem[75178] = 16'b0000000000000000;
	sram_mem[75179] = 16'b0000000000000000;
	sram_mem[75180] = 16'b0000000000000000;
	sram_mem[75181] = 16'b0000000000000000;
	sram_mem[75182] = 16'b0000000000000000;
	sram_mem[75183] = 16'b0000000000000000;
	sram_mem[75184] = 16'b0000000000000000;
	sram_mem[75185] = 16'b0000000000000000;
	sram_mem[75186] = 16'b0000000000000000;
	sram_mem[75187] = 16'b0000000000000000;
	sram_mem[75188] = 16'b0000000000000000;
	sram_mem[75189] = 16'b0000000000000000;
	sram_mem[75190] = 16'b0000000000000000;
	sram_mem[75191] = 16'b0000000000000000;
	sram_mem[75192] = 16'b0000000000000000;
	sram_mem[75193] = 16'b0000000000000000;
	sram_mem[75194] = 16'b0000000000000000;
	sram_mem[75195] = 16'b0000000000000000;
	sram_mem[75196] = 16'b0000000000000000;
	sram_mem[75197] = 16'b0000000000000000;
	sram_mem[75198] = 16'b0000000000000000;
	sram_mem[75199] = 16'b0000000000000000;
	sram_mem[75200] = 16'b0000000000000000;
	sram_mem[75201] = 16'b0000000000000000;
	sram_mem[75202] = 16'b0000000000000000;
	sram_mem[75203] = 16'b0000000000000000;
	sram_mem[75204] = 16'b0000000000000000;
	sram_mem[75205] = 16'b0000000000000000;
	sram_mem[75206] = 16'b0000000000000000;
	sram_mem[75207] = 16'b0000000000000000;
	sram_mem[75208] = 16'b0000000000000000;
	sram_mem[75209] = 16'b0000000000000000;
	sram_mem[75210] = 16'b0000000000000000;
	sram_mem[75211] = 16'b0000000000000000;
	sram_mem[75212] = 16'b0000000000000000;
	sram_mem[75213] = 16'b0000000000000000;
	sram_mem[75214] = 16'b0000000000000000;
	sram_mem[75215] = 16'b0000000000000000;
	sram_mem[75216] = 16'b0000000000000000;
	sram_mem[75217] = 16'b0000000000000000;
	sram_mem[75218] = 16'b0000000000000000;
	sram_mem[75219] = 16'b0000000000000000;
	sram_mem[75220] = 16'b0000000000000000;
	sram_mem[75221] = 16'b0000000000000000;
	sram_mem[75222] = 16'b0000000000000000;
	sram_mem[75223] = 16'b0000000000000000;
	sram_mem[75224] = 16'b0000000000000000;
	sram_mem[75225] = 16'b0000000000000000;
	sram_mem[75226] = 16'b0000000000000000;
	sram_mem[75227] = 16'b0000000000000000;
	sram_mem[75228] = 16'b0000000000000000;
	sram_mem[75229] = 16'b0000000000000000;
	sram_mem[75230] = 16'b0000000000000000;
	sram_mem[75231] = 16'b0000000000000000;
	sram_mem[75232] = 16'b0000000000000000;
	sram_mem[75233] = 16'b0000000000000000;
	sram_mem[75234] = 16'b0000000000000000;
	sram_mem[75235] = 16'b0000000000000000;
	sram_mem[75236] = 16'b0000000000000000;
	sram_mem[75237] = 16'b0000000000000000;
	sram_mem[75238] = 16'b0000000000000000;
	sram_mem[75239] = 16'b0000000000000000;
	sram_mem[75240] = 16'b0000000000000000;
	sram_mem[75241] = 16'b0000000000000000;
	sram_mem[75242] = 16'b0000000000000000;
	sram_mem[75243] = 16'b0000000000000000;
	sram_mem[75244] = 16'b0000000000000000;
	sram_mem[75245] = 16'b0000000000000000;
	sram_mem[75246] = 16'b0000000000000000;
	sram_mem[75247] = 16'b0000000000000000;
	sram_mem[75248] = 16'b0000000000000000;
	sram_mem[75249] = 16'b0000000000000000;
	sram_mem[75250] = 16'b0000000000000000;
	sram_mem[75251] = 16'b0000000000000000;
	sram_mem[75252] = 16'b0000000000000000;
	sram_mem[75253] = 16'b0000000000000000;
	sram_mem[75254] = 16'b0000000000000000;
	sram_mem[75255] = 16'b0000000000000000;
	sram_mem[75256] = 16'b0000000000000000;
	sram_mem[75257] = 16'b0000000000000000;
	sram_mem[75258] = 16'b0000000000000000;
	sram_mem[75259] = 16'b0000000000000000;
	sram_mem[75260] = 16'b0000000000000000;
	sram_mem[75261] = 16'b0000000000000000;
	sram_mem[75262] = 16'b0000000000000000;
	sram_mem[75263] = 16'b0000000000000000;
	sram_mem[75264] = 16'b0000000000000000;
	sram_mem[75265] = 16'b0000000000000000;
	sram_mem[75266] = 16'b0000000000000000;
	sram_mem[75267] = 16'b0000000000000000;
	sram_mem[75268] = 16'b0000000000000000;
	sram_mem[75269] = 16'b0000000000000000;
	sram_mem[75270] = 16'b0000000000000000;
	sram_mem[75271] = 16'b0000000000000000;
	sram_mem[75272] = 16'b0000000000000000;
	sram_mem[75273] = 16'b0000000000000000;
	sram_mem[75274] = 16'b0000000000000000;
	sram_mem[75275] = 16'b0000000000000000;
	sram_mem[75276] = 16'b0000000000000000;
	sram_mem[75277] = 16'b0000000000000000;
	sram_mem[75278] = 16'b0000000000000000;
	sram_mem[75279] = 16'b0000000000000000;
	sram_mem[75280] = 16'b0000000000000000;
	sram_mem[75281] = 16'b0000000000000000;
	sram_mem[75282] = 16'b0000000000000000;
	sram_mem[75283] = 16'b0000000000000000;
	sram_mem[75284] = 16'b0000000000000000;
	sram_mem[75285] = 16'b0000000000000000;
	sram_mem[75286] = 16'b0000000000000000;
	sram_mem[75287] = 16'b0000000000000000;
	sram_mem[75288] = 16'b0000000000000000;
	sram_mem[75289] = 16'b0000000000000000;
	sram_mem[75290] = 16'b0000000000000000;
	sram_mem[75291] = 16'b0000000000000000;
	sram_mem[75292] = 16'b0000000000000000;
	sram_mem[75293] = 16'b0000000000000000;
	sram_mem[75294] = 16'b0000000000000000;
	sram_mem[75295] = 16'b0000000000000000;
	sram_mem[75296] = 16'b0000000000000000;
	sram_mem[75297] = 16'b0000000000000000;
	sram_mem[75298] = 16'b0000000000000000;
	sram_mem[75299] = 16'b0000000000000000;
	sram_mem[75300] = 16'b0000000000000000;
	sram_mem[75301] = 16'b0000000000000000;
	sram_mem[75302] = 16'b0000000000000000;
	sram_mem[75303] = 16'b0000000000000000;
	sram_mem[75304] = 16'b0000000000000000;
	sram_mem[75305] = 16'b0000000000000000;
	sram_mem[75306] = 16'b0000000000000000;
	sram_mem[75307] = 16'b0000000000000000;
	sram_mem[75308] = 16'b0000000000000000;
	sram_mem[75309] = 16'b0000000000000000;
	sram_mem[75310] = 16'b0000000000000000;
	sram_mem[75311] = 16'b0000000000000000;
	sram_mem[75312] = 16'b0000000000000000;
	sram_mem[75313] = 16'b0000000000000000;
	sram_mem[75314] = 16'b0000000000000000;
	sram_mem[75315] = 16'b0000000000000000;
	sram_mem[75316] = 16'b0000000000000000;
	sram_mem[75317] = 16'b0000000000000000;
	sram_mem[75318] = 16'b0000000000000000;
	sram_mem[75319] = 16'b0000000000000000;
	sram_mem[75320] = 16'b0000000000000000;
	sram_mem[75321] = 16'b0000000000000000;
	sram_mem[75322] = 16'b0000000000000000;
	sram_mem[75323] = 16'b0000000000000000;
	sram_mem[75324] = 16'b0000000000000000;
	sram_mem[75325] = 16'b0000000000000000;
	sram_mem[75326] = 16'b0000000000000000;
	sram_mem[75327] = 16'b0000000000000000;
	sram_mem[75328] = 16'b0000000000000000;
	sram_mem[75329] = 16'b0000000000000000;
	sram_mem[75330] = 16'b0000000000000000;
	sram_mem[75331] = 16'b0000000000000000;
	sram_mem[75332] = 16'b0000000000000000;
	sram_mem[75333] = 16'b0000000000000000;
	sram_mem[75334] = 16'b0000000000000000;
	sram_mem[75335] = 16'b0000000000000000;
	sram_mem[75336] = 16'b0000000000000000;
	sram_mem[75337] = 16'b0000000000000000;
	sram_mem[75338] = 16'b0000000000000000;
	sram_mem[75339] = 16'b0000000000000000;
	sram_mem[75340] = 16'b0000000000000000;
	sram_mem[75341] = 16'b0000000000000000;
	sram_mem[75342] = 16'b0000000000000000;
	sram_mem[75343] = 16'b0000000000000000;
	sram_mem[75344] = 16'b0000000000000000;
	sram_mem[75345] = 16'b0000000000000000;
	sram_mem[75346] = 16'b0000000000000000;
	sram_mem[75347] = 16'b0000000000000000;
	sram_mem[75348] = 16'b0000000000000000;
	sram_mem[75349] = 16'b0000000000000000;
	sram_mem[75350] = 16'b0000000000000000;
	sram_mem[75351] = 16'b0000000000000000;
	sram_mem[75352] = 16'b0000000000000000;
	sram_mem[75353] = 16'b0000000000000000;
	sram_mem[75354] = 16'b0000000000000000;
	sram_mem[75355] = 16'b0000000000000000;
	sram_mem[75356] = 16'b0000000000000000;
	sram_mem[75357] = 16'b0000000000000000;
	sram_mem[75358] = 16'b0000000000000000;
	sram_mem[75359] = 16'b0000000000000000;
	sram_mem[75360] = 16'b0000000000000000;
	sram_mem[75361] = 16'b0000000000000000;
	sram_mem[75362] = 16'b0000000000000000;
	sram_mem[75363] = 16'b0000000000000000;
	sram_mem[75364] = 16'b0000000000000000;
	sram_mem[75365] = 16'b0000000000000000;
	sram_mem[75366] = 16'b0000000000000000;
	sram_mem[75367] = 16'b0000000000000000;
	sram_mem[75368] = 16'b0000000000000000;
	sram_mem[75369] = 16'b0000000000000000;
	sram_mem[75370] = 16'b0000000000000000;
	sram_mem[75371] = 16'b0000000000000000;
	sram_mem[75372] = 16'b0000000000000000;
	sram_mem[75373] = 16'b0000000000000000;
	sram_mem[75374] = 16'b0000000000000000;
	sram_mem[75375] = 16'b0000000000000000;
	sram_mem[75376] = 16'b0000000000000000;
	sram_mem[75377] = 16'b0000000000000000;
	sram_mem[75378] = 16'b0000000000000000;
	sram_mem[75379] = 16'b0000000000000000;
	sram_mem[75380] = 16'b0000000000000000;
	sram_mem[75381] = 16'b0000000000000000;
	sram_mem[75382] = 16'b0000000000000000;
	sram_mem[75383] = 16'b0000000000000000;
	sram_mem[75384] = 16'b0000000000000000;
	sram_mem[75385] = 16'b0000000000000000;
	sram_mem[75386] = 16'b0000000000000000;
	sram_mem[75387] = 16'b0000000000000000;
	sram_mem[75388] = 16'b0000000000000000;
	sram_mem[75389] = 16'b0000000000000000;
	sram_mem[75390] = 16'b0000000000000000;
	sram_mem[75391] = 16'b0000000000000000;
	sram_mem[75392] = 16'b0000000000000000;
	sram_mem[75393] = 16'b0000000000000000;
	sram_mem[75394] = 16'b0000000000000000;
	sram_mem[75395] = 16'b0000000000000000;
	sram_mem[75396] = 16'b0000000000000000;
	sram_mem[75397] = 16'b0000000000000000;
	sram_mem[75398] = 16'b0000000000000000;
	sram_mem[75399] = 16'b0000000000000000;
	sram_mem[75400] = 16'b0000000000000000;
	sram_mem[75401] = 16'b0000000000000000;
	sram_mem[75402] = 16'b0000000000000000;
	sram_mem[75403] = 16'b0000000000000000;
	sram_mem[75404] = 16'b0000000000000000;
	sram_mem[75405] = 16'b0000000000000000;
	sram_mem[75406] = 16'b0000000000000000;
	sram_mem[75407] = 16'b0000000000000000;
	sram_mem[75408] = 16'b0000000000000000;
	sram_mem[75409] = 16'b0000000000000000;
	sram_mem[75410] = 16'b0000000000000000;
	sram_mem[75411] = 16'b0000000000000000;
	sram_mem[75412] = 16'b0000000000000000;
	sram_mem[75413] = 16'b0000000000000000;
	sram_mem[75414] = 16'b0000000000000000;
	sram_mem[75415] = 16'b0000000000000000;
	sram_mem[75416] = 16'b0000000000000000;
	sram_mem[75417] = 16'b0000000000000000;
	sram_mem[75418] = 16'b0000000000000000;
	sram_mem[75419] = 16'b0000000000000000;
	sram_mem[75420] = 16'b0000000000000000;
	sram_mem[75421] = 16'b0000000000000000;
	sram_mem[75422] = 16'b0000000000000000;
	sram_mem[75423] = 16'b0000000000000000;
	sram_mem[75424] = 16'b0000000000000000;
	sram_mem[75425] = 16'b0000000000000000;
	sram_mem[75426] = 16'b0000000000000000;
	sram_mem[75427] = 16'b0000000000000000;
	sram_mem[75428] = 16'b0000000000000000;
	sram_mem[75429] = 16'b0000000000000000;
	sram_mem[75430] = 16'b0000000000000000;
	sram_mem[75431] = 16'b0000000000000000;
	sram_mem[75432] = 16'b0000000000000000;
	sram_mem[75433] = 16'b0000000000000000;
	sram_mem[75434] = 16'b0000000000000000;
	sram_mem[75435] = 16'b0000000000000000;
	sram_mem[75436] = 16'b0000000000000000;
	sram_mem[75437] = 16'b0000000000000000;
	sram_mem[75438] = 16'b0000000000000000;
	sram_mem[75439] = 16'b0000000000000000;
	sram_mem[75440] = 16'b0000000000000000;
	sram_mem[75441] = 16'b0000000000000000;
	sram_mem[75442] = 16'b0000000000000000;
	sram_mem[75443] = 16'b0000000000000000;
	sram_mem[75444] = 16'b0000000000000000;
	sram_mem[75445] = 16'b0000000000000000;
	sram_mem[75446] = 16'b0000000000000000;
	sram_mem[75447] = 16'b0000000000000000;
	sram_mem[75448] = 16'b0000000000000000;
	sram_mem[75449] = 16'b0000000000000000;
	sram_mem[75450] = 16'b0000000000000000;
	sram_mem[75451] = 16'b0000000000000000;
	sram_mem[75452] = 16'b0000000000000000;
	sram_mem[75453] = 16'b0000000000000000;
	sram_mem[75454] = 16'b0000000000000000;
	sram_mem[75455] = 16'b0000000000000000;
	sram_mem[75456] = 16'b0000000000000000;
	sram_mem[75457] = 16'b0000000000000000;
	sram_mem[75458] = 16'b0000000000000000;
	sram_mem[75459] = 16'b0000000000000000;
	sram_mem[75460] = 16'b0000000000000000;
	sram_mem[75461] = 16'b0000000000000000;
	sram_mem[75462] = 16'b0000000000000000;
	sram_mem[75463] = 16'b0000000000000000;
	sram_mem[75464] = 16'b0000000000000000;
	sram_mem[75465] = 16'b0000000000000000;
	sram_mem[75466] = 16'b0000000000000000;
	sram_mem[75467] = 16'b0000000000000000;
	sram_mem[75468] = 16'b0000000000000000;
	sram_mem[75469] = 16'b0000000000000000;
	sram_mem[75470] = 16'b0000000000000000;
	sram_mem[75471] = 16'b0000000000000000;
	sram_mem[75472] = 16'b0000000000000000;
	sram_mem[75473] = 16'b0000000000000000;
	sram_mem[75474] = 16'b0000000000000000;
	sram_mem[75475] = 16'b0000000000000000;
	sram_mem[75476] = 16'b0000000000000000;
	sram_mem[75477] = 16'b0000000000000000;
	sram_mem[75478] = 16'b0000000000000000;
	sram_mem[75479] = 16'b0000000000000000;
	sram_mem[75480] = 16'b0000000000000000;
	sram_mem[75481] = 16'b0000000000000000;
	sram_mem[75482] = 16'b0000000000000000;
	sram_mem[75483] = 16'b0000000000000000;
	sram_mem[75484] = 16'b0000000000000000;
	sram_mem[75485] = 16'b0000000000000000;
	sram_mem[75486] = 16'b0000000000000000;
	sram_mem[75487] = 16'b0000000000000000;
	sram_mem[75488] = 16'b0000000000000000;
	sram_mem[75489] = 16'b0000000000000000;
	sram_mem[75490] = 16'b0000000000000000;
	sram_mem[75491] = 16'b0000000000000000;
	sram_mem[75492] = 16'b0000000000000000;
	sram_mem[75493] = 16'b0000000000000000;
	sram_mem[75494] = 16'b0000000000000000;
	sram_mem[75495] = 16'b0000000000000000;
	sram_mem[75496] = 16'b0000000000000000;
	sram_mem[75497] = 16'b0000000000000000;
	sram_mem[75498] = 16'b0000000000000000;
	sram_mem[75499] = 16'b0000000000000000;
	sram_mem[75500] = 16'b0000000000000000;
	sram_mem[75501] = 16'b0000000000000000;
	sram_mem[75502] = 16'b0000000000000000;
	sram_mem[75503] = 16'b0000000000000000;
	sram_mem[75504] = 16'b0000000000000000;
	sram_mem[75505] = 16'b0000000000000000;
	sram_mem[75506] = 16'b0000000000000000;
	sram_mem[75507] = 16'b0000000000000000;
	sram_mem[75508] = 16'b0000000000000000;
	sram_mem[75509] = 16'b0000000000000000;
	sram_mem[75510] = 16'b0000000000000000;
	sram_mem[75511] = 16'b0000000000000000;
	sram_mem[75512] = 16'b0000000000000000;
	sram_mem[75513] = 16'b0000000000000000;
	sram_mem[75514] = 16'b0000000000000000;
	sram_mem[75515] = 16'b0000000000000000;
	sram_mem[75516] = 16'b0000000000000000;
	sram_mem[75517] = 16'b0000000000000000;
	sram_mem[75518] = 16'b0000000000000000;
	sram_mem[75519] = 16'b0000000000000000;
	sram_mem[75520] = 16'b0000000000000000;
	sram_mem[75521] = 16'b0000000000000000;
	sram_mem[75522] = 16'b0000000000000000;
	sram_mem[75523] = 16'b0000000000000000;
	sram_mem[75524] = 16'b0000000000000000;
	sram_mem[75525] = 16'b0000000000000000;
	sram_mem[75526] = 16'b0000000000000000;
	sram_mem[75527] = 16'b0000000000000000;
	sram_mem[75528] = 16'b0000000000000000;
	sram_mem[75529] = 16'b0000000000000000;
	sram_mem[75530] = 16'b0000000000000000;
	sram_mem[75531] = 16'b0000000000000000;
	sram_mem[75532] = 16'b0000000000000000;
	sram_mem[75533] = 16'b0000000000000000;
	sram_mem[75534] = 16'b0000000000000000;
	sram_mem[75535] = 16'b0000000000000000;
	sram_mem[75536] = 16'b0000000000000000;
	sram_mem[75537] = 16'b0000000000000000;
	sram_mem[75538] = 16'b0000000000000000;
	sram_mem[75539] = 16'b0000000000000000;
	sram_mem[75540] = 16'b0000000000000000;
	sram_mem[75541] = 16'b0000000000000000;
	sram_mem[75542] = 16'b0000000000000000;
	sram_mem[75543] = 16'b0000000000000000;
	sram_mem[75544] = 16'b0000000000000000;
	sram_mem[75545] = 16'b0000000000000000;
	sram_mem[75546] = 16'b0000000000000000;
	sram_mem[75547] = 16'b0000000000000000;
	sram_mem[75548] = 16'b0000000000000000;
	sram_mem[75549] = 16'b0000000000000000;
	sram_mem[75550] = 16'b0000000000000000;
	sram_mem[75551] = 16'b0000000000000000;
	sram_mem[75552] = 16'b0000000000000000;
	sram_mem[75553] = 16'b0000000000000000;
	sram_mem[75554] = 16'b0000000000000000;
	sram_mem[75555] = 16'b0000000000000000;
	sram_mem[75556] = 16'b0000000000000000;
	sram_mem[75557] = 16'b0000000000000000;
	sram_mem[75558] = 16'b0000000000000000;
	sram_mem[75559] = 16'b0000000000000000;
	sram_mem[75560] = 16'b0000000000000000;
	sram_mem[75561] = 16'b0000000000000000;
	sram_mem[75562] = 16'b0000000000000000;
	sram_mem[75563] = 16'b0000000000000000;
	sram_mem[75564] = 16'b0000000000000000;
	sram_mem[75565] = 16'b0000000000000000;
	sram_mem[75566] = 16'b0000000000000000;
	sram_mem[75567] = 16'b0000000000000000;
	sram_mem[75568] = 16'b0000000000000000;
	sram_mem[75569] = 16'b0000000000000000;
	sram_mem[75570] = 16'b0000000000000000;
	sram_mem[75571] = 16'b0000000000000000;
	sram_mem[75572] = 16'b0000000000000000;
	sram_mem[75573] = 16'b0000000000000000;
	sram_mem[75574] = 16'b0000000000000000;
	sram_mem[75575] = 16'b0000000000000000;
	sram_mem[75576] = 16'b0000000000000000;
	sram_mem[75577] = 16'b0000000000000000;
	sram_mem[75578] = 16'b0000000000000000;
	sram_mem[75579] = 16'b0000000000000000;
	sram_mem[75580] = 16'b0000000000000000;
	sram_mem[75581] = 16'b0000000000000000;
	sram_mem[75582] = 16'b0000000000000000;
	sram_mem[75583] = 16'b0000000000000000;
	sram_mem[75584] = 16'b0000000000000000;
	sram_mem[75585] = 16'b0000000000000000;
	sram_mem[75586] = 16'b0000000000000000;
	sram_mem[75587] = 16'b0000000000000000;
	sram_mem[75588] = 16'b0000000000000000;
	sram_mem[75589] = 16'b0000000000000000;
	sram_mem[75590] = 16'b0000000000000000;
	sram_mem[75591] = 16'b0000000000000000;
	sram_mem[75592] = 16'b0000000000000000;
	sram_mem[75593] = 16'b0000000000000000;
	sram_mem[75594] = 16'b0000000000000000;
	sram_mem[75595] = 16'b0000000000000000;
	sram_mem[75596] = 16'b0000000000000000;
	sram_mem[75597] = 16'b0000000000000000;
	sram_mem[75598] = 16'b0000000000000000;
	sram_mem[75599] = 16'b0000000000000000;
	sram_mem[75600] = 16'b0000000000000000;
	sram_mem[75601] = 16'b0000000000000000;
	sram_mem[75602] = 16'b0000000000000000;
	sram_mem[75603] = 16'b0000000000000000;
	sram_mem[75604] = 16'b0000000000000000;
	sram_mem[75605] = 16'b0000000000000000;
	sram_mem[75606] = 16'b0000000000000000;
	sram_mem[75607] = 16'b0000000000000000;
	sram_mem[75608] = 16'b0000000000000000;
	sram_mem[75609] = 16'b0000000000000000;
	sram_mem[75610] = 16'b0000000000000000;
	sram_mem[75611] = 16'b0000000000000000;
	sram_mem[75612] = 16'b0000000000000000;
	sram_mem[75613] = 16'b0000000000000000;
	sram_mem[75614] = 16'b0000000000000000;
	sram_mem[75615] = 16'b0000000000000000;
	sram_mem[75616] = 16'b0000000000000000;
	sram_mem[75617] = 16'b0000000000000000;
	sram_mem[75618] = 16'b0000000000000000;
	sram_mem[75619] = 16'b0000000000000000;
	sram_mem[75620] = 16'b0000000000000000;
	sram_mem[75621] = 16'b0000000000000000;
	sram_mem[75622] = 16'b0000000000000000;
	sram_mem[75623] = 16'b0000000000000000;
	sram_mem[75624] = 16'b0000000000000000;
	sram_mem[75625] = 16'b0000000000000000;
	sram_mem[75626] = 16'b0000000000000000;
	sram_mem[75627] = 16'b0000000000000000;
	sram_mem[75628] = 16'b0000000000000000;
	sram_mem[75629] = 16'b0000000000000000;
	sram_mem[75630] = 16'b0000000000000000;
	sram_mem[75631] = 16'b0000000000000000;
	sram_mem[75632] = 16'b0000000000000000;
	sram_mem[75633] = 16'b0000000000000000;
	sram_mem[75634] = 16'b0000000000000000;
	sram_mem[75635] = 16'b0000000000000000;
	sram_mem[75636] = 16'b0000000000000000;
	sram_mem[75637] = 16'b0000000000000000;
	sram_mem[75638] = 16'b0000000000000000;
	sram_mem[75639] = 16'b0000000000000000;
	sram_mem[75640] = 16'b0000000000000000;
	sram_mem[75641] = 16'b0000000000000000;
	sram_mem[75642] = 16'b0000000000000000;
	sram_mem[75643] = 16'b0000000000000000;
	sram_mem[75644] = 16'b0000000000000000;
	sram_mem[75645] = 16'b0000000000000000;
	sram_mem[75646] = 16'b0000000000000000;
	sram_mem[75647] = 16'b0000000000000000;
	sram_mem[75648] = 16'b0000000000000000;
	sram_mem[75649] = 16'b0000000000000000;
	sram_mem[75650] = 16'b0000000000000000;
	sram_mem[75651] = 16'b0000000000000000;
	sram_mem[75652] = 16'b0000000000000000;
	sram_mem[75653] = 16'b0000000000000000;
	sram_mem[75654] = 16'b0000000000000000;
	sram_mem[75655] = 16'b0000000000000000;
	sram_mem[75656] = 16'b0000000000000000;
	sram_mem[75657] = 16'b0000000000000000;
	sram_mem[75658] = 16'b0000000000000000;
	sram_mem[75659] = 16'b0000000000000000;
	sram_mem[75660] = 16'b0000000000000000;
	sram_mem[75661] = 16'b0000000000000000;
	sram_mem[75662] = 16'b0000000000000000;
	sram_mem[75663] = 16'b0000000000000000;
	sram_mem[75664] = 16'b0000000000000000;
	sram_mem[75665] = 16'b0000000000000000;
	sram_mem[75666] = 16'b0000000000000000;
	sram_mem[75667] = 16'b0000000000000000;
	sram_mem[75668] = 16'b0000000000000000;
	sram_mem[75669] = 16'b0000000000000000;
	sram_mem[75670] = 16'b0000000000000000;
	sram_mem[75671] = 16'b0000000000000000;
	sram_mem[75672] = 16'b0000000000000000;
	sram_mem[75673] = 16'b0000000000000000;
	sram_mem[75674] = 16'b0000000000000000;
	sram_mem[75675] = 16'b0000000000000000;
	sram_mem[75676] = 16'b0000000000000000;
	sram_mem[75677] = 16'b0000000000000000;
	sram_mem[75678] = 16'b0000000000000000;
	sram_mem[75679] = 16'b0000000000000000;
	sram_mem[75680] = 16'b0000000000000000;
	sram_mem[75681] = 16'b0000000000000000;
	sram_mem[75682] = 16'b0000000000000000;
	sram_mem[75683] = 16'b0000000000000000;
	sram_mem[75684] = 16'b0000000000000000;
	sram_mem[75685] = 16'b0000000000000000;
	sram_mem[75686] = 16'b0000000000000000;
	sram_mem[75687] = 16'b0000000000000000;
	sram_mem[75688] = 16'b0000000000000000;
	sram_mem[75689] = 16'b0000000000000000;
	sram_mem[75690] = 16'b0000000000000000;
	sram_mem[75691] = 16'b0000000000000000;
	sram_mem[75692] = 16'b0000000000000000;
	sram_mem[75693] = 16'b0000000000000000;
	sram_mem[75694] = 16'b0000000000000000;
	sram_mem[75695] = 16'b0000000000000000;
	sram_mem[75696] = 16'b0000000000000000;
	sram_mem[75697] = 16'b0000000000000000;
	sram_mem[75698] = 16'b0000000000000000;
	sram_mem[75699] = 16'b0000000000000000;
	sram_mem[75700] = 16'b0000000000000000;
	sram_mem[75701] = 16'b0000000000000000;
	sram_mem[75702] = 16'b0000000000000000;
	sram_mem[75703] = 16'b0000000000000000;
	sram_mem[75704] = 16'b0000000000000000;
	sram_mem[75705] = 16'b0000000000000000;
	sram_mem[75706] = 16'b0000000000000000;
	sram_mem[75707] = 16'b0000000000000000;
	sram_mem[75708] = 16'b0000000000000000;
	sram_mem[75709] = 16'b0000000000000000;
	sram_mem[75710] = 16'b0000000000000000;
	sram_mem[75711] = 16'b0000000000000000;
	sram_mem[75712] = 16'b0000000000000000;
	sram_mem[75713] = 16'b0000000000000000;
	sram_mem[75714] = 16'b0000000000000000;
	sram_mem[75715] = 16'b0000000000000000;
	sram_mem[75716] = 16'b0000000000000000;
	sram_mem[75717] = 16'b0000000000000000;
	sram_mem[75718] = 16'b0000000000000000;
	sram_mem[75719] = 16'b0000000000000000;
	sram_mem[75720] = 16'b0000000000000000;
	sram_mem[75721] = 16'b0000000000000000;
	sram_mem[75722] = 16'b0000000000000000;
	sram_mem[75723] = 16'b0000000000000000;
	sram_mem[75724] = 16'b0000000000000000;
	sram_mem[75725] = 16'b0000000000000000;
	sram_mem[75726] = 16'b0000000000000000;
	sram_mem[75727] = 16'b0000000000000000;
	sram_mem[75728] = 16'b0000000000000000;
	sram_mem[75729] = 16'b0000000000000000;
	sram_mem[75730] = 16'b0000000000000000;
	sram_mem[75731] = 16'b0000000000000000;
	sram_mem[75732] = 16'b0000000000000000;
	sram_mem[75733] = 16'b0000000000000000;
	sram_mem[75734] = 16'b0000000000000000;
	sram_mem[75735] = 16'b0000000000000000;
	sram_mem[75736] = 16'b0000000000000000;
	sram_mem[75737] = 16'b0000000000000000;
	sram_mem[75738] = 16'b0000000000000000;
	sram_mem[75739] = 16'b0000000000000000;
	sram_mem[75740] = 16'b0000000000000000;
	sram_mem[75741] = 16'b0000000000000000;
	sram_mem[75742] = 16'b0000000000000000;
	sram_mem[75743] = 16'b0000000000000000;
	sram_mem[75744] = 16'b0000000000000000;
	sram_mem[75745] = 16'b0000000000000000;
	sram_mem[75746] = 16'b0000000000000000;
	sram_mem[75747] = 16'b0000000000000000;
	sram_mem[75748] = 16'b0000000000000000;
	sram_mem[75749] = 16'b0000000000000000;
	sram_mem[75750] = 16'b0000000000000000;
	sram_mem[75751] = 16'b0000000000000000;
	sram_mem[75752] = 16'b0000000000000000;
	sram_mem[75753] = 16'b0000000000000000;
	sram_mem[75754] = 16'b0000000000000000;
	sram_mem[75755] = 16'b0000000000000000;
	sram_mem[75756] = 16'b0000000000000000;
	sram_mem[75757] = 16'b0000000000000000;
	sram_mem[75758] = 16'b0000000000000000;
	sram_mem[75759] = 16'b0000000000000000;
	sram_mem[75760] = 16'b0000000000000000;
	sram_mem[75761] = 16'b0000000000000000;
	sram_mem[75762] = 16'b0000000000000000;
	sram_mem[75763] = 16'b0000000000000000;
	sram_mem[75764] = 16'b0000000000000000;
	sram_mem[75765] = 16'b0000000000000000;
	sram_mem[75766] = 16'b0000000000000000;
	sram_mem[75767] = 16'b0000000000000000;
	sram_mem[75768] = 16'b0000000000000000;
	sram_mem[75769] = 16'b0000000000000000;
	sram_mem[75770] = 16'b0000000000000000;
	sram_mem[75771] = 16'b0000000000000000;
	sram_mem[75772] = 16'b0000000000000000;
	sram_mem[75773] = 16'b0000000000000000;
	sram_mem[75774] = 16'b0000000000000000;
	sram_mem[75775] = 16'b0000000000000000;
	sram_mem[75776] = 16'b0000000000000000;
	sram_mem[75777] = 16'b0000000000000000;
	sram_mem[75778] = 16'b0000000000000000;
	sram_mem[75779] = 16'b0000000000000000;
	sram_mem[75780] = 16'b0000000000000000;
	sram_mem[75781] = 16'b0000000000000000;
	sram_mem[75782] = 16'b0000000000000000;
	sram_mem[75783] = 16'b0000000000000000;
	sram_mem[75784] = 16'b0000000000000000;
	sram_mem[75785] = 16'b0000000000000000;
	sram_mem[75786] = 16'b0000000000000000;
	sram_mem[75787] = 16'b0000000000000000;
	sram_mem[75788] = 16'b0000000000000000;
	sram_mem[75789] = 16'b0000000000000000;
	sram_mem[75790] = 16'b0000000000000000;
	sram_mem[75791] = 16'b0000000000000000;
	sram_mem[75792] = 16'b0000000000000000;
	sram_mem[75793] = 16'b0000000000000000;
	sram_mem[75794] = 16'b0000000000000000;
	sram_mem[75795] = 16'b0000000000000000;
	sram_mem[75796] = 16'b0000000000000000;
	sram_mem[75797] = 16'b0000000000000000;
	sram_mem[75798] = 16'b0000000000000000;
	sram_mem[75799] = 16'b0000000000000000;
	sram_mem[75800] = 16'b0000000000000000;
	sram_mem[75801] = 16'b0000000000000000;
	sram_mem[75802] = 16'b0000000000000000;
	sram_mem[75803] = 16'b0000000000000000;
	sram_mem[75804] = 16'b0000000000000000;
	sram_mem[75805] = 16'b0000000000000000;
	sram_mem[75806] = 16'b0000000000000000;
	sram_mem[75807] = 16'b0000000000000000;
	sram_mem[75808] = 16'b0000000000000000;
	sram_mem[75809] = 16'b0000000000000000;
	sram_mem[75810] = 16'b0000000000000000;
	sram_mem[75811] = 16'b0000000000000000;
	sram_mem[75812] = 16'b0000000000000000;
	sram_mem[75813] = 16'b0000000000000000;
	sram_mem[75814] = 16'b0000000000000000;
	sram_mem[75815] = 16'b0000000000000000;
	sram_mem[75816] = 16'b0000000000000000;
	sram_mem[75817] = 16'b0000000000000000;
	sram_mem[75818] = 16'b0000000000000000;
	sram_mem[75819] = 16'b0000000000000000;
	sram_mem[75820] = 16'b0000000000000000;
	sram_mem[75821] = 16'b0000000000000000;
	sram_mem[75822] = 16'b0000000000000000;
	sram_mem[75823] = 16'b0000000000000000;
	sram_mem[75824] = 16'b0000000000000000;
	sram_mem[75825] = 16'b0000000000000000;
	sram_mem[75826] = 16'b0000000000000000;
	sram_mem[75827] = 16'b0000000000000000;
	sram_mem[75828] = 16'b0000000000000000;
	sram_mem[75829] = 16'b0000000000000000;
	sram_mem[75830] = 16'b0000000000000000;
	sram_mem[75831] = 16'b0000000000000000;
	sram_mem[75832] = 16'b0000000000000000;
	sram_mem[75833] = 16'b0000000000000000;
	sram_mem[75834] = 16'b0000000000000000;
	sram_mem[75835] = 16'b0000000000000000;
	sram_mem[75836] = 16'b0000000000000000;
	sram_mem[75837] = 16'b0000000000000000;
	sram_mem[75838] = 16'b0000000000000000;
	sram_mem[75839] = 16'b0000000000000000;
	sram_mem[75840] = 16'b0000000000000000;
	sram_mem[75841] = 16'b0000000000000000;
	sram_mem[75842] = 16'b0000000000000000;
	sram_mem[75843] = 16'b0000000000000000;
	sram_mem[75844] = 16'b0000000000000000;
	sram_mem[75845] = 16'b0000000000000000;
	sram_mem[75846] = 16'b0000000000000000;
	sram_mem[75847] = 16'b0000000000000000;
	sram_mem[75848] = 16'b0000000000000000;
	sram_mem[75849] = 16'b0000000000000000;
	sram_mem[75850] = 16'b0000000000000000;
	sram_mem[75851] = 16'b0000000000000000;
	sram_mem[75852] = 16'b0000000000000000;
	sram_mem[75853] = 16'b0000000000000000;
	sram_mem[75854] = 16'b0000000000000000;
	sram_mem[75855] = 16'b0000000000000000;
	sram_mem[75856] = 16'b0000000000000000;
	sram_mem[75857] = 16'b0000000000000000;
	sram_mem[75858] = 16'b0000000000000000;
	sram_mem[75859] = 16'b0000000000000000;
	sram_mem[75860] = 16'b0000000000000000;
	sram_mem[75861] = 16'b0000000000000000;
	sram_mem[75862] = 16'b0000000000000000;
	sram_mem[75863] = 16'b0000000000000000;
	sram_mem[75864] = 16'b0000000000000000;
	sram_mem[75865] = 16'b0000000000000000;
	sram_mem[75866] = 16'b0000000000000000;
	sram_mem[75867] = 16'b0000000000000000;
	sram_mem[75868] = 16'b0000000000000000;
	sram_mem[75869] = 16'b0000000000000000;
	sram_mem[75870] = 16'b0000000000000000;
	sram_mem[75871] = 16'b0000000000000000;
	sram_mem[75872] = 16'b0000000000000000;
	sram_mem[75873] = 16'b0000000000000000;
	sram_mem[75874] = 16'b0000000000000000;
	sram_mem[75875] = 16'b0000000000000000;
	sram_mem[75876] = 16'b0000000000000000;
	sram_mem[75877] = 16'b0000000000000000;
	sram_mem[75878] = 16'b0000000000000000;
	sram_mem[75879] = 16'b0000000000000000;
	sram_mem[75880] = 16'b0000000000000000;
	sram_mem[75881] = 16'b0000000000000000;
	sram_mem[75882] = 16'b0000000000000000;
	sram_mem[75883] = 16'b0000000000000000;
	sram_mem[75884] = 16'b0000000000000000;
	sram_mem[75885] = 16'b0000000000000000;
	sram_mem[75886] = 16'b0000000000000000;
	sram_mem[75887] = 16'b0000000000000000;
	sram_mem[75888] = 16'b0000000000000000;
	sram_mem[75889] = 16'b0000000000000000;
	sram_mem[75890] = 16'b0000000000000000;
	sram_mem[75891] = 16'b0000000000000000;
	sram_mem[75892] = 16'b0000000000000000;
	sram_mem[75893] = 16'b0000000000000000;
	sram_mem[75894] = 16'b0000000000000000;
	sram_mem[75895] = 16'b0000000000000000;
	sram_mem[75896] = 16'b0000000000000000;
	sram_mem[75897] = 16'b0000000000000000;
	sram_mem[75898] = 16'b0000000000000000;
	sram_mem[75899] = 16'b0000000000000000;
	sram_mem[75900] = 16'b0000000000000000;
	sram_mem[75901] = 16'b0000000000000000;
	sram_mem[75902] = 16'b0000000000000000;
	sram_mem[75903] = 16'b0000000000000000;
	sram_mem[75904] = 16'b0000000000000000;
	sram_mem[75905] = 16'b0000000000000000;
	sram_mem[75906] = 16'b0000000000000000;
	sram_mem[75907] = 16'b0000000000000000;
	sram_mem[75908] = 16'b0000000000000000;
	sram_mem[75909] = 16'b0000000000000000;
	sram_mem[75910] = 16'b0000000000000000;
	sram_mem[75911] = 16'b0000000000000000;
	sram_mem[75912] = 16'b0000000000000000;
	sram_mem[75913] = 16'b0000000000000000;
	sram_mem[75914] = 16'b0000000000000000;
	sram_mem[75915] = 16'b0000000000000000;
	sram_mem[75916] = 16'b0000000000000000;
	sram_mem[75917] = 16'b0000000000000000;
	sram_mem[75918] = 16'b0000000000000000;
	sram_mem[75919] = 16'b0000000000000000;
	sram_mem[75920] = 16'b0000000000000000;
	sram_mem[75921] = 16'b0000000000000000;
	sram_mem[75922] = 16'b0000000000000000;
	sram_mem[75923] = 16'b0000000000000000;
	sram_mem[75924] = 16'b0000000000000000;
	sram_mem[75925] = 16'b0000000000000000;
	sram_mem[75926] = 16'b0000000000000000;
	sram_mem[75927] = 16'b0000000000000000;
	sram_mem[75928] = 16'b0000000000000000;
	sram_mem[75929] = 16'b0000000000000000;
	sram_mem[75930] = 16'b0000000000000000;
	sram_mem[75931] = 16'b0000000000000000;
	sram_mem[75932] = 16'b0000000000000000;
	sram_mem[75933] = 16'b0000000000000000;
	sram_mem[75934] = 16'b0000000000000000;
	sram_mem[75935] = 16'b0000000000000000;
	sram_mem[75936] = 16'b0000000000000000;
	sram_mem[75937] = 16'b0000000000000000;
	sram_mem[75938] = 16'b0000000000000000;
	sram_mem[75939] = 16'b0000000000000000;
	sram_mem[75940] = 16'b0000000000000000;
	sram_mem[75941] = 16'b0000000000000000;
	sram_mem[75942] = 16'b0000000000000000;
	sram_mem[75943] = 16'b0000000000000000;
	sram_mem[75944] = 16'b0000000000000000;
	sram_mem[75945] = 16'b0000000000000000;
	sram_mem[75946] = 16'b0000000000000000;
	sram_mem[75947] = 16'b0000000000000000;
	sram_mem[75948] = 16'b0000000000000000;
	sram_mem[75949] = 16'b0000000000000000;
	sram_mem[75950] = 16'b0000000000000000;
	sram_mem[75951] = 16'b0000000000000000;
	sram_mem[75952] = 16'b0000000000000000;
	sram_mem[75953] = 16'b0000000000000000;
	sram_mem[75954] = 16'b0000000000000000;
	sram_mem[75955] = 16'b0000000000000000;
	sram_mem[75956] = 16'b0000000000000000;
	sram_mem[75957] = 16'b0000000000000000;
	sram_mem[75958] = 16'b0000000000000000;
	sram_mem[75959] = 16'b0000000000000000;
	sram_mem[75960] = 16'b0000000000000000;
	sram_mem[75961] = 16'b0000000000000000;
	sram_mem[75962] = 16'b0000000000000000;
	sram_mem[75963] = 16'b0000000000000000;
	sram_mem[75964] = 16'b0000000000000000;
	sram_mem[75965] = 16'b0000000000000000;
	sram_mem[75966] = 16'b0000000000000000;
	sram_mem[75967] = 16'b0000000000000000;
	sram_mem[75968] = 16'b0000000000000000;
	sram_mem[75969] = 16'b0000000000000000;
	sram_mem[75970] = 16'b0000000000000000;
	sram_mem[75971] = 16'b0000000000000000;
	sram_mem[75972] = 16'b0000000000000000;
	sram_mem[75973] = 16'b0000000000000000;
	sram_mem[75974] = 16'b0000000000000000;
	sram_mem[75975] = 16'b0000000000000000;
	sram_mem[75976] = 16'b0000000000000000;
	sram_mem[75977] = 16'b0000000000000000;
	sram_mem[75978] = 16'b0000000000000000;
	sram_mem[75979] = 16'b0000000000000000;
	sram_mem[75980] = 16'b0000000000000000;
	sram_mem[75981] = 16'b0000000000000000;
	sram_mem[75982] = 16'b0000000000000000;
	sram_mem[75983] = 16'b0000000000000000;
	sram_mem[75984] = 16'b0000000000000000;
	sram_mem[75985] = 16'b0000000000000000;
	sram_mem[75986] = 16'b0000000000000000;
	sram_mem[75987] = 16'b0000000000000000;
	sram_mem[75988] = 16'b0000000000000000;
	sram_mem[75989] = 16'b0000000000000000;
	sram_mem[75990] = 16'b0000000000000000;
	sram_mem[75991] = 16'b0000000000000000;
	sram_mem[75992] = 16'b0000000000000000;
	sram_mem[75993] = 16'b0000000000000000;
	sram_mem[75994] = 16'b0000000000000000;
	sram_mem[75995] = 16'b0000000000000000;
	sram_mem[75996] = 16'b0000000000000000;
	sram_mem[75997] = 16'b0000000000000000;
	sram_mem[75998] = 16'b0000000000000000;
	sram_mem[75999] = 16'b0000000000000000;
	sram_mem[76000] = 16'b0000000000000000;
	sram_mem[76001] = 16'b0000000000000000;
	sram_mem[76002] = 16'b0000000000000000;
	sram_mem[76003] = 16'b0000000000000000;
	sram_mem[76004] = 16'b0000000000000000;
	sram_mem[76005] = 16'b0000000000000000;
	sram_mem[76006] = 16'b0000000000000000;
	sram_mem[76007] = 16'b0000000000000000;
	sram_mem[76008] = 16'b0000000000000000;
	sram_mem[76009] = 16'b0000000000000000;
	sram_mem[76010] = 16'b0000000000000000;
	sram_mem[76011] = 16'b0000000000000000;
	sram_mem[76012] = 16'b0000000000000000;
	sram_mem[76013] = 16'b0000000000000000;
	sram_mem[76014] = 16'b0000000000000000;
	sram_mem[76015] = 16'b0000000000000000;
	sram_mem[76016] = 16'b0000000000000000;
	sram_mem[76017] = 16'b0000000000000000;
	sram_mem[76018] = 16'b0000000000000000;
	sram_mem[76019] = 16'b0000000000000000;
	sram_mem[76020] = 16'b0000000000000000;
	sram_mem[76021] = 16'b0000000000000000;
	sram_mem[76022] = 16'b0000000000000000;
	sram_mem[76023] = 16'b0000000000000000;
	sram_mem[76024] = 16'b0000000000000000;
	sram_mem[76025] = 16'b0000000000000000;
	sram_mem[76026] = 16'b0000000000000000;
	sram_mem[76027] = 16'b0000000000000000;
	sram_mem[76028] = 16'b0000000000000000;
	sram_mem[76029] = 16'b0000000000000000;
	sram_mem[76030] = 16'b0000000000000000;
	sram_mem[76031] = 16'b0000000000000000;
	sram_mem[76032] = 16'b0000000000000000;
	sram_mem[76033] = 16'b0000000000000000;
	sram_mem[76034] = 16'b0000000000000000;
	sram_mem[76035] = 16'b0000000000000000;
	sram_mem[76036] = 16'b0000000000000000;
	sram_mem[76037] = 16'b0000000000000000;
	sram_mem[76038] = 16'b0000000000000000;
	sram_mem[76039] = 16'b0000000000000000;
	sram_mem[76040] = 16'b0000000000000000;
	sram_mem[76041] = 16'b0000000000000000;
	sram_mem[76042] = 16'b0000000000000000;
	sram_mem[76043] = 16'b0000000000000000;
	sram_mem[76044] = 16'b0000000000000000;
	sram_mem[76045] = 16'b0000000000000000;
	sram_mem[76046] = 16'b0000000000000000;
	sram_mem[76047] = 16'b0000000000000000;
	sram_mem[76048] = 16'b0000000000000000;
	sram_mem[76049] = 16'b0000000000000000;
	sram_mem[76050] = 16'b0000000000000000;
	sram_mem[76051] = 16'b0000000000000000;
	sram_mem[76052] = 16'b0000000000000000;
	sram_mem[76053] = 16'b0000000000000000;
	sram_mem[76054] = 16'b0000000000000000;
	sram_mem[76055] = 16'b0000000000000000;
	sram_mem[76056] = 16'b0000000000000000;
	sram_mem[76057] = 16'b0000000000000000;
	sram_mem[76058] = 16'b0000000000000000;
	sram_mem[76059] = 16'b0000000000000000;
	sram_mem[76060] = 16'b0000000000000000;
	sram_mem[76061] = 16'b0000000000000000;
	sram_mem[76062] = 16'b0000000000000000;
	sram_mem[76063] = 16'b0000000000000000;
	sram_mem[76064] = 16'b0000000000000000;
	sram_mem[76065] = 16'b0000000000000000;
	sram_mem[76066] = 16'b0000000000000000;
	sram_mem[76067] = 16'b0000000000000000;
	sram_mem[76068] = 16'b0000000000000000;
	sram_mem[76069] = 16'b0000000000000000;
	sram_mem[76070] = 16'b0000000000000000;
	sram_mem[76071] = 16'b0000000000000000;
	sram_mem[76072] = 16'b0000000000000000;
	sram_mem[76073] = 16'b0000000000000000;
	sram_mem[76074] = 16'b0000000000000000;
	sram_mem[76075] = 16'b0000000000000000;
	sram_mem[76076] = 16'b0000000000000000;
	sram_mem[76077] = 16'b0000000000000000;
	sram_mem[76078] = 16'b0000000000000000;
	sram_mem[76079] = 16'b0000000000000000;
	sram_mem[76080] = 16'b0000000000000000;
	sram_mem[76081] = 16'b0000000000000000;
	sram_mem[76082] = 16'b0000000000000000;
	sram_mem[76083] = 16'b0000000000000000;
	sram_mem[76084] = 16'b0000000000000000;
	sram_mem[76085] = 16'b0000000000000000;
	sram_mem[76086] = 16'b0000000000000000;
	sram_mem[76087] = 16'b0000000000000000;
	sram_mem[76088] = 16'b0000000000000000;
	sram_mem[76089] = 16'b0000000000000000;
	sram_mem[76090] = 16'b0000000000000000;
	sram_mem[76091] = 16'b0000000000000000;
	sram_mem[76092] = 16'b0000000000000000;
	sram_mem[76093] = 16'b0000000000000000;
	sram_mem[76094] = 16'b0000000000000000;
	sram_mem[76095] = 16'b0000000000000000;
	sram_mem[76096] = 16'b0000000000000000;
	sram_mem[76097] = 16'b0000000000000000;
	sram_mem[76098] = 16'b0000000000000000;
	sram_mem[76099] = 16'b0000000000000000;
	sram_mem[76100] = 16'b0000000000000000;
	sram_mem[76101] = 16'b0000000000000000;
	sram_mem[76102] = 16'b0000000000000000;
	sram_mem[76103] = 16'b0000000000000000;
	sram_mem[76104] = 16'b0000000000000000;
	sram_mem[76105] = 16'b0000000000000000;
	sram_mem[76106] = 16'b0000000000000000;
	sram_mem[76107] = 16'b0000000000000000;
	sram_mem[76108] = 16'b0000000000000000;
	sram_mem[76109] = 16'b0000000000000000;
	sram_mem[76110] = 16'b0000000000000000;
	sram_mem[76111] = 16'b0000000000000000;
	sram_mem[76112] = 16'b0000000000000000;
	sram_mem[76113] = 16'b0000000000000000;
	sram_mem[76114] = 16'b0000000000000000;
	sram_mem[76115] = 16'b0000000000000000;
	sram_mem[76116] = 16'b0000000000000000;
	sram_mem[76117] = 16'b0000000000000000;
	sram_mem[76118] = 16'b0000000000000000;
	sram_mem[76119] = 16'b0000000000000000;
	sram_mem[76120] = 16'b0000000000000000;
	sram_mem[76121] = 16'b0000000000000000;
	sram_mem[76122] = 16'b0000000000000000;
	sram_mem[76123] = 16'b0000000000000000;
	sram_mem[76124] = 16'b0000000000000000;
	sram_mem[76125] = 16'b0000000000000000;
	sram_mem[76126] = 16'b0000000000000000;
	sram_mem[76127] = 16'b0000000000000000;
	sram_mem[76128] = 16'b0000000000000000;
	sram_mem[76129] = 16'b0000000000000000;
	sram_mem[76130] = 16'b0000000000000000;
	sram_mem[76131] = 16'b0000000000000000;
	sram_mem[76132] = 16'b0000000000000000;
	sram_mem[76133] = 16'b0000000000000000;
	sram_mem[76134] = 16'b0000000000000000;
	sram_mem[76135] = 16'b0000000000000000;
	sram_mem[76136] = 16'b0000000000000000;
	sram_mem[76137] = 16'b0000000000000000;
	sram_mem[76138] = 16'b0000000000000000;
	sram_mem[76139] = 16'b0000000000000000;
	sram_mem[76140] = 16'b0000000000000000;
	sram_mem[76141] = 16'b0000000000000000;
	sram_mem[76142] = 16'b0000000000000000;
	sram_mem[76143] = 16'b0000000000000000;
	sram_mem[76144] = 16'b0000000000000000;
	sram_mem[76145] = 16'b0000000000000000;
	sram_mem[76146] = 16'b0000000000000000;
	sram_mem[76147] = 16'b0000000000000000;
	sram_mem[76148] = 16'b0000000000000000;
	sram_mem[76149] = 16'b0000000000000000;
	sram_mem[76150] = 16'b0000000000000000;
	sram_mem[76151] = 16'b0000000000000000;
	sram_mem[76152] = 16'b0000000000000000;
	sram_mem[76153] = 16'b0000000000000000;
	sram_mem[76154] = 16'b0000000000000000;
	sram_mem[76155] = 16'b0000000000000000;
	sram_mem[76156] = 16'b0000000000000000;
	sram_mem[76157] = 16'b0000000000000000;
	sram_mem[76158] = 16'b0000000000000000;
	sram_mem[76159] = 16'b0000000000000000;
	sram_mem[76160] = 16'b0000000000000000;
	sram_mem[76161] = 16'b0000000000000000;
	sram_mem[76162] = 16'b0000000000000000;
	sram_mem[76163] = 16'b0000000000000000;
	sram_mem[76164] = 16'b0000000000000000;
	sram_mem[76165] = 16'b0000000000000000;
	sram_mem[76166] = 16'b0000000000000000;
	sram_mem[76167] = 16'b0000000000000000;
	sram_mem[76168] = 16'b0000000000000000;
	sram_mem[76169] = 16'b0000000000000000;
	sram_mem[76170] = 16'b0000000000000000;
	sram_mem[76171] = 16'b0000000000000000;
	sram_mem[76172] = 16'b0000000000000000;
	sram_mem[76173] = 16'b0000000000000000;
	sram_mem[76174] = 16'b0000000000000000;
	sram_mem[76175] = 16'b0000000000000000;
	sram_mem[76176] = 16'b0000000000000000;
	sram_mem[76177] = 16'b0000000000000000;
	sram_mem[76178] = 16'b0000000000000000;
	sram_mem[76179] = 16'b0000000000000000;
	sram_mem[76180] = 16'b0000000000000000;
	sram_mem[76181] = 16'b0000000000000000;
	sram_mem[76182] = 16'b0000000000000000;
	sram_mem[76183] = 16'b0000000000000000;
	sram_mem[76184] = 16'b0000000000000000;
	sram_mem[76185] = 16'b0000000000000000;
	sram_mem[76186] = 16'b0000000000000000;
	sram_mem[76187] = 16'b0000000000000000;
	sram_mem[76188] = 16'b0000000000000000;
	sram_mem[76189] = 16'b0000000000000000;
	sram_mem[76190] = 16'b0000000000000000;
	sram_mem[76191] = 16'b0000000000000000;
	sram_mem[76192] = 16'b0000000000000000;
	sram_mem[76193] = 16'b0000000000000000;
	sram_mem[76194] = 16'b0000000000000000;
	sram_mem[76195] = 16'b0000000000000000;
	sram_mem[76196] = 16'b0000000000000000;
	sram_mem[76197] = 16'b0000000000000000;
	sram_mem[76198] = 16'b0000000000000000;
	sram_mem[76199] = 16'b0000000000000000;
	sram_mem[76200] = 16'b0000000000000000;
	sram_mem[76201] = 16'b0000000000000000;
	sram_mem[76202] = 16'b0000000000000000;
	sram_mem[76203] = 16'b0000000000000000;
	sram_mem[76204] = 16'b0000000000000000;
	sram_mem[76205] = 16'b0000000000000000;
	sram_mem[76206] = 16'b0000000000000000;
	sram_mem[76207] = 16'b0000000000000000;
	sram_mem[76208] = 16'b0000000000000000;
	sram_mem[76209] = 16'b0000000000000000;
	sram_mem[76210] = 16'b0000000000000000;
	sram_mem[76211] = 16'b0000000000000000;
	sram_mem[76212] = 16'b0000000000000000;
	sram_mem[76213] = 16'b0000000000000000;
	sram_mem[76214] = 16'b0000000000000000;
	sram_mem[76215] = 16'b0000000000000000;
	sram_mem[76216] = 16'b0000000000000000;
	sram_mem[76217] = 16'b0000000000000000;
	sram_mem[76218] = 16'b0000000000000000;
	sram_mem[76219] = 16'b0000000000000000;
	sram_mem[76220] = 16'b0000000000000000;
	sram_mem[76221] = 16'b0000000000000000;
	sram_mem[76222] = 16'b0000000000000000;
	sram_mem[76223] = 16'b0000000000000000;
	sram_mem[76224] = 16'b0000000000000000;
	sram_mem[76225] = 16'b0000000000000000;
	sram_mem[76226] = 16'b0000000000000000;
	sram_mem[76227] = 16'b0000000000000000;
	sram_mem[76228] = 16'b0000000000000000;
	sram_mem[76229] = 16'b0000000000000000;
	sram_mem[76230] = 16'b0000000000000000;
	sram_mem[76231] = 16'b0000000000000000;
	sram_mem[76232] = 16'b0000000000000000;
	sram_mem[76233] = 16'b0000000000000000;
	sram_mem[76234] = 16'b0000000000000000;
	sram_mem[76235] = 16'b0000000000000000;
	sram_mem[76236] = 16'b0000000000000000;
	sram_mem[76237] = 16'b0000000000000000;
	sram_mem[76238] = 16'b0000000000000000;
	sram_mem[76239] = 16'b0000000000000000;
	sram_mem[76240] = 16'b0000000000000000;
	sram_mem[76241] = 16'b0000000000000000;
	sram_mem[76242] = 16'b0000000000000000;
	sram_mem[76243] = 16'b0000000000000000;
	sram_mem[76244] = 16'b0000000000000000;
	sram_mem[76245] = 16'b0000000000000000;
	sram_mem[76246] = 16'b0000000000000000;
	sram_mem[76247] = 16'b0000000000000000;
	sram_mem[76248] = 16'b0000000000000000;
	sram_mem[76249] = 16'b0000000000000000;
	sram_mem[76250] = 16'b0000000000000000;
	sram_mem[76251] = 16'b0000000000000000;
	sram_mem[76252] = 16'b0000000000000000;
	sram_mem[76253] = 16'b0000000000000000;
	sram_mem[76254] = 16'b0000000000000000;
	sram_mem[76255] = 16'b0000000000000000;
	sram_mem[76256] = 16'b0000000000000000;
	sram_mem[76257] = 16'b0000000000000000;
	sram_mem[76258] = 16'b0000000000000000;
	sram_mem[76259] = 16'b0000000000000000;
	sram_mem[76260] = 16'b0000000000000000;
	sram_mem[76261] = 16'b0000000000000000;
	sram_mem[76262] = 16'b0000000000000000;
	sram_mem[76263] = 16'b0000000000000000;
	sram_mem[76264] = 16'b0000000000000000;
	sram_mem[76265] = 16'b0000000000000000;
	sram_mem[76266] = 16'b0000000000000000;
	sram_mem[76267] = 16'b0000000000000000;
	sram_mem[76268] = 16'b0000000000000000;
	sram_mem[76269] = 16'b0000000000000000;
	sram_mem[76270] = 16'b0000000000000000;
	sram_mem[76271] = 16'b0000000000000000;
	sram_mem[76272] = 16'b0000000000000000;
	sram_mem[76273] = 16'b0000000000000000;
	sram_mem[76274] = 16'b0000000000000000;
	sram_mem[76275] = 16'b0000000000000000;
	sram_mem[76276] = 16'b0000000000000000;
	sram_mem[76277] = 16'b0000000000000000;
	sram_mem[76278] = 16'b0000000000000000;
	sram_mem[76279] = 16'b0000000000000000;
	sram_mem[76280] = 16'b0000000000000000;
	sram_mem[76281] = 16'b0000000000000000;
	sram_mem[76282] = 16'b0000000000000000;
	sram_mem[76283] = 16'b0000000000000000;
	sram_mem[76284] = 16'b0000000000000000;
	sram_mem[76285] = 16'b0000000000000000;
	sram_mem[76286] = 16'b0000000000000000;
	sram_mem[76287] = 16'b0000000000000000;
	sram_mem[76288] = 16'b0000000000000000;
	sram_mem[76289] = 16'b0000000000000000;
	sram_mem[76290] = 16'b0000000000000000;
	sram_mem[76291] = 16'b0000000000000000;
	sram_mem[76292] = 16'b0000000000000000;
	sram_mem[76293] = 16'b0000000000000000;
	sram_mem[76294] = 16'b0000000000000000;
	sram_mem[76295] = 16'b0000000000000000;
	sram_mem[76296] = 16'b0000000000000000;
	sram_mem[76297] = 16'b0000000000000000;
	sram_mem[76298] = 16'b0000000000000000;
	sram_mem[76299] = 16'b0000000000000000;
	sram_mem[76300] = 16'b0000000000000000;
	sram_mem[76301] = 16'b0000000000000000;
	sram_mem[76302] = 16'b0000000000000000;
	sram_mem[76303] = 16'b0000000000000000;
	sram_mem[76304] = 16'b0000000000000000;
	sram_mem[76305] = 16'b0000000000000000;
	sram_mem[76306] = 16'b0000000000000000;
	sram_mem[76307] = 16'b0000000000000000;
	sram_mem[76308] = 16'b0000000000000000;
	sram_mem[76309] = 16'b0000000000000000;
	sram_mem[76310] = 16'b0000000000000000;
	sram_mem[76311] = 16'b0000000000000000;
	sram_mem[76312] = 16'b0000000000000000;
	sram_mem[76313] = 16'b0000000000000000;
	sram_mem[76314] = 16'b0000000000000000;
	sram_mem[76315] = 16'b0000000000000000;
	sram_mem[76316] = 16'b0000000000000000;
	sram_mem[76317] = 16'b0000000000000000;
	sram_mem[76318] = 16'b0000000000000000;
	sram_mem[76319] = 16'b0000000000000000;
	sram_mem[76320] = 16'b0000000000000000;
	sram_mem[76321] = 16'b0000000000000000;
	sram_mem[76322] = 16'b0000000000000000;
	sram_mem[76323] = 16'b0000000000000000;
	sram_mem[76324] = 16'b0000000000000000;
	sram_mem[76325] = 16'b0000000000000000;
	sram_mem[76326] = 16'b0000000000000000;
	sram_mem[76327] = 16'b0000000000000000;
	sram_mem[76328] = 16'b0000000000000000;
	sram_mem[76329] = 16'b0000000000000000;
	sram_mem[76330] = 16'b0000000000000000;
	sram_mem[76331] = 16'b0000000000000000;
	sram_mem[76332] = 16'b0000000000000000;
	sram_mem[76333] = 16'b0000000000000000;
	sram_mem[76334] = 16'b0000000000000000;
	sram_mem[76335] = 16'b0000000000000000;
	sram_mem[76336] = 16'b0000000000000000;
	sram_mem[76337] = 16'b0000000000000000;
	sram_mem[76338] = 16'b0000000000000000;
	sram_mem[76339] = 16'b0000000000000000;
	sram_mem[76340] = 16'b0000000000000000;
	sram_mem[76341] = 16'b0000000000000000;
	sram_mem[76342] = 16'b0000000000000000;
	sram_mem[76343] = 16'b0000000000000000;
	sram_mem[76344] = 16'b0000000000000000;
	sram_mem[76345] = 16'b0000000000000000;
	sram_mem[76346] = 16'b0000000000000000;
	sram_mem[76347] = 16'b0000000000000000;
	sram_mem[76348] = 16'b0000000000000000;
	sram_mem[76349] = 16'b0000000000000000;
	sram_mem[76350] = 16'b0000000000000000;
	sram_mem[76351] = 16'b0000000000000000;
	sram_mem[76352] = 16'b0000000000000000;
	sram_mem[76353] = 16'b0000000000000000;
	sram_mem[76354] = 16'b0000000000000000;
	sram_mem[76355] = 16'b0000000000000000;
	sram_mem[76356] = 16'b0000000000000000;
	sram_mem[76357] = 16'b0000000000000000;
	sram_mem[76358] = 16'b0000000000000000;
	sram_mem[76359] = 16'b0000000000000000;
	sram_mem[76360] = 16'b0000000000000000;
	sram_mem[76361] = 16'b0000000000000000;
	sram_mem[76362] = 16'b0000000000000000;
	sram_mem[76363] = 16'b0000000000000000;
	sram_mem[76364] = 16'b0000000000000000;
	sram_mem[76365] = 16'b0000000000000000;
	sram_mem[76366] = 16'b0000000000000000;
	sram_mem[76367] = 16'b0000000000000000;
	sram_mem[76368] = 16'b0000000000000000;
	sram_mem[76369] = 16'b0000000000000000;
	sram_mem[76370] = 16'b0000000000000000;
	sram_mem[76371] = 16'b0000000000000000;
	sram_mem[76372] = 16'b0000000000000000;
	sram_mem[76373] = 16'b0000000000000000;
	sram_mem[76374] = 16'b0000000000000000;
	sram_mem[76375] = 16'b0000000000000000;
	sram_mem[76376] = 16'b0000000000000000;
	sram_mem[76377] = 16'b0000000000000000;
	sram_mem[76378] = 16'b0000000000000000;
	sram_mem[76379] = 16'b0000000000000000;
	sram_mem[76380] = 16'b0000000000000000;
	sram_mem[76381] = 16'b0000000000000000;
	sram_mem[76382] = 16'b0000000000000000;
	sram_mem[76383] = 16'b0000000000000000;
	sram_mem[76384] = 16'b0000000000000000;
	sram_mem[76385] = 16'b0000000000000000;
	sram_mem[76386] = 16'b0000000000000000;
	sram_mem[76387] = 16'b0000000000000000;
	sram_mem[76388] = 16'b0000000000000000;
	sram_mem[76389] = 16'b0000000000000000;
	sram_mem[76390] = 16'b0000000000000000;
	sram_mem[76391] = 16'b0000000000000000;
	sram_mem[76392] = 16'b0000000000000000;
	sram_mem[76393] = 16'b0000000000000000;
	sram_mem[76394] = 16'b0000000000000000;
	sram_mem[76395] = 16'b0000000000000000;
	sram_mem[76396] = 16'b0000000000000000;
	sram_mem[76397] = 16'b0000000000000000;
	sram_mem[76398] = 16'b0000000000000000;
	sram_mem[76399] = 16'b0000000000000000;
	sram_mem[76400] = 16'b0000000000000000;
	sram_mem[76401] = 16'b0000000000000000;
	sram_mem[76402] = 16'b0000000000000000;
	sram_mem[76403] = 16'b0000000000000000;
	sram_mem[76404] = 16'b0000000000000000;
	sram_mem[76405] = 16'b0000000000000000;
	sram_mem[76406] = 16'b0000000000000000;
	sram_mem[76407] = 16'b0000000000000000;
	sram_mem[76408] = 16'b0000000000000000;
	sram_mem[76409] = 16'b0000000000000000;
	sram_mem[76410] = 16'b0000000000000000;
	sram_mem[76411] = 16'b0000000000000000;
	sram_mem[76412] = 16'b0000000000000000;
	sram_mem[76413] = 16'b0000000000000000;
	sram_mem[76414] = 16'b0000000000000000;
	sram_mem[76415] = 16'b0000000000000000;
	sram_mem[76416] = 16'b0000000000000000;
	sram_mem[76417] = 16'b0000000000000000;
	sram_mem[76418] = 16'b0000000000000000;
	sram_mem[76419] = 16'b0000000000000000;
	sram_mem[76420] = 16'b0000000000000000;
	sram_mem[76421] = 16'b0000000000000000;
	sram_mem[76422] = 16'b0000000000000000;
	sram_mem[76423] = 16'b0000000000000000;
	sram_mem[76424] = 16'b0000000000000000;
	sram_mem[76425] = 16'b0000000000000000;
	sram_mem[76426] = 16'b0000000000000000;
	sram_mem[76427] = 16'b0000000000000000;
	sram_mem[76428] = 16'b0000000000000000;
	sram_mem[76429] = 16'b0000000000000000;
	sram_mem[76430] = 16'b0000000000000000;
	sram_mem[76431] = 16'b0000000000000000;
	sram_mem[76432] = 16'b0000000000000000;
	sram_mem[76433] = 16'b0000000000000000;
	sram_mem[76434] = 16'b0000000000000000;
	sram_mem[76435] = 16'b0000000000000000;
	sram_mem[76436] = 16'b0000000000000000;
	sram_mem[76437] = 16'b0000000000000000;
	sram_mem[76438] = 16'b0000000000000000;
	sram_mem[76439] = 16'b0000000000000000;
	sram_mem[76440] = 16'b0000000000000000;
	sram_mem[76441] = 16'b0000000000000000;
	sram_mem[76442] = 16'b0000000000000000;
	sram_mem[76443] = 16'b0000000000000000;
	sram_mem[76444] = 16'b0000000000000000;
	sram_mem[76445] = 16'b0000000000000000;
	sram_mem[76446] = 16'b0000000000000000;
	sram_mem[76447] = 16'b0000000000000000;
	sram_mem[76448] = 16'b0000000000000000;
	sram_mem[76449] = 16'b0000000000000000;
	sram_mem[76450] = 16'b0000000000000000;
	sram_mem[76451] = 16'b0000000000000000;
	sram_mem[76452] = 16'b0000000000000000;
	sram_mem[76453] = 16'b0000000000000000;
	sram_mem[76454] = 16'b0000000000000000;
	sram_mem[76455] = 16'b0000000000000000;
	sram_mem[76456] = 16'b0000000000000000;
	sram_mem[76457] = 16'b0000000000000000;
	sram_mem[76458] = 16'b0000000000000000;
	sram_mem[76459] = 16'b0000000000000000;
	sram_mem[76460] = 16'b0000000000000000;
	sram_mem[76461] = 16'b0000000000000000;
	sram_mem[76462] = 16'b0000000000000000;
	sram_mem[76463] = 16'b0000000000000000;
	sram_mem[76464] = 16'b0000000000000000;
	sram_mem[76465] = 16'b0000000000000000;
	sram_mem[76466] = 16'b0000000000000000;
	sram_mem[76467] = 16'b0000000000000000;
	sram_mem[76468] = 16'b0000000000000000;
	sram_mem[76469] = 16'b0000000000000000;
	sram_mem[76470] = 16'b0000000000000000;
	sram_mem[76471] = 16'b0000000000000000;
	sram_mem[76472] = 16'b0000000000000000;
	sram_mem[76473] = 16'b0000000000000000;
	sram_mem[76474] = 16'b0000000000000000;
	sram_mem[76475] = 16'b0000000000000000;
	sram_mem[76476] = 16'b0000000000000000;
	sram_mem[76477] = 16'b0000000000000000;
	sram_mem[76478] = 16'b0000000000000000;
	sram_mem[76479] = 16'b0000000000000000;
	sram_mem[76480] = 16'b0000000000000000;
	sram_mem[76481] = 16'b0000000000000000;
	sram_mem[76482] = 16'b0000000000000000;
	sram_mem[76483] = 16'b0000000000000000;
	sram_mem[76484] = 16'b0000000000000000;
	sram_mem[76485] = 16'b0000000000000000;
	sram_mem[76486] = 16'b0000000000000000;
	sram_mem[76487] = 16'b0000000000000000;
	sram_mem[76488] = 16'b0000000000000000;
	sram_mem[76489] = 16'b0000000000000000;
	sram_mem[76490] = 16'b0000000000000000;
	sram_mem[76491] = 16'b0000000000000000;
	sram_mem[76492] = 16'b0000000000000000;
	sram_mem[76493] = 16'b0000000000000000;
	sram_mem[76494] = 16'b0000000000000000;
	sram_mem[76495] = 16'b0000000000000000;
	sram_mem[76496] = 16'b0000000000000000;
	sram_mem[76497] = 16'b0000000000000000;
	sram_mem[76498] = 16'b0000000000000000;
	sram_mem[76499] = 16'b0000000000000000;
	sram_mem[76500] = 16'b0000000000000000;
	sram_mem[76501] = 16'b0000000000000000;
	sram_mem[76502] = 16'b0000000000000000;
	sram_mem[76503] = 16'b0000000000000000;
	sram_mem[76504] = 16'b0000000000000000;
	sram_mem[76505] = 16'b0000000000000000;
	sram_mem[76506] = 16'b0000000000000000;
	sram_mem[76507] = 16'b0000000000000000;
	sram_mem[76508] = 16'b0000000000000000;
	sram_mem[76509] = 16'b0000000000000000;
	sram_mem[76510] = 16'b0000000000000000;
	sram_mem[76511] = 16'b0000000000000000;
	sram_mem[76512] = 16'b0000000000000000;
	sram_mem[76513] = 16'b0000000000000000;
	sram_mem[76514] = 16'b0000000000000000;
	sram_mem[76515] = 16'b0000000000000000;
	sram_mem[76516] = 16'b0000000000000000;
	sram_mem[76517] = 16'b0000000000000000;
	sram_mem[76518] = 16'b0000000000000000;
	sram_mem[76519] = 16'b0000000000000000;
	sram_mem[76520] = 16'b0000000000000000;
	sram_mem[76521] = 16'b0000000000000000;
	sram_mem[76522] = 16'b0000000000000000;
	sram_mem[76523] = 16'b0000000000000000;
	sram_mem[76524] = 16'b0000000000000000;
	sram_mem[76525] = 16'b0000000000000000;
	sram_mem[76526] = 16'b0000000000000000;
	sram_mem[76527] = 16'b0000000000000000;
	sram_mem[76528] = 16'b0000000000000000;
	sram_mem[76529] = 16'b0000000000000000;
	sram_mem[76530] = 16'b0000000000000000;
	sram_mem[76531] = 16'b0000000000000000;
	sram_mem[76532] = 16'b0000000000000000;
	sram_mem[76533] = 16'b0000000000000000;
	sram_mem[76534] = 16'b0000000000000000;
	sram_mem[76535] = 16'b0000000000000000;
	sram_mem[76536] = 16'b0000000000000000;
	sram_mem[76537] = 16'b0000000000000000;
	sram_mem[76538] = 16'b0000000000000000;
	sram_mem[76539] = 16'b0000000000000000;
	sram_mem[76540] = 16'b0000000000000000;
	sram_mem[76541] = 16'b0000000000000000;
	sram_mem[76542] = 16'b0000000000000000;
	sram_mem[76543] = 16'b0000000000000000;
	sram_mem[76544] = 16'b0000000000000000;
	sram_mem[76545] = 16'b0000000000000000;
	sram_mem[76546] = 16'b0000000000000000;
	sram_mem[76547] = 16'b0000000000000000;
	sram_mem[76548] = 16'b0000000000000000;
	sram_mem[76549] = 16'b0000000000000000;
	sram_mem[76550] = 16'b0000000000000000;
	sram_mem[76551] = 16'b0000000000000000;
	sram_mem[76552] = 16'b0000000000000000;
	sram_mem[76553] = 16'b0000000000000000;
	sram_mem[76554] = 16'b0000000000000000;
	sram_mem[76555] = 16'b0000000000000000;
	sram_mem[76556] = 16'b0000000000000000;
	sram_mem[76557] = 16'b0000000000000000;
	sram_mem[76558] = 16'b0000000000000000;
	sram_mem[76559] = 16'b0000000000000000;
	sram_mem[76560] = 16'b0000000000000000;
	sram_mem[76561] = 16'b0000000000000000;
	sram_mem[76562] = 16'b0000000000000000;
	sram_mem[76563] = 16'b0000000000000000;
	sram_mem[76564] = 16'b0000000000000000;
	sram_mem[76565] = 16'b0000000000000000;
	sram_mem[76566] = 16'b0000000000000000;
	sram_mem[76567] = 16'b0000000000000000;
	sram_mem[76568] = 16'b0000000000000000;
	sram_mem[76569] = 16'b0000000000000000;
	sram_mem[76570] = 16'b0000000000000000;
	sram_mem[76571] = 16'b0000000000000000;
	sram_mem[76572] = 16'b0000000000000000;
	sram_mem[76573] = 16'b0000000000000000;
	sram_mem[76574] = 16'b0000000000000000;
	sram_mem[76575] = 16'b0000000000000000;
	sram_mem[76576] = 16'b0000000000000000;
	sram_mem[76577] = 16'b0000000000000000;
	sram_mem[76578] = 16'b0000000000000000;
	sram_mem[76579] = 16'b0000000000000000;
	sram_mem[76580] = 16'b0000000000000000;
	sram_mem[76581] = 16'b0000000000000000;
	sram_mem[76582] = 16'b0000000000000000;
	sram_mem[76583] = 16'b0000000000000000;
	sram_mem[76584] = 16'b0000000000000000;
	sram_mem[76585] = 16'b0000000000000000;
	sram_mem[76586] = 16'b0000000000000000;
	sram_mem[76587] = 16'b0000000000000000;
	sram_mem[76588] = 16'b0000000000000000;
	sram_mem[76589] = 16'b0000000000000000;
	sram_mem[76590] = 16'b0000000000000000;
	sram_mem[76591] = 16'b0000000000000000;
	sram_mem[76592] = 16'b0000000000000000;
	sram_mem[76593] = 16'b0000000000000000;
	sram_mem[76594] = 16'b0000000000000000;
	sram_mem[76595] = 16'b0000000000000000;
	sram_mem[76596] = 16'b0000000000000000;
	sram_mem[76597] = 16'b0000000000000000;
	sram_mem[76598] = 16'b0000000000000000;
	sram_mem[76599] = 16'b0000000000000000;
	sram_mem[76600] = 16'b0000000000000000;
	sram_mem[76601] = 16'b0000000000000000;
	sram_mem[76602] = 16'b0000000000000000;
	sram_mem[76603] = 16'b0000000000000000;
	sram_mem[76604] = 16'b0000000000000000;
	sram_mem[76605] = 16'b0000000000000000;
	sram_mem[76606] = 16'b0000000000000000;
	sram_mem[76607] = 16'b0000000000000000;
	sram_mem[76608] = 16'b0000000000000000;
	sram_mem[76609] = 16'b0000000000000000;
	sram_mem[76610] = 16'b0000000000000000;
	sram_mem[76611] = 16'b0000000000000000;
	sram_mem[76612] = 16'b0000000000000000;
	sram_mem[76613] = 16'b0000000000000000;
	sram_mem[76614] = 16'b0000000000000000;
	sram_mem[76615] = 16'b0000000000000000;
	sram_mem[76616] = 16'b0000000000000000;
	sram_mem[76617] = 16'b0000000000000000;
	sram_mem[76618] = 16'b0000000000000000;
	sram_mem[76619] = 16'b0000000000000000;
	sram_mem[76620] = 16'b0000000000000000;
	sram_mem[76621] = 16'b0000000000000000;
	sram_mem[76622] = 16'b0000000000000000;
	sram_mem[76623] = 16'b0000000000000000;
	sram_mem[76624] = 16'b0000000000000000;
	sram_mem[76625] = 16'b0000000000000000;
	sram_mem[76626] = 16'b0000000000000000;
	sram_mem[76627] = 16'b0000000000000000;
	sram_mem[76628] = 16'b0000000000000000;
	sram_mem[76629] = 16'b0000000000000000;
	sram_mem[76630] = 16'b0000000000000000;
	sram_mem[76631] = 16'b0000000000000000;
	sram_mem[76632] = 16'b0000000000000000;
	sram_mem[76633] = 16'b0000000000000000;
	sram_mem[76634] = 16'b0000000000000000;
	sram_mem[76635] = 16'b0000000000000000;
	sram_mem[76636] = 16'b0000000000000000;
	sram_mem[76637] = 16'b0000000000000000;
	sram_mem[76638] = 16'b0000000000000000;
	sram_mem[76639] = 16'b0000000000000000;
	sram_mem[76640] = 16'b0000000000000000;
	sram_mem[76641] = 16'b0000000000000000;
	sram_mem[76642] = 16'b0000000000000000;
	sram_mem[76643] = 16'b0000000000000000;
	sram_mem[76644] = 16'b0000000000000000;
	sram_mem[76645] = 16'b0000000000000000;
	sram_mem[76646] = 16'b0000000000000000;
	sram_mem[76647] = 16'b0000000000000000;
	sram_mem[76648] = 16'b0000000000000000;
	sram_mem[76649] = 16'b0000000000000000;
	sram_mem[76650] = 16'b0000000000000000;
	sram_mem[76651] = 16'b0000000000000000;
	sram_mem[76652] = 16'b0000000000000000;
	sram_mem[76653] = 16'b0000000000000000;
	sram_mem[76654] = 16'b0000000000000000;
	sram_mem[76655] = 16'b0000000000000000;
	sram_mem[76656] = 16'b0000000000000000;
	sram_mem[76657] = 16'b0000000000000000;
	sram_mem[76658] = 16'b0000000000000000;
	sram_mem[76659] = 16'b0000000000000000;
	sram_mem[76660] = 16'b0000000000000000;
	sram_mem[76661] = 16'b0000000000000000;
	sram_mem[76662] = 16'b0000000000000000;
	sram_mem[76663] = 16'b0000000000000000;
	sram_mem[76664] = 16'b0000000000000000;
	sram_mem[76665] = 16'b0000000000000000;
	sram_mem[76666] = 16'b0000000000000000;
	sram_mem[76667] = 16'b0000000000000000;
	sram_mem[76668] = 16'b0000000000000000;
	sram_mem[76669] = 16'b0000000000000000;
	sram_mem[76670] = 16'b0000000000000000;
	sram_mem[76671] = 16'b0000000000000000;
	sram_mem[76672] = 16'b0000000000000000;
	sram_mem[76673] = 16'b0000000000000000;
	sram_mem[76674] = 16'b0000000000000000;
	sram_mem[76675] = 16'b0000000000000000;
	sram_mem[76676] = 16'b0000000000000000;
	sram_mem[76677] = 16'b0000000000000000;
	sram_mem[76678] = 16'b0000000000000000;
	sram_mem[76679] = 16'b0000000000000000;
	sram_mem[76680] = 16'b0000000000000000;
	sram_mem[76681] = 16'b0000000000000000;
	sram_mem[76682] = 16'b0000000000000000;
	sram_mem[76683] = 16'b0000000000000000;
	sram_mem[76684] = 16'b0000000000000000;
	sram_mem[76685] = 16'b0000000000000000;
	sram_mem[76686] = 16'b0000000000000000;
	sram_mem[76687] = 16'b0000000000000000;
	sram_mem[76688] = 16'b0000000000000000;
	sram_mem[76689] = 16'b0000000000000000;
	sram_mem[76690] = 16'b0000000000000000;
	sram_mem[76691] = 16'b0000000000000000;
	sram_mem[76692] = 16'b0000000000000000;
	sram_mem[76693] = 16'b0000000000000000;
	sram_mem[76694] = 16'b0000000000000000;
	sram_mem[76695] = 16'b0000000000000000;
	sram_mem[76696] = 16'b0000000000000000;
	sram_mem[76697] = 16'b0000000000000000;
	sram_mem[76698] = 16'b0000000000000000;
	sram_mem[76699] = 16'b0000000000000000;
	sram_mem[76700] = 16'b0000000000000000;
	sram_mem[76701] = 16'b0000000000000000;
	sram_mem[76702] = 16'b0000000000000000;
	sram_mem[76703] = 16'b0000000000000000;
	sram_mem[76704] = 16'b0000000000000000;
	sram_mem[76705] = 16'b0000000000000000;
	sram_mem[76706] = 16'b0000000000000000;
	sram_mem[76707] = 16'b0000000000000000;
	sram_mem[76708] = 16'b0000000000000000;
	sram_mem[76709] = 16'b0000000000000000;
	sram_mem[76710] = 16'b0000000000000000;
	sram_mem[76711] = 16'b0000000000000000;
	sram_mem[76712] = 16'b0000000000000000;
	sram_mem[76713] = 16'b0000000000000000;
	sram_mem[76714] = 16'b0000000000000000;
	sram_mem[76715] = 16'b0000000000000000;
	sram_mem[76716] = 16'b0000000000000000;
	sram_mem[76717] = 16'b0000000000000000;
	sram_mem[76718] = 16'b0000000000000000;
	sram_mem[76719] = 16'b0000000000000000;
	sram_mem[76720] = 16'b0000000000000000;
	sram_mem[76721] = 16'b0000000000000000;
	sram_mem[76722] = 16'b0000000000000000;
	sram_mem[76723] = 16'b0000000000000000;
	sram_mem[76724] = 16'b0000000000000000;
	sram_mem[76725] = 16'b0000000000000000;
	sram_mem[76726] = 16'b0000000000000000;
	sram_mem[76727] = 16'b0000000000000000;
	sram_mem[76728] = 16'b0000000000000000;
	sram_mem[76729] = 16'b0000000000000000;
	sram_mem[76730] = 16'b0000000000000000;
	sram_mem[76731] = 16'b0000000000000000;
	sram_mem[76732] = 16'b0000000000000000;
	sram_mem[76733] = 16'b0000000000000000;
	sram_mem[76734] = 16'b0000000000000000;
	sram_mem[76735] = 16'b0000000000000000;
	sram_mem[76736] = 16'b0000000000000000;
	sram_mem[76737] = 16'b0000000000000000;
	sram_mem[76738] = 16'b0000000000000000;
	sram_mem[76739] = 16'b0000000000000000;
	sram_mem[76740] = 16'b0000000000000000;
	sram_mem[76741] = 16'b0000000000000000;
	sram_mem[76742] = 16'b0000000000000000;
	sram_mem[76743] = 16'b0000000000000000;
	sram_mem[76744] = 16'b0000000000000000;
	sram_mem[76745] = 16'b0000000000000000;
	sram_mem[76746] = 16'b0000000000000000;
	sram_mem[76747] = 16'b0000000000000000;
	sram_mem[76748] = 16'b0000000000000000;
	sram_mem[76749] = 16'b0000000000000000;
	sram_mem[76750] = 16'b0000000000000000;
	sram_mem[76751] = 16'b0000000000000000;
	sram_mem[76752] = 16'b0000000000000000;
	sram_mem[76753] = 16'b0000000000000000;
	sram_mem[76754] = 16'b0000000000000000;
	sram_mem[76755] = 16'b0000000000000000;
	sram_mem[76756] = 16'b0000000000000000;
	sram_mem[76757] = 16'b0000000000000000;
	sram_mem[76758] = 16'b0000000000000000;
	sram_mem[76759] = 16'b0000000000000000;
	sram_mem[76760] = 16'b0000000000000000;
	sram_mem[76761] = 16'b0000000000000000;
	sram_mem[76762] = 16'b0000000000000000;
	sram_mem[76763] = 16'b0000000000000000;
	sram_mem[76764] = 16'b0000000000000000;
	sram_mem[76765] = 16'b0000000000000000;
	sram_mem[76766] = 16'b0000000000000000;
	sram_mem[76767] = 16'b0000000000000000;
	sram_mem[76768] = 16'b0000000000000000;
	sram_mem[76769] = 16'b0000000000000000;
	sram_mem[76770] = 16'b0000000000000000;
	sram_mem[76771] = 16'b0000000000000000;
	sram_mem[76772] = 16'b0000000000000000;
	sram_mem[76773] = 16'b0000000000000000;
	sram_mem[76774] = 16'b0000000000000000;
	sram_mem[76775] = 16'b0000000000000000;
	sram_mem[76776] = 16'b0000000000000000;
	sram_mem[76777] = 16'b0000000000000000;
	sram_mem[76778] = 16'b0000000000000000;
	sram_mem[76779] = 16'b0000000000000000;
	sram_mem[76780] = 16'b0000000000000000;
	sram_mem[76781] = 16'b0000000000000000;
	sram_mem[76782] = 16'b0000000000000000;
	sram_mem[76783] = 16'b0000000000000000;
	sram_mem[76784] = 16'b0000000000000000;
	sram_mem[76785] = 16'b0000000000000000;
	sram_mem[76786] = 16'b0000000000000000;
	sram_mem[76787] = 16'b0000000000000000;
	sram_mem[76788] = 16'b0000000000000000;
	sram_mem[76789] = 16'b0000000000000000;
	sram_mem[76790] = 16'b0000000000000000;
	sram_mem[76791] = 16'b0000000000000000;
	sram_mem[76792] = 16'b0000000000000000;
	sram_mem[76793] = 16'b0000000000000000;
	sram_mem[76794] = 16'b0000000000000000;
	sram_mem[76795] = 16'b0000000000000000;
	sram_mem[76796] = 16'b0000000000000000;
	sram_mem[76797] = 16'b0000000000000000;
	sram_mem[76798] = 16'b0000000000000000;
	sram_mem[76799] = 16'b0000000000000000;
	sram_mem[76800] = 16'b0000000000000000;
	sram_mem[76801] = 16'b0000000000000000;
	sram_mem[76802] = 16'b0000000000000000;
	sram_mem[76803] = 16'b0000000000000000;
	sram_mem[76804] = 16'b0000000000000000;
	sram_mem[76805] = 16'b0000000000000000;
	sram_mem[76806] = 16'b0000000000000000;
	sram_mem[76807] = 16'b0000000000000000;
	sram_mem[76808] = 16'b0000000000000000;
	sram_mem[76809] = 16'b0000000000000000;
	sram_mem[76810] = 16'b0000000000000000;
	sram_mem[76811] = 16'b0000000000000000;
	sram_mem[76812] = 16'b0000000000000000;
	sram_mem[76813] = 16'b0000000000000000;
	sram_mem[76814] = 16'b0000000000000000;
	sram_mem[76815] = 16'b0000000000000000;
	sram_mem[76816] = 16'b0000000000000000;
	sram_mem[76817] = 16'b0000000000000000;
	sram_mem[76818] = 16'b0000000000000000;
	sram_mem[76819] = 16'b0000000000000000;
	sram_mem[76820] = 16'b0000000000000000;
	sram_mem[76821] = 16'b0000000000000000;
	sram_mem[76822] = 16'b0000000000000000;
	sram_mem[76823] = 16'b0000000000000000;
	sram_mem[76824] = 16'b0000000000000000;
	sram_mem[76825] = 16'b0000000000000000;
	sram_mem[76826] = 16'b0000000000000000;
	sram_mem[76827] = 16'b0000000000000000;
	sram_mem[76828] = 16'b0000000000000000;
	sram_mem[76829] = 16'b0000000000000000;
	sram_mem[76830] = 16'b0000000000000000;
	sram_mem[76831] = 16'b0000000000000000;
	sram_mem[76832] = 16'b0000000000000000;
	sram_mem[76833] = 16'b0000000000000000;
	sram_mem[76834] = 16'b0000000000000000;
	sram_mem[76835] = 16'b0000000000000000;
	sram_mem[76836] = 16'b0000000000000000;
	sram_mem[76837] = 16'b0000000000000000;
	sram_mem[76838] = 16'b0000000000000000;
	sram_mem[76839] = 16'b0000000000000000;
	sram_mem[76840] = 16'b0000000000000000;
	sram_mem[76841] = 16'b0000000000000000;
	sram_mem[76842] = 16'b0000000000000000;
	sram_mem[76843] = 16'b0000000000000000;
	sram_mem[76844] = 16'b0000000000000000;
	sram_mem[76845] = 16'b0000000000000000;
	sram_mem[76846] = 16'b0000000000000000;
	sram_mem[76847] = 16'b0000000000000000;
	sram_mem[76848] = 16'b0000000000000000;
	sram_mem[76849] = 16'b0000000000000000;
	sram_mem[76850] = 16'b0000000000000000;
	sram_mem[76851] = 16'b0000000000000000;
	sram_mem[76852] = 16'b0000000000000000;
	sram_mem[76853] = 16'b0000000000000000;
	sram_mem[76854] = 16'b0000000000000000;
	sram_mem[76855] = 16'b0000000000000000;
	sram_mem[76856] = 16'b0000000000000000;
	sram_mem[76857] = 16'b0000000000000000;
	sram_mem[76858] = 16'b0000000000000000;
	sram_mem[76859] = 16'b0000000000000000;
	sram_mem[76860] = 16'b0000000000000000;
	sram_mem[76861] = 16'b0000000000000000;
	sram_mem[76862] = 16'b0000000000000000;
	sram_mem[76863] = 16'b0000000000000000;
	sram_mem[76864] = 16'b0000000000000000;
	sram_mem[76865] = 16'b0000000000000000;
	sram_mem[76866] = 16'b0000000000000000;
	sram_mem[76867] = 16'b0000000000000000;
	sram_mem[76868] = 16'b0000000000000000;
	sram_mem[76869] = 16'b0000000000000000;
	sram_mem[76870] = 16'b0000000000000000;
	sram_mem[76871] = 16'b0000000000000000;
	sram_mem[76872] = 16'b0000000000000000;
	sram_mem[76873] = 16'b0000000000000000;
	sram_mem[76874] = 16'b0000000000000000;
	sram_mem[76875] = 16'b0000000000000000;
	sram_mem[76876] = 16'b0000000000000000;
	sram_mem[76877] = 16'b0000000000000000;
	sram_mem[76878] = 16'b0000000000000000;
	sram_mem[76879] = 16'b0000000000000000;
	sram_mem[76880] = 16'b0000000000000000;
	sram_mem[76881] = 16'b0000000000000000;
	sram_mem[76882] = 16'b0000000000000000;
	sram_mem[76883] = 16'b0000000000000000;
	sram_mem[76884] = 16'b0000000000000000;
	sram_mem[76885] = 16'b0000000000000000;
	sram_mem[76886] = 16'b0000000000000000;
	sram_mem[76887] = 16'b0000000000000000;
	sram_mem[76888] = 16'b0000000000000000;
	sram_mem[76889] = 16'b0000000000000000;
	sram_mem[76890] = 16'b0000000000000000;
	sram_mem[76891] = 16'b0000000000000000;
	sram_mem[76892] = 16'b0000000000000000;
	sram_mem[76893] = 16'b0000000000000000;
	sram_mem[76894] = 16'b0000000000000000;
	sram_mem[76895] = 16'b0000000000000000;
	sram_mem[76896] = 16'b0000000000000000;
	sram_mem[76897] = 16'b0000000000000000;
	sram_mem[76898] = 16'b0000000000000000;
	sram_mem[76899] = 16'b0000000000000000;
	sram_mem[76900] = 16'b0000000000000000;
	sram_mem[76901] = 16'b0000000000000000;
	sram_mem[76902] = 16'b0000000000000000;
	sram_mem[76903] = 16'b0000000000000000;
	sram_mem[76904] = 16'b0000000000000000;
	sram_mem[76905] = 16'b0000000000000000;
	sram_mem[76906] = 16'b0000000000000000;
	sram_mem[76907] = 16'b0000000000000000;
	sram_mem[76908] = 16'b0000000000000000;
	sram_mem[76909] = 16'b0000000000000000;
	sram_mem[76910] = 16'b0000000000000000;
	sram_mem[76911] = 16'b0000000000000000;
	sram_mem[76912] = 16'b0000000000000000;
	sram_mem[76913] = 16'b0000000000000000;
	sram_mem[76914] = 16'b0000000000000000;
	sram_mem[76915] = 16'b0000000000000000;
	sram_mem[76916] = 16'b0000000000000000;
	sram_mem[76917] = 16'b0000000000000000;
	sram_mem[76918] = 16'b0000000000000000;
	sram_mem[76919] = 16'b0000000000000000;
	sram_mem[76920] = 16'b0000000000000000;
	sram_mem[76921] = 16'b0000000000000000;
	sram_mem[76922] = 16'b0000000000000000;
	sram_mem[76923] = 16'b0000000000000000;
	sram_mem[76924] = 16'b0000000000000000;
	sram_mem[76925] = 16'b0000000000000000;
	sram_mem[76926] = 16'b0000000000000000;
	sram_mem[76927] = 16'b0000000000000000;
	sram_mem[76928] = 16'b0000000000000000;
	sram_mem[76929] = 16'b0000000000000000;
	sram_mem[76930] = 16'b0000000000000000;
	sram_mem[76931] = 16'b0000000000000000;
	sram_mem[76932] = 16'b0000000000000000;
	sram_mem[76933] = 16'b0000000000000000;
	sram_mem[76934] = 16'b0000000000000000;
	sram_mem[76935] = 16'b0000000000000000;
	sram_mem[76936] = 16'b0000000000000000;
	sram_mem[76937] = 16'b0000000000000000;
	sram_mem[76938] = 16'b0000000000000000;
	sram_mem[76939] = 16'b0000000000000000;
	sram_mem[76940] = 16'b0000000000000000;
	sram_mem[76941] = 16'b0000000000000000;
	sram_mem[76942] = 16'b0000000000000000;
	sram_mem[76943] = 16'b0000000000000000;
	sram_mem[76944] = 16'b0000000000000000;
	sram_mem[76945] = 16'b0000000000000000;
	sram_mem[76946] = 16'b0000000000000000;
	sram_mem[76947] = 16'b0000000000000000;
	sram_mem[76948] = 16'b0000000000000000;
	sram_mem[76949] = 16'b0000000000000000;
	sram_mem[76950] = 16'b0000000000000000;
	sram_mem[76951] = 16'b0000000000000000;
	sram_mem[76952] = 16'b0000000000000000;
	sram_mem[76953] = 16'b0000000000000000;
	sram_mem[76954] = 16'b0000000000000000;
	sram_mem[76955] = 16'b0000000000000000;
	sram_mem[76956] = 16'b0000000000000000;
	sram_mem[76957] = 16'b0000000000000000;
	sram_mem[76958] = 16'b0000000000000000;
	sram_mem[76959] = 16'b0000000000000000;
	sram_mem[76960] = 16'b0000000000000000;
	sram_mem[76961] = 16'b0000000000000000;
	sram_mem[76962] = 16'b0000000000000000;
	sram_mem[76963] = 16'b0000000000000000;
	sram_mem[76964] = 16'b0000000000000000;
	sram_mem[76965] = 16'b0000000000000000;
	sram_mem[76966] = 16'b0000000000000000;
	sram_mem[76967] = 16'b0000000000000000;
	sram_mem[76968] = 16'b0000000000000000;
	sram_mem[76969] = 16'b0000000000000000;
	sram_mem[76970] = 16'b0000000000000000;
	sram_mem[76971] = 16'b0000000000000000;
	sram_mem[76972] = 16'b0000000000000000;
	sram_mem[76973] = 16'b0000000000000000;
	sram_mem[76974] = 16'b0000000000000000;
	sram_mem[76975] = 16'b0000000000000000;
	sram_mem[76976] = 16'b0000000000000000;
	sram_mem[76977] = 16'b0000000000000000;
	sram_mem[76978] = 16'b0000000000000000;
	sram_mem[76979] = 16'b0000000000000000;
	sram_mem[76980] = 16'b0000000000000000;
	sram_mem[76981] = 16'b0000000000000000;
	sram_mem[76982] = 16'b0000000000000000;
	sram_mem[76983] = 16'b0000000000000000;
	sram_mem[76984] = 16'b0000000000000000;
	sram_mem[76985] = 16'b0000000000000000;
	sram_mem[76986] = 16'b0000000000000000;
	sram_mem[76987] = 16'b0000000000000000;
	sram_mem[76988] = 16'b0000000000000000;
	sram_mem[76989] = 16'b0000000000000000;
	sram_mem[76990] = 16'b0000000000000000;
	sram_mem[76991] = 16'b0000000000000000;
	sram_mem[76992] = 16'b0000000000000000;
	sram_mem[76993] = 16'b0000000000000000;
	sram_mem[76994] = 16'b0000000000000000;
	sram_mem[76995] = 16'b0000000000000000;
	sram_mem[76996] = 16'b0000000000000000;
	sram_mem[76997] = 16'b0000000000000000;
	sram_mem[76998] = 16'b0000000000000000;
	sram_mem[76999] = 16'b0000000000000000;
	sram_mem[77000] = 16'b0000000000000000;
	sram_mem[77001] = 16'b0000000000000000;
	sram_mem[77002] = 16'b0000000000000000;
	sram_mem[77003] = 16'b0000000000000000;
	sram_mem[77004] = 16'b0000000000000000;
	sram_mem[77005] = 16'b0000000000000000;
	sram_mem[77006] = 16'b0000000000000000;
	sram_mem[77007] = 16'b0000000000000000;
	sram_mem[77008] = 16'b0000000000000000;
	sram_mem[77009] = 16'b0000000000000000;
	sram_mem[77010] = 16'b0000000000000000;
	sram_mem[77011] = 16'b0000000000000000;
	sram_mem[77012] = 16'b0000000000000000;
	sram_mem[77013] = 16'b0000000000000000;
	sram_mem[77014] = 16'b0000000000000000;
	sram_mem[77015] = 16'b0000000000000000;
	sram_mem[77016] = 16'b0000000000000000;
	sram_mem[77017] = 16'b0000000000000000;
	sram_mem[77018] = 16'b0000000000000000;
	sram_mem[77019] = 16'b0000000000000000;
	sram_mem[77020] = 16'b0000000000000000;
	sram_mem[77021] = 16'b0000000000000000;
	sram_mem[77022] = 16'b0000000000000000;
	sram_mem[77023] = 16'b0000000000000000;
	sram_mem[77024] = 16'b0000000000000000;
	sram_mem[77025] = 16'b0000000000000000;
	sram_mem[77026] = 16'b0000000000000000;
	sram_mem[77027] = 16'b0000000000000000;
	sram_mem[77028] = 16'b0000000000000000;
	sram_mem[77029] = 16'b0000000000000000;
	sram_mem[77030] = 16'b0000000000000000;
	sram_mem[77031] = 16'b0000000000000000;
	sram_mem[77032] = 16'b0000000000000000;
	sram_mem[77033] = 16'b0000000000000000;
	sram_mem[77034] = 16'b0000000000000000;
	sram_mem[77035] = 16'b0000000000000000;
	sram_mem[77036] = 16'b0000000000000000;
	sram_mem[77037] = 16'b0000000000000000;
	sram_mem[77038] = 16'b0000000000000000;
	sram_mem[77039] = 16'b0000000000000000;
	sram_mem[77040] = 16'b0000000000000000;
	sram_mem[77041] = 16'b0000000000000000;
	sram_mem[77042] = 16'b0000000000000000;
	sram_mem[77043] = 16'b0000000000000000;
	sram_mem[77044] = 16'b0000000000000000;
	sram_mem[77045] = 16'b0000000000000000;
	sram_mem[77046] = 16'b0000000000000000;
	sram_mem[77047] = 16'b0000000000000000;
	sram_mem[77048] = 16'b0000000000000000;
	sram_mem[77049] = 16'b0000000000000000;
	sram_mem[77050] = 16'b0000000000000000;
	sram_mem[77051] = 16'b0000000000000000;
	sram_mem[77052] = 16'b0000000000000000;
	sram_mem[77053] = 16'b0000000000000000;
	sram_mem[77054] = 16'b0000000000000000;
	sram_mem[77055] = 16'b0000000000000000;
	sram_mem[77056] = 16'b0000000000000000;
	sram_mem[77057] = 16'b0000000000000000;
	sram_mem[77058] = 16'b0000000000000000;
	sram_mem[77059] = 16'b0000000000000000;
	sram_mem[77060] = 16'b0000000000000000;
	sram_mem[77061] = 16'b0000000000000000;
	sram_mem[77062] = 16'b0000000000000000;
	sram_mem[77063] = 16'b0000000000000000;
	sram_mem[77064] = 16'b0000000000000000;
	sram_mem[77065] = 16'b0000000000000000;
	sram_mem[77066] = 16'b0000000000000000;
	sram_mem[77067] = 16'b0000000000000000;
	sram_mem[77068] = 16'b0000000000000000;
	sram_mem[77069] = 16'b0000000000000000;
	sram_mem[77070] = 16'b0000000000000000;
	sram_mem[77071] = 16'b0000000000000000;
	sram_mem[77072] = 16'b0000000000000000;
	sram_mem[77073] = 16'b0000000000000000;
	sram_mem[77074] = 16'b0000000000000000;
	sram_mem[77075] = 16'b0000000000000000;
	sram_mem[77076] = 16'b0000000000000000;
	sram_mem[77077] = 16'b0000000000000000;
	sram_mem[77078] = 16'b0000000000000000;
	sram_mem[77079] = 16'b0000000000000000;
	sram_mem[77080] = 16'b0000000000000000;
	sram_mem[77081] = 16'b0000000000000000;
	sram_mem[77082] = 16'b0000000000000000;
	sram_mem[77083] = 16'b0000000000000000;
	sram_mem[77084] = 16'b0000000000000000;
	sram_mem[77085] = 16'b0000000000000000;
	sram_mem[77086] = 16'b0000000000000000;
	sram_mem[77087] = 16'b0000000000000000;
	sram_mem[77088] = 16'b0000000000000000;
	sram_mem[77089] = 16'b0000000000000000;
	sram_mem[77090] = 16'b0000000000000000;
	sram_mem[77091] = 16'b0000000000000000;
	sram_mem[77092] = 16'b0000000000000000;
	sram_mem[77093] = 16'b0000000000000000;
	sram_mem[77094] = 16'b0000000000000000;
	sram_mem[77095] = 16'b0000000000000000;
	sram_mem[77096] = 16'b0000000000000000;
	sram_mem[77097] = 16'b0000000000000000;
	sram_mem[77098] = 16'b0000000000000000;
	sram_mem[77099] = 16'b0000000000000000;
	sram_mem[77100] = 16'b0000000000000000;
	sram_mem[77101] = 16'b0000000000000000;
	sram_mem[77102] = 16'b0000000000000000;
	sram_mem[77103] = 16'b0000000000000000;
	sram_mem[77104] = 16'b0000000000000000;
	sram_mem[77105] = 16'b0000000000000000;
	sram_mem[77106] = 16'b0000000000000000;
	sram_mem[77107] = 16'b0000000000000000;
	sram_mem[77108] = 16'b0000000000000000;
	sram_mem[77109] = 16'b0000000000000000;
	sram_mem[77110] = 16'b0000000000000000;
	sram_mem[77111] = 16'b0000000000000000;
	sram_mem[77112] = 16'b0000000000000000;
	sram_mem[77113] = 16'b0000000000000000;
	sram_mem[77114] = 16'b0000000000000000;
	sram_mem[77115] = 16'b0000000000000000;
	sram_mem[77116] = 16'b0000000000000000;
	sram_mem[77117] = 16'b0000000000000000;
	sram_mem[77118] = 16'b0000000000000000;
	sram_mem[77119] = 16'b0000000000000000;
	sram_mem[77120] = 16'b0000000000000000;
	sram_mem[77121] = 16'b0000000000000000;
	sram_mem[77122] = 16'b0000000000000000;
	sram_mem[77123] = 16'b0000000000000000;
	sram_mem[77124] = 16'b0000000000000000;
	sram_mem[77125] = 16'b0000000000000000;
	sram_mem[77126] = 16'b0000000000000000;
	sram_mem[77127] = 16'b0000000000000000;
	sram_mem[77128] = 16'b0000000000000000;
	sram_mem[77129] = 16'b0000000000000000;
	sram_mem[77130] = 16'b0000000000000000;
	sram_mem[77131] = 16'b0000000000000000;
	sram_mem[77132] = 16'b0000000000000000;
	sram_mem[77133] = 16'b0000000000000000;
	sram_mem[77134] = 16'b0000000000000000;
	sram_mem[77135] = 16'b0000000000000000;
	sram_mem[77136] = 16'b0000000000000000;
	sram_mem[77137] = 16'b0000000000000000;
	sram_mem[77138] = 16'b0000000000000000;
	sram_mem[77139] = 16'b0000000000000000;
	sram_mem[77140] = 16'b0000000000000000;
	sram_mem[77141] = 16'b0000000000000000;
	sram_mem[77142] = 16'b0000000000000000;
	sram_mem[77143] = 16'b0000000000000000;
	sram_mem[77144] = 16'b0000000000000000;
	sram_mem[77145] = 16'b0000000000000000;
	sram_mem[77146] = 16'b0000000000000000;
	sram_mem[77147] = 16'b0000000000000000;
	sram_mem[77148] = 16'b0000000000000000;
	sram_mem[77149] = 16'b0000000000000000;
	sram_mem[77150] = 16'b0000000000000000;
	sram_mem[77151] = 16'b0000000000000000;
	sram_mem[77152] = 16'b0000000000000000;
	sram_mem[77153] = 16'b0000000000000000;
	sram_mem[77154] = 16'b0000000000000000;
	sram_mem[77155] = 16'b0000000000000000;
	sram_mem[77156] = 16'b0000000000000000;
	sram_mem[77157] = 16'b0000000000000000;
	sram_mem[77158] = 16'b0000000000000000;
	sram_mem[77159] = 16'b0000000000000000;
	sram_mem[77160] = 16'b0000000000000000;
	sram_mem[77161] = 16'b0000000000000000;
	sram_mem[77162] = 16'b0000000000000000;
	sram_mem[77163] = 16'b0000000000000000;
	sram_mem[77164] = 16'b0000000000000000;
	sram_mem[77165] = 16'b0000000000000000;
	sram_mem[77166] = 16'b0000000000000000;
	sram_mem[77167] = 16'b0000000000000000;
	sram_mem[77168] = 16'b0000000000000000;
	sram_mem[77169] = 16'b0000000000000000;
	sram_mem[77170] = 16'b0000000000000000;
	sram_mem[77171] = 16'b0000000000000000;
	sram_mem[77172] = 16'b0000000000000000;
	sram_mem[77173] = 16'b0000000000000000;
	sram_mem[77174] = 16'b0000000000000000;
	sram_mem[77175] = 16'b0000000000000000;
	sram_mem[77176] = 16'b0000000000000000;
	sram_mem[77177] = 16'b0000000000000000;
	sram_mem[77178] = 16'b0000000000000000;
	sram_mem[77179] = 16'b0000000000000000;
	sram_mem[77180] = 16'b0000000000000000;
	sram_mem[77181] = 16'b0000000000000000;
	sram_mem[77182] = 16'b0000000000000000;
	sram_mem[77183] = 16'b0000000000000000;
	sram_mem[77184] = 16'b0000000000000000;
	sram_mem[77185] = 16'b0000000000000000;
	sram_mem[77186] = 16'b0000000000000000;
	sram_mem[77187] = 16'b0000000000000000;
	sram_mem[77188] = 16'b0000000000000000;
	sram_mem[77189] = 16'b0000000000000000;
	sram_mem[77190] = 16'b0000000000000000;
	sram_mem[77191] = 16'b0000000000000000;
	sram_mem[77192] = 16'b0000000000000000;
	sram_mem[77193] = 16'b0000000000000000;
	sram_mem[77194] = 16'b0000000000000000;
	sram_mem[77195] = 16'b0000000000000000;
	sram_mem[77196] = 16'b0000000000000000;
	sram_mem[77197] = 16'b0000000000000000;
	sram_mem[77198] = 16'b0000000000000000;
	sram_mem[77199] = 16'b0000000000000000;
	sram_mem[77200] = 16'b0000000000000000;
	sram_mem[77201] = 16'b0000000000000000;
	sram_mem[77202] = 16'b0000000000000000;
	sram_mem[77203] = 16'b0000000000000000;
	sram_mem[77204] = 16'b0000000000000000;
	sram_mem[77205] = 16'b0000000000000000;
	sram_mem[77206] = 16'b0000000000000000;
	sram_mem[77207] = 16'b0000000000000000;
	sram_mem[77208] = 16'b0000000000000000;
	sram_mem[77209] = 16'b0000000000000000;
	sram_mem[77210] = 16'b0000000000000000;
	sram_mem[77211] = 16'b0000000000000000;
	sram_mem[77212] = 16'b0000000000000000;
	sram_mem[77213] = 16'b0000000000000000;
	sram_mem[77214] = 16'b0000000000000000;
	sram_mem[77215] = 16'b0000000000000000;
	sram_mem[77216] = 16'b0000000000000000;
	sram_mem[77217] = 16'b0000000000000000;
	sram_mem[77218] = 16'b0000000000000000;
	sram_mem[77219] = 16'b0000000000000000;
	sram_mem[77220] = 16'b0000000000000000;
	sram_mem[77221] = 16'b0000000000000000;
	sram_mem[77222] = 16'b0000000000000000;
	sram_mem[77223] = 16'b0000000000000000;
	sram_mem[77224] = 16'b0000000000000000;
	sram_mem[77225] = 16'b0000000000000000;
	sram_mem[77226] = 16'b0000000000000000;
	sram_mem[77227] = 16'b0000000000000000;
	sram_mem[77228] = 16'b0000000000000000;
	sram_mem[77229] = 16'b0000000000000000;
	sram_mem[77230] = 16'b0000000000000000;
	sram_mem[77231] = 16'b0000000000000000;
	sram_mem[77232] = 16'b0000000000000000;
	sram_mem[77233] = 16'b0000000000000000;
	sram_mem[77234] = 16'b0000000000000000;
	sram_mem[77235] = 16'b0000000000000000;
	sram_mem[77236] = 16'b0000000000000000;
	sram_mem[77237] = 16'b0000000000000000;
	sram_mem[77238] = 16'b0000000000000000;
	sram_mem[77239] = 16'b0000000000000000;
	sram_mem[77240] = 16'b0000000000000000;
	sram_mem[77241] = 16'b0000000000000000;
	sram_mem[77242] = 16'b0000000000000000;
	sram_mem[77243] = 16'b0000000000000000;
	sram_mem[77244] = 16'b0000000000000000;
	sram_mem[77245] = 16'b0000000000000000;
	sram_mem[77246] = 16'b0000000000000000;
	sram_mem[77247] = 16'b0000000000000000;
	sram_mem[77248] = 16'b0000000000000000;
	sram_mem[77249] = 16'b0000000000000000;
	sram_mem[77250] = 16'b0000000000000000;
	sram_mem[77251] = 16'b0000000000000000;
	sram_mem[77252] = 16'b0000000000000000;
	sram_mem[77253] = 16'b0000000000000000;
	sram_mem[77254] = 16'b0000000000000000;
	sram_mem[77255] = 16'b0000000000000000;
	sram_mem[77256] = 16'b0000000000000000;
	sram_mem[77257] = 16'b0000000000000000;
	sram_mem[77258] = 16'b0000000000000000;
	sram_mem[77259] = 16'b0000000000000000;
	sram_mem[77260] = 16'b0000000000000000;
	sram_mem[77261] = 16'b0000000000000000;
	sram_mem[77262] = 16'b0000000000000000;
	sram_mem[77263] = 16'b0000000000000000;
	sram_mem[77264] = 16'b0000000000000000;
	sram_mem[77265] = 16'b0000000000000000;
	sram_mem[77266] = 16'b0000000000000000;
	sram_mem[77267] = 16'b0000000000000000;
	sram_mem[77268] = 16'b0000000000000000;
	sram_mem[77269] = 16'b0000000000000000;
	sram_mem[77270] = 16'b0000000000000000;
	sram_mem[77271] = 16'b0000000000000000;
	sram_mem[77272] = 16'b0000000000000000;
	sram_mem[77273] = 16'b0000000000000000;
	sram_mem[77274] = 16'b0000000000000000;
	sram_mem[77275] = 16'b0000000000000000;
	sram_mem[77276] = 16'b0000000000000000;
	sram_mem[77277] = 16'b0000000000000000;
	sram_mem[77278] = 16'b0000000000000000;
	sram_mem[77279] = 16'b0000000000000000;
	sram_mem[77280] = 16'b0000000000000000;
	sram_mem[77281] = 16'b0000000000000000;
	sram_mem[77282] = 16'b0000000000000000;
	sram_mem[77283] = 16'b0000000000000000;
	sram_mem[77284] = 16'b0000000000000000;
	sram_mem[77285] = 16'b0000000000000000;
	sram_mem[77286] = 16'b0000000000000000;
	sram_mem[77287] = 16'b0000000000000000;
	sram_mem[77288] = 16'b0000000000000000;
	sram_mem[77289] = 16'b0000000000000000;
	sram_mem[77290] = 16'b0000000000000000;
	sram_mem[77291] = 16'b0000000000000000;
	sram_mem[77292] = 16'b0000000000000000;
	sram_mem[77293] = 16'b0000000000000000;
	sram_mem[77294] = 16'b0000000000000000;
	sram_mem[77295] = 16'b0000000000000000;
	sram_mem[77296] = 16'b0000000000000000;
	sram_mem[77297] = 16'b0000000000000000;
	sram_mem[77298] = 16'b0000000000000000;
	sram_mem[77299] = 16'b0000000000000000;
	sram_mem[77300] = 16'b0000000000000000;
	sram_mem[77301] = 16'b0000000000000000;
	sram_mem[77302] = 16'b0000000000000000;
	sram_mem[77303] = 16'b0000000000000000;
	sram_mem[77304] = 16'b0000000000000000;
	sram_mem[77305] = 16'b0000000000000000;
	sram_mem[77306] = 16'b0000000000000000;
	sram_mem[77307] = 16'b0000000000000000;
	sram_mem[77308] = 16'b0000000000000000;
	sram_mem[77309] = 16'b0000000000000000;
	sram_mem[77310] = 16'b0000000000000000;
	sram_mem[77311] = 16'b0000000000000000;
	sram_mem[77312] = 16'b0000000000000000;
	sram_mem[77313] = 16'b0000000000000000;
	sram_mem[77314] = 16'b0000000000000000;
	sram_mem[77315] = 16'b0000000000000000;
	sram_mem[77316] = 16'b0000000000000000;
	sram_mem[77317] = 16'b0000000000000000;
	sram_mem[77318] = 16'b0000000000000000;
	sram_mem[77319] = 16'b0000000000000000;
	sram_mem[77320] = 16'b0000000000000000;
	sram_mem[77321] = 16'b0000000000000000;
	sram_mem[77322] = 16'b0000000000000000;
	sram_mem[77323] = 16'b0000000000000000;
	sram_mem[77324] = 16'b0000000000000000;
	sram_mem[77325] = 16'b0000000000000000;
	sram_mem[77326] = 16'b0000000000000000;
	sram_mem[77327] = 16'b0000000000000000;
	sram_mem[77328] = 16'b0000000000000000;
	sram_mem[77329] = 16'b0000000000000000;
	sram_mem[77330] = 16'b0000000000000000;
	sram_mem[77331] = 16'b0000000000000000;
	sram_mem[77332] = 16'b0000000000000000;
	sram_mem[77333] = 16'b0000000000000000;
	sram_mem[77334] = 16'b0000000000000000;
	sram_mem[77335] = 16'b0000000000000000;
	sram_mem[77336] = 16'b0000000000000000;
	sram_mem[77337] = 16'b0000000000000000;
	sram_mem[77338] = 16'b0000000000000000;
	sram_mem[77339] = 16'b0000000000000000;
	sram_mem[77340] = 16'b0000000000000000;
	sram_mem[77341] = 16'b0000000000000000;
	sram_mem[77342] = 16'b0000000000000000;
	sram_mem[77343] = 16'b0000000000000000;
	sram_mem[77344] = 16'b0000000000000000;
	sram_mem[77345] = 16'b0000000000000000;
	sram_mem[77346] = 16'b0000000000000000;
	sram_mem[77347] = 16'b0000000000000000;
	sram_mem[77348] = 16'b0000000000000000;
	sram_mem[77349] = 16'b0000000000000000;
	sram_mem[77350] = 16'b0000000000000000;
	sram_mem[77351] = 16'b0000000000000000;
	sram_mem[77352] = 16'b0000000000000000;
	sram_mem[77353] = 16'b0000000000000000;
	sram_mem[77354] = 16'b0000000000000000;
	sram_mem[77355] = 16'b0000000000000000;
	sram_mem[77356] = 16'b0000000000000000;
	sram_mem[77357] = 16'b0000000000000000;
	sram_mem[77358] = 16'b0000000000000000;
	sram_mem[77359] = 16'b0000000000000000;
	sram_mem[77360] = 16'b0000000000000000;
	sram_mem[77361] = 16'b0000000000000000;
	sram_mem[77362] = 16'b0000000000000000;
	sram_mem[77363] = 16'b0000000000000000;
	sram_mem[77364] = 16'b0000000000000000;
	sram_mem[77365] = 16'b0000000000000000;
	sram_mem[77366] = 16'b0000000000000000;
	sram_mem[77367] = 16'b0000000000000000;
	sram_mem[77368] = 16'b0000000000000000;
	sram_mem[77369] = 16'b0000000000000000;
	sram_mem[77370] = 16'b0000000000000000;
	sram_mem[77371] = 16'b0000000000000000;
	sram_mem[77372] = 16'b0000000000000000;
	sram_mem[77373] = 16'b0000000000000000;
	sram_mem[77374] = 16'b0000000000000000;
	sram_mem[77375] = 16'b0000000000000000;
	sram_mem[77376] = 16'b0000000000000000;
	sram_mem[77377] = 16'b0000000000000000;
	sram_mem[77378] = 16'b0000000000000000;
	sram_mem[77379] = 16'b0000000000000000;
	sram_mem[77380] = 16'b0000000000000000;
	sram_mem[77381] = 16'b0000000000000000;
	sram_mem[77382] = 16'b0000000000000000;
	sram_mem[77383] = 16'b0000000000000000;
	sram_mem[77384] = 16'b0000000000000000;
	sram_mem[77385] = 16'b0000000000000000;
	sram_mem[77386] = 16'b0000000000000000;
	sram_mem[77387] = 16'b0000000000000000;
	sram_mem[77388] = 16'b0000000000000000;
	sram_mem[77389] = 16'b0000000000000000;
	sram_mem[77390] = 16'b0000000000000000;
	sram_mem[77391] = 16'b0000000000000000;
	sram_mem[77392] = 16'b0000000000000000;
	sram_mem[77393] = 16'b0000000000000000;
	sram_mem[77394] = 16'b0000000000000000;
	sram_mem[77395] = 16'b0000000000000000;
	sram_mem[77396] = 16'b0000000000000000;
	sram_mem[77397] = 16'b0000000000000000;
	sram_mem[77398] = 16'b0000000000000000;
	sram_mem[77399] = 16'b0000000000000000;
	sram_mem[77400] = 16'b0000000000000000;
	sram_mem[77401] = 16'b0000000000000000;
	sram_mem[77402] = 16'b0000000000000000;
	sram_mem[77403] = 16'b0000000000000000;
	sram_mem[77404] = 16'b0000000000000000;
	sram_mem[77405] = 16'b0000000000000000;
	sram_mem[77406] = 16'b0000000000000000;
	sram_mem[77407] = 16'b0000000000000000;
	sram_mem[77408] = 16'b0000000000000000;
	sram_mem[77409] = 16'b0000000000000000;
	sram_mem[77410] = 16'b0000000000000000;
	sram_mem[77411] = 16'b0000000000000000;
	sram_mem[77412] = 16'b0000000000000000;
	sram_mem[77413] = 16'b0000000000000000;
	sram_mem[77414] = 16'b0000000000000000;
	sram_mem[77415] = 16'b0000000000000000;
	sram_mem[77416] = 16'b0000000000000000;
	sram_mem[77417] = 16'b0000000000000000;
	sram_mem[77418] = 16'b0000000000000000;
	sram_mem[77419] = 16'b0000000000000000;
	sram_mem[77420] = 16'b0000000000000000;
	sram_mem[77421] = 16'b0000000000000000;
	sram_mem[77422] = 16'b0000000000000000;
	sram_mem[77423] = 16'b0000000000000000;
	sram_mem[77424] = 16'b0000000000000000;
	sram_mem[77425] = 16'b0000000000000000;
	sram_mem[77426] = 16'b0000000000000000;
	sram_mem[77427] = 16'b0000000000000000;
	sram_mem[77428] = 16'b0000000000000000;
	sram_mem[77429] = 16'b0000000000000000;
	sram_mem[77430] = 16'b0000000000000000;
	sram_mem[77431] = 16'b0000000000000000;
	sram_mem[77432] = 16'b0000000000000000;
	sram_mem[77433] = 16'b0000000000000000;
	sram_mem[77434] = 16'b0000000000000000;
	sram_mem[77435] = 16'b0000000000000000;
	sram_mem[77436] = 16'b0000000000000000;
	sram_mem[77437] = 16'b0000000000000000;
	sram_mem[77438] = 16'b0000000000000000;
	sram_mem[77439] = 16'b0000000000000000;
	sram_mem[77440] = 16'b0000000000000000;
	sram_mem[77441] = 16'b0000000000000000;
	sram_mem[77442] = 16'b0000000000000000;
	sram_mem[77443] = 16'b0000000000000000;
	sram_mem[77444] = 16'b0000000000000000;
	sram_mem[77445] = 16'b0000000000000000;
	sram_mem[77446] = 16'b0000000000000000;
	sram_mem[77447] = 16'b0000000000000000;
	sram_mem[77448] = 16'b0000000000000000;
	sram_mem[77449] = 16'b0000000000000000;
	sram_mem[77450] = 16'b0000000000000000;
	sram_mem[77451] = 16'b0000000000000000;
	sram_mem[77452] = 16'b0000000000000000;
	sram_mem[77453] = 16'b0000000000000000;
	sram_mem[77454] = 16'b0000000000000000;
	sram_mem[77455] = 16'b0000000000000000;
	sram_mem[77456] = 16'b0000000000000000;
	sram_mem[77457] = 16'b0000000000000000;
	sram_mem[77458] = 16'b0000000000000000;
	sram_mem[77459] = 16'b0000000000000000;
	sram_mem[77460] = 16'b0000000000000000;
	sram_mem[77461] = 16'b0000000000000000;
	sram_mem[77462] = 16'b0000000000000000;
	sram_mem[77463] = 16'b0000000000000000;
	sram_mem[77464] = 16'b0000000000000000;
	sram_mem[77465] = 16'b0000000000000000;
	sram_mem[77466] = 16'b0000000000000000;
	sram_mem[77467] = 16'b0000000000000000;
	sram_mem[77468] = 16'b0000000000000000;
	sram_mem[77469] = 16'b0000000000000000;
	sram_mem[77470] = 16'b0000000000000000;
	sram_mem[77471] = 16'b0000000000000000;
	sram_mem[77472] = 16'b0000000000000000;
	sram_mem[77473] = 16'b0000000000000000;
	sram_mem[77474] = 16'b0000000000000000;
	sram_mem[77475] = 16'b0000000000000000;
	sram_mem[77476] = 16'b0000000000000000;
	sram_mem[77477] = 16'b0000000000000000;
	sram_mem[77478] = 16'b0000000000000000;
	sram_mem[77479] = 16'b0000000000000000;
	sram_mem[77480] = 16'b0000000000000000;
	sram_mem[77481] = 16'b0000000000000000;
	sram_mem[77482] = 16'b0000000000000000;
	sram_mem[77483] = 16'b0000000000000000;
	sram_mem[77484] = 16'b0000000000000000;
	sram_mem[77485] = 16'b0000000000000000;
	sram_mem[77486] = 16'b0000000000000000;
	sram_mem[77487] = 16'b0000000000000000;
	sram_mem[77488] = 16'b0000000000000000;
	sram_mem[77489] = 16'b0000000000000000;
	sram_mem[77490] = 16'b0000000000000000;
	sram_mem[77491] = 16'b0000000000000000;
	sram_mem[77492] = 16'b0000000000000000;
	sram_mem[77493] = 16'b0000000000000000;
	sram_mem[77494] = 16'b0000000000000000;
	sram_mem[77495] = 16'b0000000000000000;
	sram_mem[77496] = 16'b0000000000000000;
	sram_mem[77497] = 16'b0000000000000000;
	sram_mem[77498] = 16'b0000000000000000;
	sram_mem[77499] = 16'b0000000000000000;
	sram_mem[77500] = 16'b0000000000000000;
	sram_mem[77501] = 16'b0000000000000000;
	sram_mem[77502] = 16'b0000000000000000;
	sram_mem[77503] = 16'b0000000000000000;
	sram_mem[77504] = 16'b0000000000000000;
	sram_mem[77505] = 16'b0000000000000000;
	sram_mem[77506] = 16'b0000000000000000;
	sram_mem[77507] = 16'b0000000000000000;
	sram_mem[77508] = 16'b0000000000000000;
	sram_mem[77509] = 16'b0000000000000000;
	sram_mem[77510] = 16'b0000000000000000;
	sram_mem[77511] = 16'b0000000000000000;
	sram_mem[77512] = 16'b0000000000000000;
	sram_mem[77513] = 16'b0000000000000000;
	sram_mem[77514] = 16'b0000000000000000;
	sram_mem[77515] = 16'b0000000000000000;
	sram_mem[77516] = 16'b0000000000000000;
	sram_mem[77517] = 16'b0000000000000000;
	sram_mem[77518] = 16'b0000000000000000;
	sram_mem[77519] = 16'b0000000000000000;
	sram_mem[77520] = 16'b0000000000000000;
	sram_mem[77521] = 16'b0000000000000000;
	sram_mem[77522] = 16'b0000000000000000;
	sram_mem[77523] = 16'b0000000000000000;
	sram_mem[77524] = 16'b0000000000000000;
	sram_mem[77525] = 16'b0000000000000000;
	sram_mem[77526] = 16'b0000000000000000;
	sram_mem[77527] = 16'b0000000000000000;
	sram_mem[77528] = 16'b0000000000000000;
	sram_mem[77529] = 16'b0000000000000000;
	sram_mem[77530] = 16'b0000000000000000;
	sram_mem[77531] = 16'b0000000000000000;
	sram_mem[77532] = 16'b0000000000000000;
	sram_mem[77533] = 16'b0000000000000000;
	sram_mem[77534] = 16'b0000000000000000;
	sram_mem[77535] = 16'b0000000000000000;
	sram_mem[77536] = 16'b0000000000000000;
	sram_mem[77537] = 16'b0000000000000000;
	sram_mem[77538] = 16'b0000000000000000;
	sram_mem[77539] = 16'b0000000000000000;
	sram_mem[77540] = 16'b0000000000000000;
	sram_mem[77541] = 16'b0000000000000000;
	sram_mem[77542] = 16'b0000000000000000;
	sram_mem[77543] = 16'b0000000000000000;
	sram_mem[77544] = 16'b0000000000000000;
	sram_mem[77545] = 16'b0000000000000000;
	sram_mem[77546] = 16'b0000000000000000;
	sram_mem[77547] = 16'b0000000000000000;
	sram_mem[77548] = 16'b0000000000000000;
	sram_mem[77549] = 16'b0000000000000000;
	sram_mem[77550] = 16'b0000000000000000;
	sram_mem[77551] = 16'b0000000000000000;
	sram_mem[77552] = 16'b0000000000000000;
	sram_mem[77553] = 16'b0000000000000000;
	sram_mem[77554] = 16'b0000000000000000;
	sram_mem[77555] = 16'b0000000000000000;
	sram_mem[77556] = 16'b0000000000000000;
	sram_mem[77557] = 16'b0000000000000000;
	sram_mem[77558] = 16'b0000000000000000;
	sram_mem[77559] = 16'b0000000000000000;
	sram_mem[77560] = 16'b0000000000000000;
	sram_mem[77561] = 16'b0000000000000000;
	sram_mem[77562] = 16'b0000000000000000;
	sram_mem[77563] = 16'b0000000000000000;
	sram_mem[77564] = 16'b0000000000000000;
	sram_mem[77565] = 16'b0000000000000000;
	sram_mem[77566] = 16'b0000000000000000;
	sram_mem[77567] = 16'b0000000000000000;
	sram_mem[77568] = 16'b0000000000000000;
	sram_mem[77569] = 16'b0000000000000000;
	sram_mem[77570] = 16'b0000000000000000;
	sram_mem[77571] = 16'b0000000000000000;
	sram_mem[77572] = 16'b0000000000000000;
	sram_mem[77573] = 16'b0000000000000000;
	sram_mem[77574] = 16'b0000000000000000;
	sram_mem[77575] = 16'b0000000000000000;
	sram_mem[77576] = 16'b0000000000000000;
	sram_mem[77577] = 16'b0000000000000000;
	sram_mem[77578] = 16'b0000000000000000;
	sram_mem[77579] = 16'b0000000000000000;
	sram_mem[77580] = 16'b0000000000000000;
	sram_mem[77581] = 16'b0000000000000000;
	sram_mem[77582] = 16'b0000000000000000;
	sram_mem[77583] = 16'b0000000000000000;
	sram_mem[77584] = 16'b0000000000000000;
	sram_mem[77585] = 16'b0000000000000000;
	sram_mem[77586] = 16'b0000000000000000;
	sram_mem[77587] = 16'b0000000000000000;
	sram_mem[77588] = 16'b0000000000000000;
	sram_mem[77589] = 16'b0000000000000000;
	sram_mem[77590] = 16'b0000000000000000;
	sram_mem[77591] = 16'b0000000000000000;
	sram_mem[77592] = 16'b0000000000000000;
	sram_mem[77593] = 16'b0000000000000000;
	sram_mem[77594] = 16'b0000000000000000;
	sram_mem[77595] = 16'b0000000000000000;
	sram_mem[77596] = 16'b0000000000000000;
	sram_mem[77597] = 16'b0000000000000000;
	sram_mem[77598] = 16'b0000000000000000;
	sram_mem[77599] = 16'b0000000000000000;
	sram_mem[77600] = 16'b0000000000000000;
	sram_mem[77601] = 16'b0000000000000000;
	sram_mem[77602] = 16'b0000000000000000;
	sram_mem[77603] = 16'b0000000000000000;
	sram_mem[77604] = 16'b0000000000000000;
	sram_mem[77605] = 16'b0000000000000000;
	sram_mem[77606] = 16'b0000000000000000;
	sram_mem[77607] = 16'b0000000000000000;
	sram_mem[77608] = 16'b0000000000000000;
	sram_mem[77609] = 16'b0000000000000000;
	sram_mem[77610] = 16'b0000000000000000;
	sram_mem[77611] = 16'b0000000000000000;
	sram_mem[77612] = 16'b0000000000000000;
	sram_mem[77613] = 16'b0000000000000000;
	sram_mem[77614] = 16'b0000000000000000;
	sram_mem[77615] = 16'b0000000000000000;
	sram_mem[77616] = 16'b0000000000000000;
	sram_mem[77617] = 16'b0000000000000000;
	sram_mem[77618] = 16'b0000000000000000;
	sram_mem[77619] = 16'b0000000000000000;
	sram_mem[77620] = 16'b0000000000000000;
	sram_mem[77621] = 16'b0000000000000000;
	sram_mem[77622] = 16'b0000000000000000;
	sram_mem[77623] = 16'b0000000000000000;
	sram_mem[77624] = 16'b0000000000000000;
	sram_mem[77625] = 16'b0000000000000000;
	sram_mem[77626] = 16'b0000000000000000;
	sram_mem[77627] = 16'b0000000000000000;
	sram_mem[77628] = 16'b0000000000000000;
	sram_mem[77629] = 16'b0000000000000000;
	sram_mem[77630] = 16'b0000000000000000;
	sram_mem[77631] = 16'b0000000000000000;
	sram_mem[77632] = 16'b0000000000000000;
	sram_mem[77633] = 16'b0000000000000000;
	sram_mem[77634] = 16'b0000000000000000;
	sram_mem[77635] = 16'b0000000000000000;
	sram_mem[77636] = 16'b0000000000000000;
	sram_mem[77637] = 16'b0000000000000000;
	sram_mem[77638] = 16'b0000000000000000;
	sram_mem[77639] = 16'b0000000000000000;
	sram_mem[77640] = 16'b0000000000000000;
	sram_mem[77641] = 16'b0000000000000000;
	sram_mem[77642] = 16'b0000000000000000;
	sram_mem[77643] = 16'b0000000000000000;
	sram_mem[77644] = 16'b0000000000000000;
	sram_mem[77645] = 16'b0000000000000000;
	sram_mem[77646] = 16'b0000000000000000;
	sram_mem[77647] = 16'b0000000000000000;
	sram_mem[77648] = 16'b0000000000000000;
	sram_mem[77649] = 16'b0000000000000000;
	sram_mem[77650] = 16'b0000000000000000;
	sram_mem[77651] = 16'b0000000000000000;
	sram_mem[77652] = 16'b0000000000000000;
	sram_mem[77653] = 16'b0000000000000000;
	sram_mem[77654] = 16'b0000000000000000;
	sram_mem[77655] = 16'b0000000000000000;
	sram_mem[77656] = 16'b0000000000000000;
	sram_mem[77657] = 16'b0000000000000000;
	sram_mem[77658] = 16'b0000000000000000;
	sram_mem[77659] = 16'b0000000000000000;
	sram_mem[77660] = 16'b0000000000000000;
	sram_mem[77661] = 16'b0000000000000000;
	sram_mem[77662] = 16'b0000000000000000;
	sram_mem[77663] = 16'b0000000000000000;
	sram_mem[77664] = 16'b0000000000000000;
	sram_mem[77665] = 16'b0000000000000000;
	sram_mem[77666] = 16'b0000000000000000;
	sram_mem[77667] = 16'b0000000000000000;
	sram_mem[77668] = 16'b0000000000000000;
	sram_mem[77669] = 16'b0000000000000000;
	sram_mem[77670] = 16'b0000000000000000;
	sram_mem[77671] = 16'b0000000000000000;
	sram_mem[77672] = 16'b0000000000000000;
	sram_mem[77673] = 16'b0000000000000000;
	sram_mem[77674] = 16'b0000000000000000;
	sram_mem[77675] = 16'b0000000000000000;
	sram_mem[77676] = 16'b0000000000000000;
	sram_mem[77677] = 16'b0000000000000000;
	sram_mem[77678] = 16'b0000000000000000;
	sram_mem[77679] = 16'b0000000000000000;
	sram_mem[77680] = 16'b0000000000000000;
	sram_mem[77681] = 16'b0000000000000000;
	sram_mem[77682] = 16'b0000000000000000;
	sram_mem[77683] = 16'b0000000000000000;
	sram_mem[77684] = 16'b0000000000000000;
	sram_mem[77685] = 16'b0000000000000000;
	sram_mem[77686] = 16'b0000000000000000;
	sram_mem[77687] = 16'b0000000000000000;
	sram_mem[77688] = 16'b0000000000000000;
	sram_mem[77689] = 16'b0000000000000000;
	sram_mem[77690] = 16'b0000000000000000;
	sram_mem[77691] = 16'b0000000000000000;
	sram_mem[77692] = 16'b0000000000000000;
	sram_mem[77693] = 16'b0000000000000000;
	sram_mem[77694] = 16'b0000000000000000;
	sram_mem[77695] = 16'b0000000000000000;
	sram_mem[77696] = 16'b0000000000000000;
	sram_mem[77697] = 16'b0000000000000000;
	sram_mem[77698] = 16'b0000000000000000;
	sram_mem[77699] = 16'b0000000000000000;
	sram_mem[77700] = 16'b0000000000000000;
	sram_mem[77701] = 16'b0000000000000000;
	sram_mem[77702] = 16'b0000000000000000;
	sram_mem[77703] = 16'b0000000000000000;
	sram_mem[77704] = 16'b0000000000000000;
	sram_mem[77705] = 16'b0000000000000000;
	sram_mem[77706] = 16'b0000000000000000;
	sram_mem[77707] = 16'b0000000000000000;
	sram_mem[77708] = 16'b0000000000000000;
	sram_mem[77709] = 16'b0000000000000000;
	sram_mem[77710] = 16'b0000000000000000;
	sram_mem[77711] = 16'b0000000000000000;
	sram_mem[77712] = 16'b0000000000000000;
	sram_mem[77713] = 16'b0000000000000000;
	sram_mem[77714] = 16'b0000000000000000;
	sram_mem[77715] = 16'b0000000000000000;
	sram_mem[77716] = 16'b0000000000000000;
	sram_mem[77717] = 16'b0000000000000000;
	sram_mem[77718] = 16'b0000000000000000;
	sram_mem[77719] = 16'b0000000000000000;
	sram_mem[77720] = 16'b0000000000000000;
	sram_mem[77721] = 16'b0000000000000000;
	sram_mem[77722] = 16'b0000000000000000;
	sram_mem[77723] = 16'b0000000000000000;
	sram_mem[77724] = 16'b0000000000000000;
	sram_mem[77725] = 16'b0000000000000000;
	sram_mem[77726] = 16'b0000000000000000;
	sram_mem[77727] = 16'b0000000000000000;
	sram_mem[77728] = 16'b0000000000000000;
	sram_mem[77729] = 16'b0000000000000000;
	sram_mem[77730] = 16'b0000000000000000;
	sram_mem[77731] = 16'b0000000000000000;
	sram_mem[77732] = 16'b0000000000000000;
	sram_mem[77733] = 16'b0000000000000000;
	sram_mem[77734] = 16'b0000000000000000;
	sram_mem[77735] = 16'b0000000000000000;
	sram_mem[77736] = 16'b0000000000000000;
	sram_mem[77737] = 16'b0000000000000000;
	sram_mem[77738] = 16'b0000000000000000;
	sram_mem[77739] = 16'b0000000000000000;
	sram_mem[77740] = 16'b0000000000000000;
	sram_mem[77741] = 16'b0000000000000000;
	sram_mem[77742] = 16'b0000000000000000;
	sram_mem[77743] = 16'b0000000000000000;
	sram_mem[77744] = 16'b0000000000000000;
	sram_mem[77745] = 16'b0000000000000000;
	sram_mem[77746] = 16'b0000000000000000;
	sram_mem[77747] = 16'b0000000000000000;
	sram_mem[77748] = 16'b0000000000000000;
	sram_mem[77749] = 16'b0000000000000000;
	sram_mem[77750] = 16'b0000000000000000;
	sram_mem[77751] = 16'b0000000000000000;
	sram_mem[77752] = 16'b0000000000000000;
	sram_mem[77753] = 16'b0000000000000000;
	sram_mem[77754] = 16'b0000000000000000;
	sram_mem[77755] = 16'b0000000000000000;
	sram_mem[77756] = 16'b0000000000000000;
	sram_mem[77757] = 16'b0000000000000000;
	sram_mem[77758] = 16'b0000000000000000;
	sram_mem[77759] = 16'b0000000000000000;
	sram_mem[77760] = 16'b0000000000000000;
	sram_mem[77761] = 16'b0000000000000000;
	sram_mem[77762] = 16'b0000000000000000;
	sram_mem[77763] = 16'b0000000000000000;
	sram_mem[77764] = 16'b0000000000000000;
	sram_mem[77765] = 16'b0000000000000000;
	sram_mem[77766] = 16'b0000000000000000;
	sram_mem[77767] = 16'b0000000000000000;
	sram_mem[77768] = 16'b0000000000000000;
	sram_mem[77769] = 16'b0000000000000000;
	sram_mem[77770] = 16'b0000000000000000;
	sram_mem[77771] = 16'b0000000000000000;
	sram_mem[77772] = 16'b0000000000000000;
	sram_mem[77773] = 16'b0000000000000000;
	sram_mem[77774] = 16'b0000000000000000;
	sram_mem[77775] = 16'b0000000000000000;
	sram_mem[77776] = 16'b0000000000000000;
	sram_mem[77777] = 16'b0000000000000000;
	sram_mem[77778] = 16'b0000000000000000;
	sram_mem[77779] = 16'b0000000000000000;
	sram_mem[77780] = 16'b0000000000000000;
	sram_mem[77781] = 16'b0000000000000000;
	sram_mem[77782] = 16'b0000000000000000;
	sram_mem[77783] = 16'b0000000000000000;
	sram_mem[77784] = 16'b0000000000000000;
	sram_mem[77785] = 16'b0000000000000000;
	sram_mem[77786] = 16'b0000000000000000;
	sram_mem[77787] = 16'b0000000000000000;
	sram_mem[77788] = 16'b0000000000000000;
	sram_mem[77789] = 16'b0000000000000000;
	sram_mem[77790] = 16'b0000000000000000;
	sram_mem[77791] = 16'b0000000000000000;
	sram_mem[77792] = 16'b0000000000000000;
	sram_mem[77793] = 16'b0000000000000000;
	sram_mem[77794] = 16'b0000000000000000;
	sram_mem[77795] = 16'b0000000000000000;
	sram_mem[77796] = 16'b0000000000000000;
	sram_mem[77797] = 16'b0000000000000000;
	sram_mem[77798] = 16'b0000000000000000;
	sram_mem[77799] = 16'b0000000000000000;
	sram_mem[77800] = 16'b0000000000000000;
	sram_mem[77801] = 16'b0000000000000000;
	sram_mem[77802] = 16'b0000000000000000;
	sram_mem[77803] = 16'b0000000000000000;
	sram_mem[77804] = 16'b0000000000000000;
	sram_mem[77805] = 16'b0000000000000000;
	sram_mem[77806] = 16'b0000000000000000;
	sram_mem[77807] = 16'b0000000000000000;
	sram_mem[77808] = 16'b0000000000000000;
	sram_mem[77809] = 16'b0000000000000000;
	sram_mem[77810] = 16'b0000000000000000;
	sram_mem[77811] = 16'b0000000000000000;
	sram_mem[77812] = 16'b0000000000000000;
	sram_mem[77813] = 16'b0000000000000000;
	sram_mem[77814] = 16'b0000000000000000;
	sram_mem[77815] = 16'b0000000000000000;
	sram_mem[77816] = 16'b0000000000000000;
	sram_mem[77817] = 16'b0000000000000000;
	sram_mem[77818] = 16'b0000000000000000;
	sram_mem[77819] = 16'b0000000000000000;
	sram_mem[77820] = 16'b0000000000000000;
	sram_mem[77821] = 16'b0000000000000000;
	sram_mem[77822] = 16'b0000000000000000;
	sram_mem[77823] = 16'b0000000000000000;
	sram_mem[77824] = 16'b0000000000000000;
	sram_mem[77825] = 16'b0000000000000000;
	sram_mem[77826] = 16'b0000000000000000;
	sram_mem[77827] = 16'b0000000000000000;
	sram_mem[77828] = 16'b0000000000000000;
	sram_mem[77829] = 16'b0000000000000000;
	sram_mem[77830] = 16'b0000000000000000;
	sram_mem[77831] = 16'b0000000000000000;
	sram_mem[77832] = 16'b0000000000000000;
	sram_mem[77833] = 16'b0000000000000000;
	sram_mem[77834] = 16'b0000000000000000;
	sram_mem[77835] = 16'b0000000000000000;
	sram_mem[77836] = 16'b0000000000000000;
	sram_mem[77837] = 16'b0000000000000000;
	sram_mem[77838] = 16'b0000000000000000;
	sram_mem[77839] = 16'b0000000000000000;
	sram_mem[77840] = 16'b0000000000000000;
	sram_mem[77841] = 16'b0000000000000000;
	sram_mem[77842] = 16'b0000000000000000;
	sram_mem[77843] = 16'b0000000000000000;
	sram_mem[77844] = 16'b0000000000000000;
	sram_mem[77845] = 16'b0000000000000000;
	sram_mem[77846] = 16'b0000000000000000;
	sram_mem[77847] = 16'b0000000000000000;
	sram_mem[77848] = 16'b0000000000000000;
	sram_mem[77849] = 16'b0000000000000000;
	sram_mem[77850] = 16'b0000000000000000;
	sram_mem[77851] = 16'b0000000000000000;
	sram_mem[77852] = 16'b0000000000000000;
	sram_mem[77853] = 16'b0000000000000000;
	sram_mem[77854] = 16'b0000000000000000;
	sram_mem[77855] = 16'b0000000000000000;
	sram_mem[77856] = 16'b0000000000000000;
	sram_mem[77857] = 16'b0000000000000000;
	sram_mem[77858] = 16'b0000000000000000;
	sram_mem[77859] = 16'b0000000000000000;
	sram_mem[77860] = 16'b0000000000000000;
	sram_mem[77861] = 16'b0000000000000000;
	sram_mem[77862] = 16'b0000000000000000;
	sram_mem[77863] = 16'b0000000000000000;
	sram_mem[77864] = 16'b0000000000000000;
	sram_mem[77865] = 16'b0000000000000000;
	sram_mem[77866] = 16'b0000000000000000;
	sram_mem[77867] = 16'b0000000000000000;
	sram_mem[77868] = 16'b0000000000000000;
	sram_mem[77869] = 16'b0000000000000000;
	sram_mem[77870] = 16'b0000000000000000;
	sram_mem[77871] = 16'b0000000000000000;
	sram_mem[77872] = 16'b0000000000000000;
	sram_mem[77873] = 16'b0000000000000000;
	sram_mem[77874] = 16'b0000000000000000;
	sram_mem[77875] = 16'b0000000000000000;
	sram_mem[77876] = 16'b0000000000000000;
	sram_mem[77877] = 16'b0000000000000000;
	sram_mem[77878] = 16'b0000000000000000;
	sram_mem[77879] = 16'b0000000000000000;
	sram_mem[77880] = 16'b0000000000000000;
	sram_mem[77881] = 16'b0000000000000000;
	sram_mem[77882] = 16'b0000000000000000;
	sram_mem[77883] = 16'b0000000000000000;
	sram_mem[77884] = 16'b0000000000000000;
	sram_mem[77885] = 16'b0000000000000000;
	sram_mem[77886] = 16'b0000000000000000;
	sram_mem[77887] = 16'b0000000000000000;
	sram_mem[77888] = 16'b0000000000000000;
	sram_mem[77889] = 16'b0000000000000000;
	sram_mem[77890] = 16'b0000000000000000;
	sram_mem[77891] = 16'b0000000000000000;
	sram_mem[77892] = 16'b0000000000000000;
	sram_mem[77893] = 16'b0000000000000000;
	sram_mem[77894] = 16'b0000000000000000;
	sram_mem[77895] = 16'b0000000000000000;
	sram_mem[77896] = 16'b0000000000000000;
	sram_mem[77897] = 16'b0000000000000000;
	sram_mem[77898] = 16'b0000000000000000;
	sram_mem[77899] = 16'b0000000000000000;
	sram_mem[77900] = 16'b0000000000000000;
	sram_mem[77901] = 16'b0000000000000000;
	sram_mem[77902] = 16'b0000000000000000;
	sram_mem[77903] = 16'b0000000000000000;
	sram_mem[77904] = 16'b0000000000000000;
	sram_mem[77905] = 16'b0000000000000000;
	sram_mem[77906] = 16'b0000000000000000;
	sram_mem[77907] = 16'b0000000000000000;
	sram_mem[77908] = 16'b0000000000000000;
	sram_mem[77909] = 16'b0000000000000000;
	sram_mem[77910] = 16'b0000000000000000;
	sram_mem[77911] = 16'b0000000000000000;
	sram_mem[77912] = 16'b0000000000000000;
	sram_mem[77913] = 16'b0000000000000000;
	sram_mem[77914] = 16'b0000000000000000;
	sram_mem[77915] = 16'b0000000000000000;
	sram_mem[77916] = 16'b0000000000000000;
	sram_mem[77917] = 16'b0000000000000000;
	sram_mem[77918] = 16'b0000000000000000;
	sram_mem[77919] = 16'b0000000000000000;
	sram_mem[77920] = 16'b0000000000000000;
	sram_mem[77921] = 16'b0000000000000000;
	sram_mem[77922] = 16'b0000000000000000;
	sram_mem[77923] = 16'b0000000000000000;
	sram_mem[77924] = 16'b0000000000000000;
	sram_mem[77925] = 16'b0000000000000000;
	sram_mem[77926] = 16'b0000000000000000;
	sram_mem[77927] = 16'b0000000000000000;
	sram_mem[77928] = 16'b0000000000000000;
	sram_mem[77929] = 16'b0000000000000000;
	sram_mem[77930] = 16'b0000000000000000;
	sram_mem[77931] = 16'b0000000000000000;
	sram_mem[77932] = 16'b0000000000000000;
	sram_mem[77933] = 16'b0000000000000000;
	sram_mem[77934] = 16'b0000000000000000;
	sram_mem[77935] = 16'b0000000000000000;
	sram_mem[77936] = 16'b0000000000000000;
	sram_mem[77937] = 16'b0000000000000000;
	sram_mem[77938] = 16'b0000000000000000;
	sram_mem[77939] = 16'b0000000000000000;
	sram_mem[77940] = 16'b0000000000000000;
	sram_mem[77941] = 16'b0000000000000000;
	sram_mem[77942] = 16'b0000000000000000;
	sram_mem[77943] = 16'b0000000000000000;
	sram_mem[77944] = 16'b0000000000000000;
	sram_mem[77945] = 16'b0000000000000000;
	sram_mem[77946] = 16'b0000000000000000;
	sram_mem[77947] = 16'b0000000000000000;
	sram_mem[77948] = 16'b0000000000000000;
	sram_mem[77949] = 16'b0000000000000000;
	sram_mem[77950] = 16'b0000000000000000;
	sram_mem[77951] = 16'b0000000000000000;
	sram_mem[77952] = 16'b0000000000000000;
	sram_mem[77953] = 16'b0000000000000000;
	sram_mem[77954] = 16'b0000000000000000;
	sram_mem[77955] = 16'b0000000000000000;
	sram_mem[77956] = 16'b0000000000000000;
	sram_mem[77957] = 16'b0000000000000000;
	sram_mem[77958] = 16'b0000000000000000;
	sram_mem[77959] = 16'b0000000000000000;
	sram_mem[77960] = 16'b0000000000000000;
	sram_mem[77961] = 16'b0000000000000000;
	sram_mem[77962] = 16'b0000000000000000;
	sram_mem[77963] = 16'b0000000000000000;
	sram_mem[77964] = 16'b0000000000000000;
	sram_mem[77965] = 16'b0000000000000000;
	sram_mem[77966] = 16'b0000000000000000;
	sram_mem[77967] = 16'b0000000000000000;
	sram_mem[77968] = 16'b0000000000000000;
	sram_mem[77969] = 16'b0000000000000000;
	sram_mem[77970] = 16'b0000000000000000;
	sram_mem[77971] = 16'b0000000000000000;
	sram_mem[77972] = 16'b0000000000000000;
	sram_mem[77973] = 16'b0000000000000000;
	sram_mem[77974] = 16'b0000000000000000;
	sram_mem[77975] = 16'b0000000000000000;
	sram_mem[77976] = 16'b0000000000000000;
	sram_mem[77977] = 16'b0000000000000000;
	sram_mem[77978] = 16'b0000000000000000;
	sram_mem[77979] = 16'b0000000000000000;
	sram_mem[77980] = 16'b0000000000000000;
	sram_mem[77981] = 16'b0000000000000000;
	sram_mem[77982] = 16'b0000000000000000;
	sram_mem[77983] = 16'b0000000000000000;
	sram_mem[77984] = 16'b0000000000000000;
	sram_mem[77985] = 16'b0000000000000000;
	sram_mem[77986] = 16'b0000000000000000;
	sram_mem[77987] = 16'b0000000000000000;
	sram_mem[77988] = 16'b0000000000000000;
	sram_mem[77989] = 16'b0000000000000000;
	sram_mem[77990] = 16'b0000000000000000;
	sram_mem[77991] = 16'b0000000000000000;
	sram_mem[77992] = 16'b0000000000000000;
	sram_mem[77993] = 16'b0000000000000000;
	sram_mem[77994] = 16'b0000000000000000;
	sram_mem[77995] = 16'b0000000000000000;
	sram_mem[77996] = 16'b0000000000000000;
	sram_mem[77997] = 16'b0000000000000000;
	sram_mem[77998] = 16'b0000000000000000;
	sram_mem[77999] = 16'b0000000000000000;
	sram_mem[78000] = 16'b0000000000000000;
	sram_mem[78001] = 16'b0000000000000000;
	sram_mem[78002] = 16'b0000000000000000;
	sram_mem[78003] = 16'b0000000000000000;
	sram_mem[78004] = 16'b0000000000000000;
	sram_mem[78005] = 16'b0000000000000000;
	sram_mem[78006] = 16'b0000000000000000;
	sram_mem[78007] = 16'b0000000000000000;
	sram_mem[78008] = 16'b0000000000000000;
	sram_mem[78009] = 16'b0000000000000000;
	sram_mem[78010] = 16'b0000000000000000;
	sram_mem[78011] = 16'b0000000000000000;
	sram_mem[78012] = 16'b0000000000000000;
	sram_mem[78013] = 16'b0000000000000000;
	sram_mem[78014] = 16'b0000000000000000;
	sram_mem[78015] = 16'b0000000000000000;
	sram_mem[78016] = 16'b0000000000000000;
	sram_mem[78017] = 16'b0000000000000000;
	sram_mem[78018] = 16'b0000000000000000;
	sram_mem[78019] = 16'b0000000000000000;
	sram_mem[78020] = 16'b0000000000000000;
	sram_mem[78021] = 16'b0000000000000000;
	sram_mem[78022] = 16'b0000000000000000;
	sram_mem[78023] = 16'b0000000000000000;
	sram_mem[78024] = 16'b0000000000000000;
	sram_mem[78025] = 16'b0000000000000000;
	sram_mem[78026] = 16'b0000000000000000;
	sram_mem[78027] = 16'b0000000000000000;
	sram_mem[78028] = 16'b0000000000000000;
	sram_mem[78029] = 16'b0000000000000000;
	sram_mem[78030] = 16'b0000000000000000;
	sram_mem[78031] = 16'b0000000000000000;
	sram_mem[78032] = 16'b0000000000000000;
	sram_mem[78033] = 16'b0000000000000000;
	sram_mem[78034] = 16'b0000000000000000;
	sram_mem[78035] = 16'b0000000000000000;
	sram_mem[78036] = 16'b0000000000000000;
	sram_mem[78037] = 16'b0000000000000000;
	sram_mem[78038] = 16'b0000000000000000;
	sram_mem[78039] = 16'b0000000000000000;
	sram_mem[78040] = 16'b0000000000000000;
	sram_mem[78041] = 16'b0000000000000000;
	sram_mem[78042] = 16'b0000000000000000;
	sram_mem[78043] = 16'b0000000000000000;
	sram_mem[78044] = 16'b0000000000000000;
	sram_mem[78045] = 16'b0000000000000000;
	sram_mem[78046] = 16'b0000000000000000;
	sram_mem[78047] = 16'b0000000000000000;
	sram_mem[78048] = 16'b0000000000000000;
	sram_mem[78049] = 16'b0000000000000000;
	sram_mem[78050] = 16'b0000000000000000;
	sram_mem[78051] = 16'b0000000000000000;
	sram_mem[78052] = 16'b0000000000000000;
	sram_mem[78053] = 16'b0000000000000000;
	sram_mem[78054] = 16'b0000000000000000;
	sram_mem[78055] = 16'b0000000000000000;
	sram_mem[78056] = 16'b0000000000000000;
	sram_mem[78057] = 16'b0000000000000000;
	sram_mem[78058] = 16'b0000000000000000;
	sram_mem[78059] = 16'b0000000000000000;
	sram_mem[78060] = 16'b0000000000000000;
	sram_mem[78061] = 16'b0000000000000000;
	sram_mem[78062] = 16'b0000000000000000;
	sram_mem[78063] = 16'b0000000000000000;
	sram_mem[78064] = 16'b0000000000000000;
	sram_mem[78065] = 16'b0000000000000000;
	sram_mem[78066] = 16'b0000000000000000;
	sram_mem[78067] = 16'b0000000000000000;
	sram_mem[78068] = 16'b0000000000000000;
	sram_mem[78069] = 16'b0000000000000000;
	sram_mem[78070] = 16'b0000000000000000;
	sram_mem[78071] = 16'b0000000000000000;
	sram_mem[78072] = 16'b0000000000000000;
	sram_mem[78073] = 16'b0000000000000000;
	sram_mem[78074] = 16'b0000000000000000;
	sram_mem[78075] = 16'b0000000000000000;
	sram_mem[78076] = 16'b0000000000000000;
	sram_mem[78077] = 16'b0000000000000000;
	sram_mem[78078] = 16'b0000000000000000;
	sram_mem[78079] = 16'b0000000000000000;
	sram_mem[78080] = 16'b0000000000000000;
	sram_mem[78081] = 16'b0000000000000000;
	sram_mem[78082] = 16'b0000000000000000;
	sram_mem[78083] = 16'b0000000000000000;
	sram_mem[78084] = 16'b0000000000000000;
	sram_mem[78085] = 16'b0000000000000000;
	sram_mem[78086] = 16'b0000000000000000;
	sram_mem[78087] = 16'b0000000000000000;
	sram_mem[78088] = 16'b0000000000000000;
	sram_mem[78089] = 16'b0000000000000000;
	sram_mem[78090] = 16'b0000000000000000;
	sram_mem[78091] = 16'b0000000000000000;
	sram_mem[78092] = 16'b0000000000000000;
	sram_mem[78093] = 16'b0000000000000000;
	sram_mem[78094] = 16'b0000000000000000;
	sram_mem[78095] = 16'b0000000000000000;
	sram_mem[78096] = 16'b0000000000000000;
	sram_mem[78097] = 16'b0000000000000000;
	sram_mem[78098] = 16'b0000000000000000;
	sram_mem[78099] = 16'b0000000000000000;
	sram_mem[78100] = 16'b0000000000000000;
	sram_mem[78101] = 16'b0000000000000000;
	sram_mem[78102] = 16'b0000000000000000;
	sram_mem[78103] = 16'b0000000000000000;
	sram_mem[78104] = 16'b0000000000000000;
	sram_mem[78105] = 16'b0000000000000000;
	sram_mem[78106] = 16'b0000000000000000;
	sram_mem[78107] = 16'b0000000000000000;
	sram_mem[78108] = 16'b0000000000000000;
	sram_mem[78109] = 16'b0000000000000000;
	sram_mem[78110] = 16'b0000000000000000;
	sram_mem[78111] = 16'b0000000000000000;
	sram_mem[78112] = 16'b0000000000000000;
	sram_mem[78113] = 16'b0000000000000000;
	sram_mem[78114] = 16'b0000000000000000;
	sram_mem[78115] = 16'b0000000000000000;
	sram_mem[78116] = 16'b0000000000000000;
	sram_mem[78117] = 16'b0000000000000000;
	sram_mem[78118] = 16'b0000000000000000;
	sram_mem[78119] = 16'b0000000000000000;
	sram_mem[78120] = 16'b0000000000000000;
	sram_mem[78121] = 16'b0000000000000000;
	sram_mem[78122] = 16'b0000000000000000;
	sram_mem[78123] = 16'b0000000000000000;
	sram_mem[78124] = 16'b0000000000000000;
	sram_mem[78125] = 16'b0000000000000000;
	sram_mem[78126] = 16'b0000000000000000;
	sram_mem[78127] = 16'b0000000000000000;
	sram_mem[78128] = 16'b0000000000000000;
	sram_mem[78129] = 16'b0000000000000000;
	sram_mem[78130] = 16'b0000000000000000;
	sram_mem[78131] = 16'b0000000000000000;
	sram_mem[78132] = 16'b0000000000000000;
	sram_mem[78133] = 16'b0000000000000000;
	sram_mem[78134] = 16'b0000000000000000;
	sram_mem[78135] = 16'b0000000000000000;
	sram_mem[78136] = 16'b0000000000000000;
	sram_mem[78137] = 16'b0000000000000000;
	sram_mem[78138] = 16'b0000000000000000;
	sram_mem[78139] = 16'b0000000000000000;
	sram_mem[78140] = 16'b0000000000000000;
	sram_mem[78141] = 16'b0000000000000000;
	sram_mem[78142] = 16'b0000000000000000;
	sram_mem[78143] = 16'b0000000000000000;
	sram_mem[78144] = 16'b0000000000000000;
	sram_mem[78145] = 16'b0000000000000000;
	sram_mem[78146] = 16'b0000000000000000;
	sram_mem[78147] = 16'b0000000000000000;
	sram_mem[78148] = 16'b0000000000000000;
	sram_mem[78149] = 16'b0000000000000000;
	sram_mem[78150] = 16'b0000000000000000;
	sram_mem[78151] = 16'b0000000000000000;
	sram_mem[78152] = 16'b0000000000000000;
	sram_mem[78153] = 16'b0000000000000000;
	sram_mem[78154] = 16'b0000000000000000;
	sram_mem[78155] = 16'b0000000000000000;
	sram_mem[78156] = 16'b0000000000000000;
	sram_mem[78157] = 16'b0000000000000000;
	sram_mem[78158] = 16'b0000000000000000;
	sram_mem[78159] = 16'b0000000000000000;
	sram_mem[78160] = 16'b0000000000000000;
	sram_mem[78161] = 16'b0000000000000000;
	sram_mem[78162] = 16'b0000000000000000;
	sram_mem[78163] = 16'b0000000000000000;
	sram_mem[78164] = 16'b0000000000000000;
	sram_mem[78165] = 16'b0000000000000000;
	sram_mem[78166] = 16'b0000000000000000;
	sram_mem[78167] = 16'b0000000000000000;
	sram_mem[78168] = 16'b0000000000000000;
	sram_mem[78169] = 16'b0000000000000000;
	sram_mem[78170] = 16'b0000000000000000;
	sram_mem[78171] = 16'b0000000000000000;
	sram_mem[78172] = 16'b0000000000000000;
	sram_mem[78173] = 16'b0000000000000000;
	sram_mem[78174] = 16'b0000000000000000;
	sram_mem[78175] = 16'b0000000000000000;
	sram_mem[78176] = 16'b0000000000000000;
	sram_mem[78177] = 16'b0000000000000000;
	sram_mem[78178] = 16'b0000000000000000;
	sram_mem[78179] = 16'b0000000000000000;
	sram_mem[78180] = 16'b0000000000000000;
	sram_mem[78181] = 16'b0000000000000000;
	sram_mem[78182] = 16'b0000000000000000;
	sram_mem[78183] = 16'b0000000000000000;
	sram_mem[78184] = 16'b0000000000000000;
	sram_mem[78185] = 16'b0000000000000000;
	sram_mem[78186] = 16'b0000000000000000;
	sram_mem[78187] = 16'b0000000000000000;
	sram_mem[78188] = 16'b0000000000000000;
	sram_mem[78189] = 16'b0000000000000000;
	sram_mem[78190] = 16'b0000000000000000;
	sram_mem[78191] = 16'b0000000000000000;
	sram_mem[78192] = 16'b0000000000000000;
	sram_mem[78193] = 16'b0000000000000000;
	sram_mem[78194] = 16'b0000000000000000;
	sram_mem[78195] = 16'b0000000000000000;
	sram_mem[78196] = 16'b0000000000000000;
	sram_mem[78197] = 16'b0000000000000000;
	sram_mem[78198] = 16'b0000000000000000;
	sram_mem[78199] = 16'b0000000000000000;
	sram_mem[78200] = 16'b0000000000000000;
	sram_mem[78201] = 16'b0000000000000000;
	sram_mem[78202] = 16'b0000000000000000;
	sram_mem[78203] = 16'b0000000000000000;
	sram_mem[78204] = 16'b0000000000000000;
	sram_mem[78205] = 16'b0000000000000000;
	sram_mem[78206] = 16'b0000000000000000;
	sram_mem[78207] = 16'b0000000000000000;
	sram_mem[78208] = 16'b0000000000000000;
	sram_mem[78209] = 16'b0000000000000000;
	sram_mem[78210] = 16'b0000000000000000;
	sram_mem[78211] = 16'b0000000000000000;
	sram_mem[78212] = 16'b0000000000000000;
	sram_mem[78213] = 16'b0000000000000000;
	sram_mem[78214] = 16'b0000000000000000;
	sram_mem[78215] = 16'b0000000000000000;
	sram_mem[78216] = 16'b0000000000000000;
	sram_mem[78217] = 16'b0000000000000000;
	sram_mem[78218] = 16'b0000000000000000;
	sram_mem[78219] = 16'b0000000000000000;
	sram_mem[78220] = 16'b0000000000000000;
	sram_mem[78221] = 16'b0000000000000000;
	sram_mem[78222] = 16'b0000000000000000;
	sram_mem[78223] = 16'b0000000000000000;
	sram_mem[78224] = 16'b0000000000000000;
	sram_mem[78225] = 16'b0000000000000000;
	sram_mem[78226] = 16'b0000000000000000;
	sram_mem[78227] = 16'b0000000000000000;
	sram_mem[78228] = 16'b0000000000000000;
	sram_mem[78229] = 16'b0000000000000000;
	sram_mem[78230] = 16'b0000000000000000;
	sram_mem[78231] = 16'b0000000000000000;
	sram_mem[78232] = 16'b0000000000000000;
	sram_mem[78233] = 16'b0000000000000000;
	sram_mem[78234] = 16'b0000000000000000;
	sram_mem[78235] = 16'b0000000000000000;
	sram_mem[78236] = 16'b0000000000000000;
	sram_mem[78237] = 16'b0000000000000000;
	sram_mem[78238] = 16'b0000000000000000;
	sram_mem[78239] = 16'b0000000000000000;
	sram_mem[78240] = 16'b0000000000000000;
	sram_mem[78241] = 16'b0000000000000000;
	sram_mem[78242] = 16'b0000000000000000;
	sram_mem[78243] = 16'b0000000000000000;
	sram_mem[78244] = 16'b0000000000000000;
	sram_mem[78245] = 16'b0000000000000000;
	sram_mem[78246] = 16'b0000000000000000;
	sram_mem[78247] = 16'b0000000000000000;
	sram_mem[78248] = 16'b0000000000000000;
	sram_mem[78249] = 16'b0000000000000000;
	sram_mem[78250] = 16'b0000000000000000;
	sram_mem[78251] = 16'b0000000000000000;
	sram_mem[78252] = 16'b0000000000000000;
	sram_mem[78253] = 16'b0000000000000000;
	sram_mem[78254] = 16'b0000000000000000;
	sram_mem[78255] = 16'b0000000000000000;
	sram_mem[78256] = 16'b0000000000000000;
	sram_mem[78257] = 16'b0000000000000000;
	sram_mem[78258] = 16'b0000000000000000;
	sram_mem[78259] = 16'b0000000000000000;
	sram_mem[78260] = 16'b0000000000000000;
	sram_mem[78261] = 16'b0000000000000000;
	sram_mem[78262] = 16'b0000000000000000;
	sram_mem[78263] = 16'b0000000000000000;
	sram_mem[78264] = 16'b0000000000000000;
	sram_mem[78265] = 16'b0000000000000000;
	sram_mem[78266] = 16'b0000000000000000;
	sram_mem[78267] = 16'b0000000000000000;
	sram_mem[78268] = 16'b0000000000000000;
	sram_mem[78269] = 16'b0000000000000000;
	sram_mem[78270] = 16'b0000000000000000;
	sram_mem[78271] = 16'b0000000000000000;
	sram_mem[78272] = 16'b0000000000000000;
	sram_mem[78273] = 16'b0000000000000000;
	sram_mem[78274] = 16'b0000000000000000;
	sram_mem[78275] = 16'b0000000000000000;
	sram_mem[78276] = 16'b0000000000000000;
	sram_mem[78277] = 16'b0000000000000000;
	sram_mem[78278] = 16'b0000000000000000;
	sram_mem[78279] = 16'b0000000000000000;
	sram_mem[78280] = 16'b0000000000000000;
	sram_mem[78281] = 16'b0000000000000000;
	sram_mem[78282] = 16'b0000000000000000;
	sram_mem[78283] = 16'b0000000000000000;
	sram_mem[78284] = 16'b0000000000000000;
	sram_mem[78285] = 16'b0000000000000000;
	sram_mem[78286] = 16'b0000000000000000;
	sram_mem[78287] = 16'b0000000000000000;
	sram_mem[78288] = 16'b0000000000000000;
	sram_mem[78289] = 16'b0000000000000000;
	sram_mem[78290] = 16'b0000000000000000;
	sram_mem[78291] = 16'b0000000000000000;
	sram_mem[78292] = 16'b0000000000000000;
	sram_mem[78293] = 16'b0000000000000000;
	sram_mem[78294] = 16'b0000000000000000;
	sram_mem[78295] = 16'b0000000000000000;
	sram_mem[78296] = 16'b0000000000000000;
	sram_mem[78297] = 16'b0000000000000000;
	sram_mem[78298] = 16'b0000000000000000;
	sram_mem[78299] = 16'b0000000000000000;
	sram_mem[78300] = 16'b0000000000000000;
	sram_mem[78301] = 16'b0000000000000000;
	sram_mem[78302] = 16'b0000000000000000;
	sram_mem[78303] = 16'b0000000000000000;
	sram_mem[78304] = 16'b0000000000000000;
	sram_mem[78305] = 16'b0000000000000000;
	sram_mem[78306] = 16'b0000000000000000;
	sram_mem[78307] = 16'b0000000000000000;
	sram_mem[78308] = 16'b0000000000000000;
	sram_mem[78309] = 16'b0000000000000000;
	sram_mem[78310] = 16'b0000000000000000;
	sram_mem[78311] = 16'b0000000000000000;
	sram_mem[78312] = 16'b0000000000000000;
	sram_mem[78313] = 16'b0000000000000000;
	sram_mem[78314] = 16'b0000000000000000;
	sram_mem[78315] = 16'b0000000000000000;
	sram_mem[78316] = 16'b0000000000000000;
	sram_mem[78317] = 16'b0000000000000000;
	sram_mem[78318] = 16'b0000000000000000;
	sram_mem[78319] = 16'b0000000000000000;
	sram_mem[78320] = 16'b0000000000000000;
	sram_mem[78321] = 16'b0000000000000000;
	sram_mem[78322] = 16'b0000000000000000;
	sram_mem[78323] = 16'b0000000000000000;
	sram_mem[78324] = 16'b0000000000000000;
	sram_mem[78325] = 16'b0000000000000000;
	sram_mem[78326] = 16'b0000000000000000;
	sram_mem[78327] = 16'b0000000000000000;
	sram_mem[78328] = 16'b0000000000000000;
	sram_mem[78329] = 16'b0000000000000000;
	sram_mem[78330] = 16'b0000000000000000;
	sram_mem[78331] = 16'b0000000000000000;
	sram_mem[78332] = 16'b0000000000000000;
	sram_mem[78333] = 16'b0000000000000000;
	sram_mem[78334] = 16'b0000000000000000;
	sram_mem[78335] = 16'b0000000000000000;
	sram_mem[78336] = 16'b0000000000000000;
	sram_mem[78337] = 16'b0000000000000000;
	sram_mem[78338] = 16'b0000000000000000;
	sram_mem[78339] = 16'b0000000000000000;
	sram_mem[78340] = 16'b0000000000000000;
	sram_mem[78341] = 16'b0000000000000000;
	sram_mem[78342] = 16'b0000000000000000;
	sram_mem[78343] = 16'b0000000000000000;
	sram_mem[78344] = 16'b0000000000000000;
	sram_mem[78345] = 16'b0000000000000000;
	sram_mem[78346] = 16'b0000000000000000;
	sram_mem[78347] = 16'b0000000000000000;
	sram_mem[78348] = 16'b0000000000000000;
	sram_mem[78349] = 16'b0000000000000000;
	sram_mem[78350] = 16'b0000000000000000;
	sram_mem[78351] = 16'b0000000000000000;
	sram_mem[78352] = 16'b0000000000000000;
	sram_mem[78353] = 16'b0000000000000000;
	sram_mem[78354] = 16'b0000000000000000;
	sram_mem[78355] = 16'b0000000000000000;
	sram_mem[78356] = 16'b0000000000000000;
	sram_mem[78357] = 16'b0000000000000000;
	sram_mem[78358] = 16'b0000000000000000;
	sram_mem[78359] = 16'b0000000000000000;
	sram_mem[78360] = 16'b0000000000000000;
	sram_mem[78361] = 16'b0000000000000000;
	sram_mem[78362] = 16'b0000000000000000;
	sram_mem[78363] = 16'b0000000000000000;
	sram_mem[78364] = 16'b0000000000000000;
	sram_mem[78365] = 16'b0000000000000000;
	sram_mem[78366] = 16'b0000000000000000;
	sram_mem[78367] = 16'b0000000000000000;
	sram_mem[78368] = 16'b0000000000000000;
	sram_mem[78369] = 16'b0000000000000000;
	sram_mem[78370] = 16'b0000000000000000;
	sram_mem[78371] = 16'b0000000000000000;
	sram_mem[78372] = 16'b0000000000000000;
	sram_mem[78373] = 16'b0000000000000000;
	sram_mem[78374] = 16'b0000000000000000;
	sram_mem[78375] = 16'b0000000000000000;
	sram_mem[78376] = 16'b0000000000000000;
	sram_mem[78377] = 16'b0000000000000000;
	sram_mem[78378] = 16'b0000000000000000;
	sram_mem[78379] = 16'b0000000000000000;
	sram_mem[78380] = 16'b0000000000000000;
	sram_mem[78381] = 16'b0000000000000000;
	sram_mem[78382] = 16'b0000000000000000;
	sram_mem[78383] = 16'b0000000000000000;
	sram_mem[78384] = 16'b0000000000000000;
	sram_mem[78385] = 16'b0000000000000000;
	sram_mem[78386] = 16'b0000000000000000;
	sram_mem[78387] = 16'b0000000000000000;
	sram_mem[78388] = 16'b0000000000000000;
	sram_mem[78389] = 16'b0000000000000000;
	sram_mem[78390] = 16'b0000000000000000;
	sram_mem[78391] = 16'b0000000000000000;
	sram_mem[78392] = 16'b0000000000000000;
	sram_mem[78393] = 16'b0000000000000000;
	sram_mem[78394] = 16'b0000000000000000;
	sram_mem[78395] = 16'b0000000000000000;
	sram_mem[78396] = 16'b0000000000000000;
	sram_mem[78397] = 16'b0000000000000000;
	sram_mem[78398] = 16'b0000000000000000;
	sram_mem[78399] = 16'b0000000000000000;
	sram_mem[78400] = 16'b0000000000000000;
	sram_mem[78401] = 16'b0000000000000000;
	sram_mem[78402] = 16'b0000000000000000;
	sram_mem[78403] = 16'b0000000000000000;
	sram_mem[78404] = 16'b0000000000000000;
	sram_mem[78405] = 16'b0000000000000000;
	sram_mem[78406] = 16'b0000000000000000;
	sram_mem[78407] = 16'b0000000000000000;
	sram_mem[78408] = 16'b0000000000000000;
	sram_mem[78409] = 16'b0000000000000000;
	sram_mem[78410] = 16'b0000000000000000;
	sram_mem[78411] = 16'b0000000000000000;
	sram_mem[78412] = 16'b0000000000000000;
	sram_mem[78413] = 16'b0000000000000000;
	sram_mem[78414] = 16'b0000000000000000;
	sram_mem[78415] = 16'b0000000000000000;
	sram_mem[78416] = 16'b0000000000000000;
	sram_mem[78417] = 16'b0000000000000000;
	sram_mem[78418] = 16'b0000000000000000;
	sram_mem[78419] = 16'b0000000000000000;
	sram_mem[78420] = 16'b0000000000000000;
	sram_mem[78421] = 16'b0000000000000000;
	sram_mem[78422] = 16'b0000000000000000;
	sram_mem[78423] = 16'b0000000000000000;
	sram_mem[78424] = 16'b0000000000000000;
	sram_mem[78425] = 16'b0000000000000000;
	sram_mem[78426] = 16'b0000000000000000;
	sram_mem[78427] = 16'b0000000000000000;
	sram_mem[78428] = 16'b0000000000000000;
	sram_mem[78429] = 16'b0000000000000000;
	sram_mem[78430] = 16'b0000000000000000;
	sram_mem[78431] = 16'b0000000000000000;
	sram_mem[78432] = 16'b0000000000000000;
	sram_mem[78433] = 16'b0000000000000000;
	sram_mem[78434] = 16'b0000000000000000;
	sram_mem[78435] = 16'b0000000000000000;
	sram_mem[78436] = 16'b0000000000000000;
	sram_mem[78437] = 16'b0000000000000000;
	sram_mem[78438] = 16'b0000000000000000;
	sram_mem[78439] = 16'b0000000000000000;
	sram_mem[78440] = 16'b0000000000000000;
	sram_mem[78441] = 16'b0000000000000000;
	sram_mem[78442] = 16'b0000000000000000;
	sram_mem[78443] = 16'b0000000000000000;
	sram_mem[78444] = 16'b0000000000000000;
	sram_mem[78445] = 16'b0000000000000000;
	sram_mem[78446] = 16'b0000000000000000;
	sram_mem[78447] = 16'b0000000000000000;
	sram_mem[78448] = 16'b0000000000000000;
	sram_mem[78449] = 16'b0000000000000000;
	sram_mem[78450] = 16'b0000000000000000;
	sram_mem[78451] = 16'b0000000000000000;
	sram_mem[78452] = 16'b0000000000000000;
	sram_mem[78453] = 16'b0000000000000000;
	sram_mem[78454] = 16'b0000000000000000;
	sram_mem[78455] = 16'b0000000000000000;
	sram_mem[78456] = 16'b0000000000000000;
	sram_mem[78457] = 16'b0000000000000000;
	sram_mem[78458] = 16'b0000000000000000;
	sram_mem[78459] = 16'b0000000000000000;
	sram_mem[78460] = 16'b0000000000000000;
	sram_mem[78461] = 16'b0000000000000000;
	sram_mem[78462] = 16'b0000000000000000;
	sram_mem[78463] = 16'b0000000000000000;
	sram_mem[78464] = 16'b0000000000000000;
	sram_mem[78465] = 16'b0000000000000000;
	sram_mem[78466] = 16'b0000000000000000;
	sram_mem[78467] = 16'b0000000000000000;
	sram_mem[78468] = 16'b0000000000000000;
	sram_mem[78469] = 16'b0000000000000000;
	sram_mem[78470] = 16'b0000000000000000;
	sram_mem[78471] = 16'b0000000000000000;
	sram_mem[78472] = 16'b0000000000000000;
	sram_mem[78473] = 16'b0000000000000000;
	sram_mem[78474] = 16'b0000000000000000;
	sram_mem[78475] = 16'b0000000000000000;
	sram_mem[78476] = 16'b0000000000000000;
	sram_mem[78477] = 16'b0000000000000000;
	sram_mem[78478] = 16'b0000000000000000;
	sram_mem[78479] = 16'b0000000000000000;
	sram_mem[78480] = 16'b0000000000000000;
	sram_mem[78481] = 16'b0000000000000000;
	sram_mem[78482] = 16'b0000000000000000;
	sram_mem[78483] = 16'b0000000000000000;
	sram_mem[78484] = 16'b0000000000000000;
	sram_mem[78485] = 16'b0000000000000000;
	sram_mem[78486] = 16'b0000000000000000;
	sram_mem[78487] = 16'b0000000000000000;
	sram_mem[78488] = 16'b0000000000000000;
	sram_mem[78489] = 16'b0000000000000000;
	sram_mem[78490] = 16'b0000000000000000;
	sram_mem[78491] = 16'b0000000000000000;
	sram_mem[78492] = 16'b0000000000000000;
	sram_mem[78493] = 16'b0000000000000000;
	sram_mem[78494] = 16'b0000000000000000;
	sram_mem[78495] = 16'b0000000000000000;
	sram_mem[78496] = 16'b0000000000000000;
	sram_mem[78497] = 16'b0000000000000000;
	sram_mem[78498] = 16'b0000000000000000;
	sram_mem[78499] = 16'b0000000000000000;
	sram_mem[78500] = 16'b0000000000000000;
	sram_mem[78501] = 16'b0000000000000000;
	sram_mem[78502] = 16'b0000000000000000;
	sram_mem[78503] = 16'b0000000000000000;
	sram_mem[78504] = 16'b0000000000000000;
	sram_mem[78505] = 16'b0000000000000000;
	sram_mem[78506] = 16'b0000000000000000;
	sram_mem[78507] = 16'b0000000000000000;
	sram_mem[78508] = 16'b0000000000000000;
	sram_mem[78509] = 16'b0000000000000000;
	sram_mem[78510] = 16'b0000000000000000;
	sram_mem[78511] = 16'b0000000000000000;
	sram_mem[78512] = 16'b0000000000000000;
	sram_mem[78513] = 16'b0000000000000000;
	sram_mem[78514] = 16'b0000000000000000;
	sram_mem[78515] = 16'b0000000000000000;
	sram_mem[78516] = 16'b0000000000000000;
	sram_mem[78517] = 16'b0000000000000000;
	sram_mem[78518] = 16'b0000000000000000;
	sram_mem[78519] = 16'b0000000000000000;
	sram_mem[78520] = 16'b0000000000000000;
	sram_mem[78521] = 16'b0000000000000000;
	sram_mem[78522] = 16'b0000000000000000;
	sram_mem[78523] = 16'b0000000000000000;
	sram_mem[78524] = 16'b0000000000000000;
	sram_mem[78525] = 16'b0000000000000000;
	sram_mem[78526] = 16'b0000000000000000;
	sram_mem[78527] = 16'b0000000000000000;
	sram_mem[78528] = 16'b0000000000000000;
	sram_mem[78529] = 16'b0000000000000000;
	sram_mem[78530] = 16'b0000000000000000;
	sram_mem[78531] = 16'b0000000000000000;
	sram_mem[78532] = 16'b0000000000000000;
	sram_mem[78533] = 16'b0000000000000000;
	sram_mem[78534] = 16'b0000000000000000;
	sram_mem[78535] = 16'b0000000000000000;
	sram_mem[78536] = 16'b0000000000000000;
	sram_mem[78537] = 16'b0000000000000000;
	sram_mem[78538] = 16'b0000000000000000;
	sram_mem[78539] = 16'b0000000000000000;
	sram_mem[78540] = 16'b0000000000000000;
	sram_mem[78541] = 16'b0000000000000000;
	sram_mem[78542] = 16'b0000000000000000;
	sram_mem[78543] = 16'b0000000000000000;
	sram_mem[78544] = 16'b0000000000000000;
	sram_mem[78545] = 16'b0000000000000000;
	sram_mem[78546] = 16'b0000000000000000;
	sram_mem[78547] = 16'b0000000000000000;
	sram_mem[78548] = 16'b0000000000000000;
	sram_mem[78549] = 16'b0000000000000000;
	sram_mem[78550] = 16'b0000000000000000;
	sram_mem[78551] = 16'b0000000000000000;
	sram_mem[78552] = 16'b0000000000000000;
	sram_mem[78553] = 16'b0000000000000000;
	sram_mem[78554] = 16'b0000000000000000;
	sram_mem[78555] = 16'b0000000000000000;
	sram_mem[78556] = 16'b0000000000000000;
	sram_mem[78557] = 16'b0000000000000000;
	sram_mem[78558] = 16'b0000000000000000;
	sram_mem[78559] = 16'b0000000000000000;
	sram_mem[78560] = 16'b0000000000000000;
	sram_mem[78561] = 16'b0000000000000000;
	sram_mem[78562] = 16'b0000000000000000;
	sram_mem[78563] = 16'b0000000000000000;
	sram_mem[78564] = 16'b0000000000000000;
	sram_mem[78565] = 16'b0000000000000000;
	sram_mem[78566] = 16'b0000000000000000;
	sram_mem[78567] = 16'b0000000000000000;
	sram_mem[78568] = 16'b0000000000000000;
	sram_mem[78569] = 16'b0000000000000000;
	sram_mem[78570] = 16'b0000000000000000;
	sram_mem[78571] = 16'b0000000000000000;
	sram_mem[78572] = 16'b0000000000000000;
	sram_mem[78573] = 16'b0000000000000000;
	sram_mem[78574] = 16'b0000000000000000;
	sram_mem[78575] = 16'b0000000000000000;
	sram_mem[78576] = 16'b0000000000000000;
	sram_mem[78577] = 16'b0000000000000000;
	sram_mem[78578] = 16'b0000000000000000;
	sram_mem[78579] = 16'b0000000000000000;
	sram_mem[78580] = 16'b0000000000000000;
	sram_mem[78581] = 16'b0000000000000000;
	sram_mem[78582] = 16'b0000000000000000;
	sram_mem[78583] = 16'b0000000000000000;
	sram_mem[78584] = 16'b0000000000000000;
	sram_mem[78585] = 16'b0000000000000000;
	sram_mem[78586] = 16'b0000000000000000;
	sram_mem[78587] = 16'b0000000000000000;
	sram_mem[78588] = 16'b0000000000000000;
	sram_mem[78589] = 16'b0000000000000000;
	sram_mem[78590] = 16'b0000000000000000;
	sram_mem[78591] = 16'b0000000000000000;
	sram_mem[78592] = 16'b0000000000000000;
	sram_mem[78593] = 16'b0000000000000000;
	sram_mem[78594] = 16'b0000000000000000;
	sram_mem[78595] = 16'b0000000000000000;
	sram_mem[78596] = 16'b0000000000000000;
	sram_mem[78597] = 16'b0000000000000000;
	sram_mem[78598] = 16'b0000000000000000;
	sram_mem[78599] = 16'b0000000000000000;
	sram_mem[78600] = 16'b0000000000000000;
	sram_mem[78601] = 16'b0000000000000000;
	sram_mem[78602] = 16'b0000000000000000;
	sram_mem[78603] = 16'b0000000000000000;
	sram_mem[78604] = 16'b0000000000000000;
	sram_mem[78605] = 16'b0000000000000000;
	sram_mem[78606] = 16'b0000000000000000;
	sram_mem[78607] = 16'b0000000000000000;
	sram_mem[78608] = 16'b0000000000000000;
	sram_mem[78609] = 16'b0000000000000000;
	sram_mem[78610] = 16'b0000000000000000;
	sram_mem[78611] = 16'b0000000000000000;
	sram_mem[78612] = 16'b0000000000000000;
	sram_mem[78613] = 16'b0000000000000000;
	sram_mem[78614] = 16'b0000000000000000;
	sram_mem[78615] = 16'b0000000000000000;
	sram_mem[78616] = 16'b0000000000000000;
	sram_mem[78617] = 16'b0000000000000000;
	sram_mem[78618] = 16'b0000000000000000;
	sram_mem[78619] = 16'b0000000000000000;
	sram_mem[78620] = 16'b0000000000000000;
	sram_mem[78621] = 16'b0000000000000000;
	sram_mem[78622] = 16'b0000000000000000;
	sram_mem[78623] = 16'b0000000000000000;
	sram_mem[78624] = 16'b0000000000000000;
	sram_mem[78625] = 16'b0000000000000000;
	sram_mem[78626] = 16'b0000000000000000;
	sram_mem[78627] = 16'b0000000000000000;
	sram_mem[78628] = 16'b0000000000000000;
	sram_mem[78629] = 16'b0000000000000000;
	sram_mem[78630] = 16'b0000000000000000;
	sram_mem[78631] = 16'b0000000000000000;
	sram_mem[78632] = 16'b0000000000000000;
	sram_mem[78633] = 16'b0000000000000000;
	sram_mem[78634] = 16'b0000000000000000;
	sram_mem[78635] = 16'b0000000000000000;
	sram_mem[78636] = 16'b0000000000000000;
	sram_mem[78637] = 16'b0000000000000000;
	sram_mem[78638] = 16'b0000000000000000;
	sram_mem[78639] = 16'b0000000000000000;
	sram_mem[78640] = 16'b0000000000000000;
	sram_mem[78641] = 16'b0000000000000000;
	sram_mem[78642] = 16'b0000000000000000;
	sram_mem[78643] = 16'b0000000000000000;
	sram_mem[78644] = 16'b0000000000000000;
	sram_mem[78645] = 16'b0000000000000000;
	sram_mem[78646] = 16'b0000000000000000;
	sram_mem[78647] = 16'b0000000000000000;
	sram_mem[78648] = 16'b0000000000000000;
	sram_mem[78649] = 16'b0000000000000000;
	sram_mem[78650] = 16'b0000000000000000;
	sram_mem[78651] = 16'b0000000000000000;
	sram_mem[78652] = 16'b0000000000000000;
	sram_mem[78653] = 16'b0000000000000000;
	sram_mem[78654] = 16'b0000000000000000;
	sram_mem[78655] = 16'b0000000000000000;
	sram_mem[78656] = 16'b0000000000000000;
	sram_mem[78657] = 16'b0000000000000000;
	sram_mem[78658] = 16'b0000000000000000;
	sram_mem[78659] = 16'b0000000000000000;
	sram_mem[78660] = 16'b0000000000000000;
	sram_mem[78661] = 16'b0000000000000000;
	sram_mem[78662] = 16'b0000000000000000;
	sram_mem[78663] = 16'b0000000000000000;
	sram_mem[78664] = 16'b0000000000000000;
	sram_mem[78665] = 16'b0000000000000000;
	sram_mem[78666] = 16'b0000000000000000;
	sram_mem[78667] = 16'b0000000000000000;
	sram_mem[78668] = 16'b0000000000000000;
	sram_mem[78669] = 16'b0000000000000000;
	sram_mem[78670] = 16'b0000000000000000;
	sram_mem[78671] = 16'b0000000000000000;
	sram_mem[78672] = 16'b0000000000000000;
	sram_mem[78673] = 16'b0000000000000000;
	sram_mem[78674] = 16'b0000000000000000;
	sram_mem[78675] = 16'b0000000000000000;
	sram_mem[78676] = 16'b0000000000000000;
	sram_mem[78677] = 16'b0000000000000000;
	sram_mem[78678] = 16'b0000000000000000;
	sram_mem[78679] = 16'b0000000000000000;
	sram_mem[78680] = 16'b0000000000000000;
	sram_mem[78681] = 16'b0000000000000000;
	sram_mem[78682] = 16'b0000000000000000;
	sram_mem[78683] = 16'b0000000000000000;
	sram_mem[78684] = 16'b0000000000000000;
	sram_mem[78685] = 16'b0000000000000000;
	sram_mem[78686] = 16'b0000000000000000;
	sram_mem[78687] = 16'b0000000000000000;
	sram_mem[78688] = 16'b0000000000000000;
	sram_mem[78689] = 16'b0000000000000000;
	sram_mem[78690] = 16'b0000000000000000;
	sram_mem[78691] = 16'b0000000000000000;
	sram_mem[78692] = 16'b0000000000000000;
	sram_mem[78693] = 16'b0000000000000000;
	sram_mem[78694] = 16'b0000000000000000;
	sram_mem[78695] = 16'b0000000000000000;
	sram_mem[78696] = 16'b0000000000000000;
	sram_mem[78697] = 16'b0000000000000000;
	sram_mem[78698] = 16'b0000000000000000;
	sram_mem[78699] = 16'b0000000000000000;
	sram_mem[78700] = 16'b0000000000000000;
	sram_mem[78701] = 16'b0000000000000000;
	sram_mem[78702] = 16'b0000000000000000;
	sram_mem[78703] = 16'b0000000000000000;
	sram_mem[78704] = 16'b0000000000000000;
	sram_mem[78705] = 16'b0000000000000000;
	sram_mem[78706] = 16'b0000000000000000;
	sram_mem[78707] = 16'b0000000000000000;
	sram_mem[78708] = 16'b0000000000000000;
	sram_mem[78709] = 16'b0000000000000000;
	sram_mem[78710] = 16'b0000000000000000;
	sram_mem[78711] = 16'b0000000000000000;
	sram_mem[78712] = 16'b0000000000000000;
	sram_mem[78713] = 16'b0000000000000000;
	sram_mem[78714] = 16'b0000000000000000;
	sram_mem[78715] = 16'b0000000000000000;
	sram_mem[78716] = 16'b0000000000000000;
	sram_mem[78717] = 16'b0000000000000000;
	sram_mem[78718] = 16'b0000000000000000;
	sram_mem[78719] = 16'b0000000000000000;
	sram_mem[78720] = 16'b0000000000000000;
	sram_mem[78721] = 16'b0000000000000000;
	sram_mem[78722] = 16'b0000000000000000;
	sram_mem[78723] = 16'b0000000000000000;
	sram_mem[78724] = 16'b0000000000000000;
	sram_mem[78725] = 16'b0000000000000000;
	sram_mem[78726] = 16'b0000000000000000;
	sram_mem[78727] = 16'b0000000000000000;
	sram_mem[78728] = 16'b0000000000000000;
	sram_mem[78729] = 16'b0000000000000000;
	sram_mem[78730] = 16'b0000000000000000;
	sram_mem[78731] = 16'b0000000000000000;
	sram_mem[78732] = 16'b0000000000000000;
	sram_mem[78733] = 16'b0000000000000000;
	sram_mem[78734] = 16'b0000000000000000;
	sram_mem[78735] = 16'b0000000000000000;
	sram_mem[78736] = 16'b0000000000000000;
	sram_mem[78737] = 16'b0000000000000000;
	sram_mem[78738] = 16'b0000000000000000;
	sram_mem[78739] = 16'b0000000000000000;
	sram_mem[78740] = 16'b0000000000000000;
	sram_mem[78741] = 16'b0000000000000000;
	sram_mem[78742] = 16'b0000000000000000;
	sram_mem[78743] = 16'b0000000000000000;
	sram_mem[78744] = 16'b0000000000000000;
	sram_mem[78745] = 16'b0000000000000000;
	sram_mem[78746] = 16'b0000000000000000;
	sram_mem[78747] = 16'b0000000000000000;
	sram_mem[78748] = 16'b0000000000000000;
	sram_mem[78749] = 16'b0000000000000000;
	sram_mem[78750] = 16'b0000000000000000;
	sram_mem[78751] = 16'b0000000000000000;
	sram_mem[78752] = 16'b0000000000000000;
	sram_mem[78753] = 16'b0000000000000000;
	sram_mem[78754] = 16'b0000000000000000;
	sram_mem[78755] = 16'b0000000000000000;
	sram_mem[78756] = 16'b0000000000000000;
	sram_mem[78757] = 16'b0000000000000000;
	sram_mem[78758] = 16'b0000000000000000;
	sram_mem[78759] = 16'b0000000000000000;
	sram_mem[78760] = 16'b0000000000000000;
	sram_mem[78761] = 16'b0000000000000000;
	sram_mem[78762] = 16'b0000000000000000;
	sram_mem[78763] = 16'b0000000000000000;
	sram_mem[78764] = 16'b0000000000000000;
	sram_mem[78765] = 16'b0000000000000000;
	sram_mem[78766] = 16'b0000000000000000;
	sram_mem[78767] = 16'b0000000000000000;
	sram_mem[78768] = 16'b0000000000000000;
	sram_mem[78769] = 16'b0000000000000000;
	sram_mem[78770] = 16'b0000000000000000;
	sram_mem[78771] = 16'b0000000000000000;
	sram_mem[78772] = 16'b0000000000000000;
	sram_mem[78773] = 16'b0000000000000000;
	sram_mem[78774] = 16'b0000000000000000;
	sram_mem[78775] = 16'b0000000000000000;
	sram_mem[78776] = 16'b0000000000000000;
	sram_mem[78777] = 16'b0000000000000000;
	sram_mem[78778] = 16'b0000000000000000;
	sram_mem[78779] = 16'b0000000000000000;
	sram_mem[78780] = 16'b0000000000000000;
	sram_mem[78781] = 16'b0000000000000000;
	sram_mem[78782] = 16'b0000000000000000;
	sram_mem[78783] = 16'b0000000000000000;
	sram_mem[78784] = 16'b0000000000000000;
	sram_mem[78785] = 16'b0000000000000000;
	sram_mem[78786] = 16'b0000000000000000;
	sram_mem[78787] = 16'b0000000000000000;
	sram_mem[78788] = 16'b0000000000000000;
	sram_mem[78789] = 16'b0000000000000000;
	sram_mem[78790] = 16'b0000000000000000;
	sram_mem[78791] = 16'b0000000000000000;
	sram_mem[78792] = 16'b0000000000000000;
	sram_mem[78793] = 16'b0000000000000000;
	sram_mem[78794] = 16'b0000000000000000;
	sram_mem[78795] = 16'b0000000000000000;
	sram_mem[78796] = 16'b0000000000000000;
	sram_mem[78797] = 16'b0000000000000000;
	sram_mem[78798] = 16'b0000000000000000;
	sram_mem[78799] = 16'b0000000000000000;
	sram_mem[78800] = 16'b0000000000000000;
	sram_mem[78801] = 16'b0000000000000000;
	sram_mem[78802] = 16'b0000000000000000;
	sram_mem[78803] = 16'b0000000000000000;
	sram_mem[78804] = 16'b0000000000000000;
	sram_mem[78805] = 16'b0000000000000000;
	sram_mem[78806] = 16'b0000000000000000;
	sram_mem[78807] = 16'b0000000000000000;
	sram_mem[78808] = 16'b0000000000000000;
	sram_mem[78809] = 16'b0000000000000000;
	sram_mem[78810] = 16'b0000000000000000;
	sram_mem[78811] = 16'b0000000000000000;
	sram_mem[78812] = 16'b0000000000000000;
	sram_mem[78813] = 16'b0000000000000000;
	sram_mem[78814] = 16'b0000000000000000;
	sram_mem[78815] = 16'b0000000000000000;
	sram_mem[78816] = 16'b0000000000000000;
	sram_mem[78817] = 16'b0000000000000000;
	sram_mem[78818] = 16'b0000000000000000;
	sram_mem[78819] = 16'b0000000000000000;
	sram_mem[78820] = 16'b0000000000000000;
	sram_mem[78821] = 16'b0000000000000000;
	sram_mem[78822] = 16'b0000000000000000;
	sram_mem[78823] = 16'b0000000000000000;
	sram_mem[78824] = 16'b0000000000000000;
	sram_mem[78825] = 16'b0000000000000000;
	sram_mem[78826] = 16'b0000000000000000;
	sram_mem[78827] = 16'b0000000000000000;
	sram_mem[78828] = 16'b0000000000000000;
	sram_mem[78829] = 16'b0000000000000000;
	sram_mem[78830] = 16'b0000000000000000;
	sram_mem[78831] = 16'b0000000000000000;
	sram_mem[78832] = 16'b0000000000000000;
	sram_mem[78833] = 16'b0000000000000000;
	sram_mem[78834] = 16'b0000000000000000;
	sram_mem[78835] = 16'b0000000000000000;
	sram_mem[78836] = 16'b0000000000000000;
	sram_mem[78837] = 16'b0000000000000000;
	sram_mem[78838] = 16'b0000000000000000;
	sram_mem[78839] = 16'b0000000000000000;
	sram_mem[78840] = 16'b0000000000000000;
	sram_mem[78841] = 16'b0000000000000000;
	sram_mem[78842] = 16'b0000000000000000;
	sram_mem[78843] = 16'b0000000000000000;
	sram_mem[78844] = 16'b0000000000000000;
	sram_mem[78845] = 16'b0000000000000000;
	sram_mem[78846] = 16'b0000000000000000;
	sram_mem[78847] = 16'b0000000000000000;
	sram_mem[78848] = 16'b0000000000000000;
	sram_mem[78849] = 16'b0000000000000000;
	sram_mem[78850] = 16'b0000000000000000;
	sram_mem[78851] = 16'b0000000000000000;
	sram_mem[78852] = 16'b0000000000000000;
	sram_mem[78853] = 16'b0000000000000000;
	sram_mem[78854] = 16'b0000000000000000;
	sram_mem[78855] = 16'b0000000000000000;
	sram_mem[78856] = 16'b0000000000000000;
	sram_mem[78857] = 16'b0000000000000000;
	sram_mem[78858] = 16'b0000000000000000;
	sram_mem[78859] = 16'b0000000000000000;
	sram_mem[78860] = 16'b0000000000000000;
	sram_mem[78861] = 16'b0000000000000000;
	sram_mem[78862] = 16'b0000000000000000;
	sram_mem[78863] = 16'b0000000000000000;
	sram_mem[78864] = 16'b0000000000000000;
	sram_mem[78865] = 16'b0000000000000000;
	sram_mem[78866] = 16'b0000000000000000;
	sram_mem[78867] = 16'b0000000000000000;
	sram_mem[78868] = 16'b0000000000000000;
	sram_mem[78869] = 16'b0000000000000000;
	sram_mem[78870] = 16'b0000000000000000;
	sram_mem[78871] = 16'b0000000000000000;
	sram_mem[78872] = 16'b0000000000000000;
	sram_mem[78873] = 16'b0000000000000000;
	sram_mem[78874] = 16'b0000000000000000;
	sram_mem[78875] = 16'b0000000000000000;
	sram_mem[78876] = 16'b0000000000000000;
	sram_mem[78877] = 16'b0000000000000000;
	sram_mem[78878] = 16'b0000000000000000;
	sram_mem[78879] = 16'b0000000000000000;
	sram_mem[78880] = 16'b0000000000000000;
	sram_mem[78881] = 16'b0000000000000000;
	sram_mem[78882] = 16'b0000000000000000;
	sram_mem[78883] = 16'b0000000000000000;
	sram_mem[78884] = 16'b0000000000000000;
	sram_mem[78885] = 16'b0000000000000000;
	sram_mem[78886] = 16'b0000000000000000;
	sram_mem[78887] = 16'b0000000000000000;
	sram_mem[78888] = 16'b0000000000000000;
	sram_mem[78889] = 16'b0000000000000000;
	sram_mem[78890] = 16'b0000000000000000;
	sram_mem[78891] = 16'b0000000000000000;
	sram_mem[78892] = 16'b0000000000000000;
	sram_mem[78893] = 16'b0000000000000000;
	sram_mem[78894] = 16'b0000000000000000;
	sram_mem[78895] = 16'b0000000000000000;
	sram_mem[78896] = 16'b0000000000000000;
	sram_mem[78897] = 16'b0000000000000000;
	sram_mem[78898] = 16'b0000000000000000;
	sram_mem[78899] = 16'b0000000000000000;
	sram_mem[78900] = 16'b0000000000000000;
	sram_mem[78901] = 16'b0000000000000000;
	sram_mem[78902] = 16'b0000000000000000;
	sram_mem[78903] = 16'b0000000000000000;
	sram_mem[78904] = 16'b0000000000000000;
	sram_mem[78905] = 16'b0000000000000000;
	sram_mem[78906] = 16'b0000000000000000;
	sram_mem[78907] = 16'b0000000000000000;
	sram_mem[78908] = 16'b0000000000000000;
	sram_mem[78909] = 16'b0000000000000000;
	sram_mem[78910] = 16'b0000000000000000;
	sram_mem[78911] = 16'b0000000000000000;
	sram_mem[78912] = 16'b0000000000000000;
	sram_mem[78913] = 16'b0000000000000000;
	sram_mem[78914] = 16'b0000000000000000;
	sram_mem[78915] = 16'b0000000000000000;
	sram_mem[78916] = 16'b0000000000000000;
	sram_mem[78917] = 16'b0000000000000000;
	sram_mem[78918] = 16'b0000000000000000;
	sram_mem[78919] = 16'b0000000000000000;
	sram_mem[78920] = 16'b0000000000000000;
	sram_mem[78921] = 16'b0000000000000000;
	sram_mem[78922] = 16'b0000000000000000;
	sram_mem[78923] = 16'b0000000000000000;
	sram_mem[78924] = 16'b0000000000000000;
	sram_mem[78925] = 16'b0000000000000000;
	sram_mem[78926] = 16'b0000000000000000;
	sram_mem[78927] = 16'b0000000000000000;
	sram_mem[78928] = 16'b0000000000000000;
	sram_mem[78929] = 16'b0000000000000000;
	sram_mem[78930] = 16'b0000000000000000;
	sram_mem[78931] = 16'b0000000000000000;
	sram_mem[78932] = 16'b0000000000000000;
	sram_mem[78933] = 16'b0000000000000000;
	sram_mem[78934] = 16'b0000000000000000;
	sram_mem[78935] = 16'b0000000000000000;
	sram_mem[78936] = 16'b0000000000000000;
	sram_mem[78937] = 16'b0000000000000000;
	sram_mem[78938] = 16'b0000000000000000;
	sram_mem[78939] = 16'b0000000000000000;
	sram_mem[78940] = 16'b0000000000000000;
	sram_mem[78941] = 16'b0000000000000000;
	sram_mem[78942] = 16'b0000000000000000;
	sram_mem[78943] = 16'b0000000000000000;
	sram_mem[78944] = 16'b0000000000000000;
	sram_mem[78945] = 16'b0000000000000000;
	sram_mem[78946] = 16'b0000000000000000;
	sram_mem[78947] = 16'b0000000000000000;
	sram_mem[78948] = 16'b0000000000000000;
	sram_mem[78949] = 16'b0000000000000000;
	sram_mem[78950] = 16'b0000000000000000;
	sram_mem[78951] = 16'b0000000000000000;
	sram_mem[78952] = 16'b0000000000000000;
	sram_mem[78953] = 16'b0000000000000000;
	sram_mem[78954] = 16'b0000000000000000;
	sram_mem[78955] = 16'b0000000000000000;
	sram_mem[78956] = 16'b0000000000000000;
	sram_mem[78957] = 16'b0000000000000000;
	sram_mem[78958] = 16'b0000000000000000;
	sram_mem[78959] = 16'b0000000000000000;
	sram_mem[78960] = 16'b0000000000000000;
	sram_mem[78961] = 16'b0000000000000000;
	sram_mem[78962] = 16'b0000000000000000;
	sram_mem[78963] = 16'b0000000000000000;
	sram_mem[78964] = 16'b0000000000000000;
	sram_mem[78965] = 16'b0000000000000000;
	sram_mem[78966] = 16'b0000000000000000;
	sram_mem[78967] = 16'b0000000000000000;
	sram_mem[78968] = 16'b0000000000000000;
	sram_mem[78969] = 16'b0000000000000000;
	sram_mem[78970] = 16'b0000000000000000;
	sram_mem[78971] = 16'b0000000000000000;
	sram_mem[78972] = 16'b0000000000000000;
	sram_mem[78973] = 16'b0000000000000000;
	sram_mem[78974] = 16'b0000000000000000;
	sram_mem[78975] = 16'b0000000000000000;
	sram_mem[78976] = 16'b0000000000000000;
	sram_mem[78977] = 16'b0000000000000000;
	sram_mem[78978] = 16'b0000000000000000;
	sram_mem[78979] = 16'b0000000000000000;
	sram_mem[78980] = 16'b0000000000000000;
	sram_mem[78981] = 16'b0000000000000000;
	sram_mem[78982] = 16'b0000000000000000;
	sram_mem[78983] = 16'b0000000000000000;
	sram_mem[78984] = 16'b0000000000000000;
	sram_mem[78985] = 16'b0000000000000000;
	sram_mem[78986] = 16'b0000000000000000;
	sram_mem[78987] = 16'b0000000000000000;
	sram_mem[78988] = 16'b0000000000000000;
	sram_mem[78989] = 16'b0000000000000000;
	sram_mem[78990] = 16'b0000000000000000;
	sram_mem[78991] = 16'b0000000000000000;
	sram_mem[78992] = 16'b0000000000000000;
	sram_mem[78993] = 16'b0000000000000000;
	sram_mem[78994] = 16'b0000000000000000;
	sram_mem[78995] = 16'b0000000000000000;
	sram_mem[78996] = 16'b0000000000000000;
	sram_mem[78997] = 16'b0000000000000000;
	sram_mem[78998] = 16'b0000000000000000;
	sram_mem[78999] = 16'b0000000000000000;
	sram_mem[79000] = 16'b0000000000000000;
	sram_mem[79001] = 16'b0000000000000000;
	sram_mem[79002] = 16'b0000000000000000;
	sram_mem[79003] = 16'b0000000000000000;
	sram_mem[79004] = 16'b0000000000000000;
	sram_mem[79005] = 16'b0000000000000000;
	sram_mem[79006] = 16'b0000000000000000;
	sram_mem[79007] = 16'b0000000000000000;
	sram_mem[79008] = 16'b0000000000000000;
	sram_mem[79009] = 16'b0000000000000000;
	sram_mem[79010] = 16'b0000000000000000;
	sram_mem[79011] = 16'b0000000000000000;
	sram_mem[79012] = 16'b0000000000000000;
	sram_mem[79013] = 16'b0000000000000000;
	sram_mem[79014] = 16'b0000000000000000;
	sram_mem[79015] = 16'b0000000000000000;
	sram_mem[79016] = 16'b0000000000000000;
	sram_mem[79017] = 16'b0000000000000000;
	sram_mem[79018] = 16'b0000000000000000;
	sram_mem[79019] = 16'b0000000000000000;
	sram_mem[79020] = 16'b0000000000000000;
	sram_mem[79021] = 16'b0000000000000000;
	sram_mem[79022] = 16'b0000000000000000;
	sram_mem[79023] = 16'b0000000000000000;
	sram_mem[79024] = 16'b0000000000000000;
	sram_mem[79025] = 16'b0000000000000000;
	sram_mem[79026] = 16'b0000000000000000;
	sram_mem[79027] = 16'b0000000000000000;
	sram_mem[79028] = 16'b0000000000000000;
	sram_mem[79029] = 16'b0000000000000000;
	sram_mem[79030] = 16'b0000000000000000;
	sram_mem[79031] = 16'b0000000000000000;
	sram_mem[79032] = 16'b0000000000000000;
	sram_mem[79033] = 16'b0000000000000000;
	sram_mem[79034] = 16'b0000000000000000;
	sram_mem[79035] = 16'b0000000000000000;
	sram_mem[79036] = 16'b0000000000000000;
	sram_mem[79037] = 16'b0000000000000000;
	sram_mem[79038] = 16'b0000000000000000;
	sram_mem[79039] = 16'b0000000000000000;
	sram_mem[79040] = 16'b0000000000000000;
	sram_mem[79041] = 16'b0000000000000000;
	sram_mem[79042] = 16'b0000000000000000;
	sram_mem[79043] = 16'b0000000000000000;
	sram_mem[79044] = 16'b0000000000000000;
	sram_mem[79045] = 16'b0000000000000000;
	sram_mem[79046] = 16'b0000000000000000;
	sram_mem[79047] = 16'b0000000000000000;
	sram_mem[79048] = 16'b0000000000000000;
	sram_mem[79049] = 16'b0000000000000000;
	sram_mem[79050] = 16'b0000000000000000;
	sram_mem[79051] = 16'b0000000000000000;
	sram_mem[79052] = 16'b0000000000000000;
	sram_mem[79053] = 16'b0000000000000000;
	sram_mem[79054] = 16'b0000000000000000;
	sram_mem[79055] = 16'b0000000000000000;
	sram_mem[79056] = 16'b0000000000000000;
	sram_mem[79057] = 16'b0000000000000000;
	sram_mem[79058] = 16'b0000000000000000;
	sram_mem[79059] = 16'b0000000000000000;
	sram_mem[79060] = 16'b0000000000000000;
	sram_mem[79061] = 16'b0000000000000000;
	sram_mem[79062] = 16'b0000000000000000;
	sram_mem[79063] = 16'b0000000000000000;
	sram_mem[79064] = 16'b0000000000000000;
	sram_mem[79065] = 16'b0000000000000000;
	sram_mem[79066] = 16'b0000000000000000;
	sram_mem[79067] = 16'b0000000000000000;
	sram_mem[79068] = 16'b0000000000000000;
	sram_mem[79069] = 16'b0000000000000000;
	sram_mem[79070] = 16'b0000000000000000;
	sram_mem[79071] = 16'b0000000000000000;
	sram_mem[79072] = 16'b0000000000000000;
	sram_mem[79073] = 16'b0000000000000000;
	sram_mem[79074] = 16'b0000000000000000;
	sram_mem[79075] = 16'b0000000000000000;
	sram_mem[79076] = 16'b0000000000000000;
	sram_mem[79077] = 16'b0000000000000000;
	sram_mem[79078] = 16'b0000000000000000;
	sram_mem[79079] = 16'b0000000000000000;
	sram_mem[79080] = 16'b0000000000000000;
	sram_mem[79081] = 16'b0000000000000000;
	sram_mem[79082] = 16'b0000000000000000;
	sram_mem[79083] = 16'b0000000000000000;
	sram_mem[79084] = 16'b0000000000000000;
	sram_mem[79085] = 16'b0000000000000000;
	sram_mem[79086] = 16'b0000000000000000;
	sram_mem[79087] = 16'b0000000000000000;
	sram_mem[79088] = 16'b0000000000000000;
	sram_mem[79089] = 16'b0000000000000000;
	sram_mem[79090] = 16'b0000000000000000;
	sram_mem[79091] = 16'b0000000000000000;
	sram_mem[79092] = 16'b0000000000000000;
	sram_mem[79093] = 16'b0000000000000000;
	sram_mem[79094] = 16'b0000000000000000;
	sram_mem[79095] = 16'b0000000000000000;
	sram_mem[79096] = 16'b0000000000000000;
	sram_mem[79097] = 16'b0000000000000000;
	sram_mem[79098] = 16'b0000000000000000;
	sram_mem[79099] = 16'b0000000000000000;
	sram_mem[79100] = 16'b0000000000000000;
	sram_mem[79101] = 16'b0000000000000000;
	sram_mem[79102] = 16'b0000000000000000;
	sram_mem[79103] = 16'b0000000000000000;
	sram_mem[79104] = 16'b0000000000000000;
	sram_mem[79105] = 16'b0000000000000000;
	sram_mem[79106] = 16'b0000000000000000;
	sram_mem[79107] = 16'b0000000000000000;
	sram_mem[79108] = 16'b0000000000000000;
	sram_mem[79109] = 16'b0000000000000000;
	sram_mem[79110] = 16'b0000000000000000;
	sram_mem[79111] = 16'b0000000000000000;
	sram_mem[79112] = 16'b0000000000000000;
	sram_mem[79113] = 16'b0000000000000000;
	sram_mem[79114] = 16'b0000000000000000;
	sram_mem[79115] = 16'b0000000000000000;
	sram_mem[79116] = 16'b0000000000000000;
	sram_mem[79117] = 16'b0000000000000000;
	sram_mem[79118] = 16'b0000000000000000;
	sram_mem[79119] = 16'b0000000000000000;
	sram_mem[79120] = 16'b0000000000000000;
	sram_mem[79121] = 16'b0000000000000000;
	sram_mem[79122] = 16'b0000000000000000;
	sram_mem[79123] = 16'b0000000000000000;
	sram_mem[79124] = 16'b0000000000000000;
	sram_mem[79125] = 16'b0000000000000000;
	sram_mem[79126] = 16'b0000000000000000;
	sram_mem[79127] = 16'b0000000000000000;
	sram_mem[79128] = 16'b0000000000000000;
	sram_mem[79129] = 16'b0000000000000000;
	sram_mem[79130] = 16'b0000000000000000;
	sram_mem[79131] = 16'b0000000000000000;
	sram_mem[79132] = 16'b0000000000000000;
	sram_mem[79133] = 16'b0000000000000000;
	sram_mem[79134] = 16'b0000000000000000;
	sram_mem[79135] = 16'b0000000000000000;
	sram_mem[79136] = 16'b0000000000000000;
	sram_mem[79137] = 16'b0000000000000000;
	sram_mem[79138] = 16'b0000000000000000;
	sram_mem[79139] = 16'b0000000000000000;
	sram_mem[79140] = 16'b0000000000000000;
	sram_mem[79141] = 16'b0000000000000000;
	sram_mem[79142] = 16'b0000000000000000;
	sram_mem[79143] = 16'b0000000000000000;
	sram_mem[79144] = 16'b0000000000000000;
	sram_mem[79145] = 16'b0000000000000000;
	sram_mem[79146] = 16'b0000000000000000;
	sram_mem[79147] = 16'b0000000000000000;
	sram_mem[79148] = 16'b0000000000000000;
	sram_mem[79149] = 16'b0000000000000000;
	sram_mem[79150] = 16'b0000000000000000;
	sram_mem[79151] = 16'b0000000000000000;
	sram_mem[79152] = 16'b0000000000000000;
	sram_mem[79153] = 16'b0000000000000000;
	sram_mem[79154] = 16'b0000000000000000;
	sram_mem[79155] = 16'b0000000000000000;
	sram_mem[79156] = 16'b0000000000000000;
	sram_mem[79157] = 16'b0000000000000000;
	sram_mem[79158] = 16'b0000000000000000;
	sram_mem[79159] = 16'b0000000000000000;
	sram_mem[79160] = 16'b0000000000000000;
	sram_mem[79161] = 16'b0000000000000000;
	sram_mem[79162] = 16'b0000000000000000;
	sram_mem[79163] = 16'b0000000000000000;
	sram_mem[79164] = 16'b0000000000000000;
	sram_mem[79165] = 16'b0000000000000000;
	sram_mem[79166] = 16'b0000000000000000;
	sram_mem[79167] = 16'b0000000000000000;
	sram_mem[79168] = 16'b0000000000000000;
	sram_mem[79169] = 16'b0000000000000000;
	sram_mem[79170] = 16'b0000000000000000;
	sram_mem[79171] = 16'b0000000000000000;
	sram_mem[79172] = 16'b0000000000000000;
	sram_mem[79173] = 16'b0000000000000000;
	sram_mem[79174] = 16'b0000000000000000;
	sram_mem[79175] = 16'b0000000000000000;
	sram_mem[79176] = 16'b0000000000000000;
	sram_mem[79177] = 16'b0000000000000000;
	sram_mem[79178] = 16'b0000000000000000;
	sram_mem[79179] = 16'b0000000000000000;
	sram_mem[79180] = 16'b0000000000000000;
	sram_mem[79181] = 16'b0000000000000000;
	sram_mem[79182] = 16'b0000000000000000;
	sram_mem[79183] = 16'b0000000000000000;
	sram_mem[79184] = 16'b0000000000000000;
	sram_mem[79185] = 16'b0000000000000000;
	sram_mem[79186] = 16'b0000000000000000;
	sram_mem[79187] = 16'b0000000000000000;
	sram_mem[79188] = 16'b0000000000000000;
	sram_mem[79189] = 16'b0000000000000000;
	sram_mem[79190] = 16'b0000000000000000;
	sram_mem[79191] = 16'b0000000000000000;
	sram_mem[79192] = 16'b0000000000000000;
	sram_mem[79193] = 16'b0000000000000000;
	sram_mem[79194] = 16'b0000000000000000;
	sram_mem[79195] = 16'b0000000000000000;
	sram_mem[79196] = 16'b0000000000000000;
	sram_mem[79197] = 16'b0000000000000000;
	sram_mem[79198] = 16'b0000000000000000;
	sram_mem[79199] = 16'b0000000000000000;
	sram_mem[79200] = 16'b0000000000000000;
	sram_mem[79201] = 16'b0000000000000000;
	sram_mem[79202] = 16'b0000000000000000;
	sram_mem[79203] = 16'b0000000000000000;
	sram_mem[79204] = 16'b0000000000000000;
	sram_mem[79205] = 16'b0000000000000000;
	sram_mem[79206] = 16'b0000000000000000;
	sram_mem[79207] = 16'b0000000000000000;
	sram_mem[79208] = 16'b0000000000000000;
	sram_mem[79209] = 16'b0000000000000000;
	sram_mem[79210] = 16'b0000000000000000;
	sram_mem[79211] = 16'b0000000000000000;
	sram_mem[79212] = 16'b0000000000000000;
	sram_mem[79213] = 16'b0000000000000000;
	sram_mem[79214] = 16'b0000000000000000;
	sram_mem[79215] = 16'b0000000000000000;
	sram_mem[79216] = 16'b0000000000000000;
	sram_mem[79217] = 16'b0000000000000000;
	sram_mem[79218] = 16'b0000000000000000;
	sram_mem[79219] = 16'b0000000000000000;
	sram_mem[79220] = 16'b0000000000000000;
	sram_mem[79221] = 16'b0000000000000000;
	sram_mem[79222] = 16'b0000000000000000;
	sram_mem[79223] = 16'b0000000000000000;
	sram_mem[79224] = 16'b0000000000000000;
	sram_mem[79225] = 16'b0000000000000000;
	sram_mem[79226] = 16'b0000000000000000;
	sram_mem[79227] = 16'b0000000000000000;
	sram_mem[79228] = 16'b0000000000000000;
	sram_mem[79229] = 16'b0000000000000000;
	sram_mem[79230] = 16'b0000000000000000;
	sram_mem[79231] = 16'b0000000000000000;
	sram_mem[79232] = 16'b0000000000000000;
	sram_mem[79233] = 16'b0000000000000000;
	sram_mem[79234] = 16'b0000000000000000;
	sram_mem[79235] = 16'b0000000000000000;
	sram_mem[79236] = 16'b0000000000000000;
	sram_mem[79237] = 16'b0000000000000000;
	sram_mem[79238] = 16'b0000000000000000;
	sram_mem[79239] = 16'b0000000000000000;
	sram_mem[79240] = 16'b0000000000000000;
	sram_mem[79241] = 16'b0000000000000000;
	sram_mem[79242] = 16'b0000000000000000;
	sram_mem[79243] = 16'b0000000000000000;
	sram_mem[79244] = 16'b0000000000000000;
	sram_mem[79245] = 16'b0000000000000000;
	sram_mem[79246] = 16'b0000000000000000;
	sram_mem[79247] = 16'b0000000000000000;
	sram_mem[79248] = 16'b0000000000000000;
	sram_mem[79249] = 16'b0000000000000000;
	sram_mem[79250] = 16'b0000000000000000;
	sram_mem[79251] = 16'b0000000000000000;
	sram_mem[79252] = 16'b0000000000000000;
	sram_mem[79253] = 16'b0000000000000000;
	sram_mem[79254] = 16'b0000000000000000;
	sram_mem[79255] = 16'b0000000000000000;
	sram_mem[79256] = 16'b0000000000000000;
	sram_mem[79257] = 16'b0000000000000000;
	sram_mem[79258] = 16'b0000000000000000;
	sram_mem[79259] = 16'b0000000000000000;
	sram_mem[79260] = 16'b0000000000000000;
	sram_mem[79261] = 16'b0000000000000000;
	sram_mem[79262] = 16'b0000000000000000;
	sram_mem[79263] = 16'b0000000000000000;
	sram_mem[79264] = 16'b0000000000000000;
	sram_mem[79265] = 16'b0000000000000000;
	sram_mem[79266] = 16'b0000000000000000;
	sram_mem[79267] = 16'b0000000000000000;
	sram_mem[79268] = 16'b0000000000000000;
	sram_mem[79269] = 16'b0000000000000000;
	sram_mem[79270] = 16'b0000000000000000;
	sram_mem[79271] = 16'b0000000000000000;
	sram_mem[79272] = 16'b0000000000000000;
	sram_mem[79273] = 16'b0000000000000000;
	sram_mem[79274] = 16'b0000000000000000;
	sram_mem[79275] = 16'b0000000000000000;
	sram_mem[79276] = 16'b0000000000000000;
	sram_mem[79277] = 16'b0000000000000000;
	sram_mem[79278] = 16'b0000000000000000;
	sram_mem[79279] = 16'b0000000000000000;
	sram_mem[79280] = 16'b0000000000000000;
	sram_mem[79281] = 16'b0000000000000000;
	sram_mem[79282] = 16'b0000000000000000;
	sram_mem[79283] = 16'b0000000000000000;
	sram_mem[79284] = 16'b0000000000000000;
	sram_mem[79285] = 16'b0000000000000000;
	sram_mem[79286] = 16'b0000000000000000;
	sram_mem[79287] = 16'b0000000000000000;
	sram_mem[79288] = 16'b0000000000000000;
	sram_mem[79289] = 16'b0000000000000000;
	sram_mem[79290] = 16'b0000000000000000;
	sram_mem[79291] = 16'b0000000000000000;
	sram_mem[79292] = 16'b0000000000000000;
	sram_mem[79293] = 16'b0000000000000000;
	sram_mem[79294] = 16'b0000000000000000;
	sram_mem[79295] = 16'b0000000000000000;
	sram_mem[79296] = 16'b0000000000000000;
	sram_mem[79297] = 16'b0000000000000000;
	sram_mem[79298] = 16'b0000000000000000;
	sram_mem[79299] = 16'b0000000000000000;
	sram_mem[79300] = 16'b0000000000000000;
	sram_mem[79301] = 16'b0000000000000000;
	sram_mem[79302] = 16'b0000000000000000;
	sram_mem[79303] = 16'b0000000000000000;
	sram_mem[79304] = 16'b0000000000000000;
	sram_mem[79305] = 16'b0000000000000000;
	sram_mem[79306] = 16'b0000000000000000;
	sram_mem[79307] = 16'b0000000000000000;
	sram_mem[79308] = 16'b0000000000000000;
	sram_mem[79309] = 16'b0000000000000000;
	sram_mem[79310] = 16'b0000000000000000;
	sram_mem[79311] = 16'b0000000000000000;
	sram_mem[79312] = 16'b0000000000000000;
	sram_mem[79313] = 16'b0000000000000000;
	sram_mem[79314] = 16'b0000000000000000;
	sram_mem[79315] = 16'b0000000000000000;
	sram_mem[79316] = 16'b0000000000000000;
	sram_mem[79317] = 16'b0000000000000000;
	sram_mem[79318] = 16'b0000000000000000;
	sram_mem[79319] = 16'b0000000000000000;
	sram_mem[79320] = 16'b0000000000000000;
	sram_mem[79321] = 16'b0000000000000000;
	sram_mem[79322] = 16'b0000000000000000;
	sram_mem[79323] = 16'b0000000000000000;
	sram_mem[79324] = 16'b0000000000000000;
	sram_mem[79325] = 16'b0000000000000000;
	sram_mem[79326] = 16'b0000000000000000;
	sram_mem[79327] = 16'b0000000000000000;
	sram_mem[79328] = 16'b0000000000000000;
	sram_mem[79329] = 16'b0000000000000000;
	sram_mem[79330] = 16'b0000000000000000;
	sram_mem[79331] = 16'b0000000000000000;
	sram_mem[79332] = 16'b0000000000000000;
	sram_mem[79333] = 16'b0000000000000000;
	sram_mem[79334] = 16'b0000000000000000;
	sram_mem[79335] = 16'b0000000000000000;
	sram_mem[79336] = 16'b0000000000000000;
	sram_mem[79337] = 16'b0000000000000000;
	sram_mem[79338] = 16'b0000000000000000;
	sram_mem[79339] = 16'b0000000000000000;
	sram_mem[79340] = 16'b0000000000000000;
	sram_mem[79341] = 16'b0000000000000000;
	sram_mem[79342] = 16'b0000000000000000;
	sram_mem[79343] = 16'b0000000000000000;
	sram_mem[79344] = 16'b0000000000000000;
	sram_mem[79345] = 16'b0000000000000000;
	sram_mem[79346] = 16'b0000000000000000;
	sram_mem[79347] = 16'b0000000000000000;
	sram_mem[79348] = 16'b0000000000000000;
	sram_mem[79349] = 16'b0000000000000000;
	sram_mem[79350] = 16'b0000000000000000;
	sram_mem[79351] = 16'b0000000000000000;
	sram_mem[79352] = 16'b0000000000000000;
	sram_mem[79353] = 16'b0000000000000000;
	sram_mem[79354] = 16'b0000000000000000;
	sram_mem[79355] = 16'b0000000000000000;
	sram_mem[79356] = 16'b0000000000000000;
	sram_mem[79357] = 16'b0000000000000000;
	sram_mem[79358] = 16'b0000000000000000;
	sram_mem[79359] = 16'b0000000000000000;
	sram_mem[79360] = 16'b0000000000000000;
	sram_mem[79361] = 16'b0000000000000000;
	sram_mem[79362] = 16'b0000000000000000;
	sram_mem[79363] = 16'b0000000000000000;
	sram_mem[79364] = 16'b0000000000000000;
	sram_mem[79365] = 16'b0000000000000000;
	sram_mem[79366] = 16'b0000000000000000;
	sram_mem[79367] = 16'b0000000000000000;
	sram_mem[79368] = 16'b0000000000000000;
	sram_mem[79369] = 16'b0000000000000000;
	sram_mem[79370] = 16'b0000000000000000;
	sram_mem[79371] = 16'b0000000000000000;
	sram_mem[79372] = 16'b0000000000000000;
	sram_mem[79373] = 16'b0000000000000000;
	sram_mem[79374] = 16'b0000000000000000;
	sram_mem[79375] = 16'b0000000000000000;
	sram_mem[79376] = 16'b0000000000000000;
	sram_mem[79377] = 16'b0000000000000000;
	sram_mem[79378] = 16'b0000000000000000;
	sram_mem[79379] = 16'b0000000000000000;
	sram_mem[79380] = 16'b0000000000000000;
	sram_mem[79381] = 16'b0000000000000000;
	sram_mem[79382] = 16'b0000000000000000;
	sram_mem[79383] = 16'b0000000000000000;
	sram_mem[79384] = 16'b0000000000000000;
	sram_mem[79385] = 16'b0000000000000000;
	sram_mem[79386] = 16'b0000000000000000;
	sram_mem[79387] = 16'b0000000000000000;
	sram_mem[79388] = 16'b0000000000000000;
	sram_mem[79389] = 16'b0000000000000000;
	sram_mem[79390] = 16'b0000000000000000;
	sram_mem[79391] = 16'b0000000000000000;
	sram_mem[79392] = 16'b0000000000000000;
	sram_mem[79393] = 16'b0000000000000000;
	sram_mem[79394] = 16'b0000000000000000;
	sram_mem[79395] = 16'b0000000000000000;
	sram_mem[79396] = 16'b0000000000000000;
	sram_mem[79397] = 16'b0000000000000000;
	sram_mem[79398] = 16'b0000000000000000;
	sram_mem[79399] = 16'b0000000000000000;
	sram_mem[79400] = 16'b0000000000000000;
	sram_mem[79401] = 16'b0000000000000000;
	sram_mem[79402] = 16'b0000000000000000;
	sram_mem[79403] = 16'b0000000000000000;
	sram_mem[79404] = 16'b0000000000000000;
	sram_mem[79405] = 16'b0000000000000000;
	sram_mem[79406] = 16'b0000000000000000;
	sram_mem[79407] = 16'b0000000000000000;
	sram_mem[79408] = 16'b0000000000000000;
	sram_mem[79409] = 16'b0000000000000000;
	sram_mem[79410] = 16'b0000000000000000;
	sram_mem[79411] = 16'b0000000000000000;
	sram_mem[79412] = 16'b0000000000000000;
	sram_mem[79413] = 16'b0000000000000000;
	sram_mem[79414] = 16'b0000000000000000;
	sram_mem[79415] = 16'b0000000000000000;
	sram_mem[79416] = 16'b0000000000000000;
	sram_mem[79417] = 16'b0000000000000000;
	sram_mem[79418] = 16'b0000000000000000;
	sram_mem[79419] = 16'b0000000000000000;
	sram_mem[79420] = 16'b0000000000000000;
	sram_mem[79421] = 16'b0000000000000000;
	sram_mem[79422] = 16'b0000000000000000;
	sram_mem[79423] = 16'b0000000000000000;
	sram_mem[79424] = 16'b0000000000000000;
	sram_mem[79425] = 16'b0000000000000000;
	sram_mem[79426] = 16'b0000000000000000;
	sram_mem[79427] = 16'b0000000000000000;
	sram_mem[79428] = 16'b0000000000000000;
	sram_mem[79429] = 16'b0000000000000000;
	sram_mem[79430] = 16'b0000000000000000;
	sram_mem[79431] = 16'b0000000000000000;
	sram_mem[79432] = 16'b0000000000000000;
	sram_mem[79433] = 16'b0000000000000000;
	sram_mem[79434] = 16'b0000000000000000;
	sram_mem[79435] = 16'b0000000000000000;
	sram_mem[79436] = 16'b0000000000000000;
	sram_mem[79437] = 16'b0000000000000000;
	sram_mem[79438] = 16'b0000000000000000;
	sram_mem[79439] = 16'b0000000000000000;
	sram_mem[79440] = 16'b0000000000000000;
	sram_mem[79441] = 16'b0000000000000000;
	sram_mem[79442] = 16'b0000000000000000;
	sram_mem[79443] = 16'b0000000000000000;
	sram_mem[79444] = 16'b0000000000000000;
	sram_mem[79445] = 16'b0000000000000000;
	sram_mem[79446] = 16'b0000000000000000;
	sram_mem[79447] = 16'b0000000000000000;
	sram_mem[79448] = 16'b0000000000000000;
	sram_mem[79449] = 16'b0000000000000000;
	sram_mem[79450] = 16'b0000000000000000;
	sram_mem[79451] = 16'b0000000000000000;
	sram_mem[79452] = 16'b0000000000000000;
	sram_mem[79453] = 16'b0000000000000000;
	sram_mem[79454] = 16'b0000000000000000;
	sram_mem[79455] = 16'b0000000000000000;
	sram_mem[79456] = 16'b0000000000000000;
	sram_mem[79457] = 16'b0000000000000000;
	sram_mem[79458] = 16'b0000000000000000;
	sram_mem[79459] = 16'b0000000000000000;
	sram_mem[79460] = 16'b0000000000000000;
	sram_mem[79461] = 16'b0000000000000000;
	sram_mem[79462] = 16'b0000000000000000;
	sram_mem[79463] = 16'b0000000000000000;
	sram_mem[79464] = 16'b0000000000000000;
	sram_mem[79465] = 16'b0000000000000000;
	sram_mem[79466] = 16'b0000000000000000;
	sram_mem[79467] = 16'b0000000000000000;
	sram_mem[79468] = 16'b0000000000000000;
	sram_mem[79469] = 16'b0000000000000000;
	sram_mem[79470] = 16'b0000000000000000;
	sram_mem[79471] = 16'b0000000000000000;
	sram_mem[79472] = 16'b0000000000000000;
	sram_mem[79473] = 16'b0000000000000000;
	sram_mem[79474] = 16'b0000000000000000;
	sram_mem[79475] = 16'b0000000000000000;
	sram_mem[79476] = 16'b0000000000000000;
	sram_mem[79477] = 16'b0000000000000000;
	sram_mem[79478] = 16'b0000000000000000;
	sram_mem[79479] = 16'b0000000000000000;
	sram_mem[79480] = 16'b0000000000000000;
	sram_mem[79481] = 16'b0000000000000000;
	sram_mem[79482] = 16'b0000000000000000;
	sram_mem[79483] = 16'b0000000000000000;
	sram_mem[79484] = 16'b0000000000000000;
	sram_mem[79485] = 16'b0000000000000000;
	sram_mem[79486] = 16'b0000000000000000;
	sram_mem[79487] = 16'b0000000000000000;
	sram_mem[79488] = 16'b0000000000000000;
	sram_mem[79489] = 16'b0000000000000000;
	sram_mem[79490] = 16'b0000000000000000;
	sram_mem[79491] = 16'b0000000000000000;
	sram_mem[79492] = 16'b0000000000000000;
	sram_mem[79493] = 16'b0000000000000000;
	sram_mem[79494] = 16'b0000000000000000;
	sram_mem[79495] = 16'b0000000000000000;
	sram_mem[79496] = 16'b0000000000000000;
	sram_mem[79497] = 16'b0000000000000000;
	sram_mem[79498] = 16'b0000000000000000;
	sram_mem[79499] = 16'b0000000000000000;
	sram_mem[79500] = 16'b0000000000000000;
	sram_mem[79501] = 16'b0000000000000000;
	sram_mem[79502] = 16'b0000000000000000;
	sram_mem[79503] = 16'b0000000000000000;
	sram_mem[79504] = 16'b0000000000000000;
	sram_mem[79505] = 16'b0000000000000000;
	sram_mem[79506] = 16'b0000000000000000;
	sram_mem[79507] = 16'b0000000000000000;
	sram_mem[79508] = 16'b0000000000000000;
	sram_mem[79509] = 16'b0000000000000000;
	sram_mem[79510] = 16'b0000000000000000;
	sram_mem[79511] = 16'b0000000000000000;
	sram_mem[79512] = 16'b0000000000000000;
	sram_mem[79513] = 16'b0000000000000000;
	sram_mem[79514] = 16'b0000000000000000;
	sram_mem[79515] = 16'b0000000000000000;
	sram_mem[79516] = 16'b0000000000000000;
	sram_mem[79517] = 16'b0000000000000000;
	sram_mem[79518] = 16'b0000000000000000;
	sram_mem[79519] = 16'b0000000000000000;
	sram_mem[79520] = 16'b0000000000000000;
	sram_mem[79521] = 16'b0000000000000000;
	sram_mem[79522] = 16'b0000000000000000;
	sram_mem[79523] = 16'b0000000000000000;
	sram_mem[79524] = 16'b0000000000000000;
	sram_mem[79525] = 16'b0000000000000000;
	sram_mem[79526] = 16'b0000000000000000;
	sram_mem[79527] = 16'b0000000000000000;
	sram_mem[79528] = 16'b0000000000000000;
	sram_mem[79529] = 16'b0000000000000000;
	sram_mem[79530] = 16'b0000000000000000;
	sram_mem[79531] = 16'b0000000000000000;
	sram_mem[79532] = 16'b0000000000000000;
	sram_mem[79533] = 16'b0000000000000000;
	sram_mem[79534] = 16'b0000000000000000;
	sram_mem[79535] = 16'b0000000000000000;
	sram_mem[79536] = 16'b0000000000000000;
	sram_mem[79537] = 16'b0000000000000000;
	sram_mem[79538] = 16'b0000000000000000;
	sram_mem[79539] = 16'b0000000000000000;
	sram_mem[79540] = 16'b0000000000000000;
	sram_mem[79541] = 16'b0000000000000000;
	sram_mem[79542] = 16'b0000000000000000;
	sram_mem[79543] = 16'b0000000000000000;
	sram_mem[79544] = 16'b0000000000000000;
	sram_mem[79545] = 16'b0000000000000000;
	sram_mem[79546] = 16'b0000000000000000;
	sram_mem[79547] = 16'b0000000000000000;
	sram_mem[79548] = 16'b0000000000000000;
	sram_mem[79549] = 16'b0000000000000000;
	sram_mem[79550] = 16'b0000000000000000;
	sram_mem[79551] = 16'b0000000000000000;
	sram_mem[79552] = 16'b0000000000000000;
	sram_mem[79553] = 16'b0000000000000000;
	sram_mem[79554] = 16'b0000000000000000;
	sram_mem[79555] = 16'b0000000000000000;
	sram_mem[79556] = 16'b0000000000000000;
	sram_mem[79557] = 16'b0000000000000000;
	sram_mem[79558] = 16'b0000000000000000;
	sram_mem[79559] = 16'b0000000000000000;
	sram_mem[79560] = 16'b0000000000000000;
	sram_mem[79561] = 16'b0000000000000000;
	sram_mem[79562] = 16'b0000000000000000;
	sram_mem[79563] = 16'b0000000000000000;
	sram_mem[79564] = 16'b0000000000000000;
	sram_mem[79565] = 16'b0000000000000000;
	sram_mem[79566] = 16'b0000000000000000;
	sram_mem[79567] = 16'b0000000000000000;
	sram_mem[79568] = 16'b0000000000000000;
	sram_mem[79569] = 16'b0000000000000000;
	sram_mem[79570] = 16'b0000000000000000;
	sram_mem[79571] = 16'b0000000000000000;
	sram_mem[79572] = 16'b0000000000000000;
	sram_mem[79573] = 16'b0000000000000000;
	sram_mem[79574] = 16'b0000000000000000;
	sram_mem[79575] = 16'b0000000000000000;
	sram_mem[79576] = 16'b0000000000000000;
	sram_mem[79577] = 16'b0000000000000000;
	sram_mem[79578] = 16'b0000000000000000;
	sram_mem[79579] = 16'b0000000000000000;
	sram_mem[79580] = 16'b0000000000000000;
	sram_mem[79581] = 16'b0000000000000000;
	sram_mem[79582] = 16'b0000000000000000;
	sram_mem[79583] = 16'b0000000000000000;
	sram_mem[79584] = 16'b0000000000000000;
	sram_mem[79585] = 16'b0000000000000000;
	sram_mem[79586] = 16'b0000000000000000;
	sram_mem[79587] = 16'b0000000000000000;
	sram_mem[79588] = 16'b0000000000000000;
	sram_mem[79589] = 16'b0000000000000000;
	sram_mem[79590] = 16'b0000000000000000;
	sram_mem[79591] = 16'b0000000000000000;
	sram_mem[79592] = 16'b0000000000000000;
	sram_mem[79593] = 16'b0000000000000000;
	sram_mem[79594] = 16'b0000000000000000;
	sram_mem[79595] = 16'b0000000000000000;
	sram_mem[79596] = 16'b0000000000000000;
	sram_mem[79597] = 16'b0000000000000000;
	sram_mem[79598] = 16'b0000000000000000;
	sram_mem[79599] = 16'b0000000000000000;
	sram_mem[79600] = 16'b0000000000000000;
	sram_mem[79601] = 16'b0000000000000000;
	sram_mem[79602] = 16'b0000000000000000;
	sram_mem[79603] = 16'b0000000000000000;
	sram_mem[79604] = 16'b0000000000000000;
	sram_mem[79605] = 16'b0000000000000000;
	sram_mem[79606] = 16'b0000000000000000;
	sram_mem[79607] = 16'b0000000000000000;
	sram_mem[79608] = 16'b0000000000000000;
	sram_mem[79609] = 16'b0000000000000000;
	sram_mem[79610] = 16'b0000000000000000;
	sram_mem[79611] = 16'b0000000000000000;
	sram_mem[79612] = 16'b0000000000000000;
	sram_mem[79613] = 16'b0000000000000000;
	sram_mem[79614] = 16'b0000000000000000;
	sram_mem[79615] = 16'b0000000000000000;
	sram_mem[79616] = 16'b0000000000000000;
	sram_mem[79617] = 16'b0000000000000000;
	sram_mem[79618] = 16'b0000000000000000;
	sram_mem[79619] = 16'b0000000000000000;
	sram_mem[79620] = 16'b0000000000000000;
	sram_mem[79621] = 16'b0000000000000000;
	sram_mem[79622] = 16'b0000000000000000;
	sram_mem[79623] = 16'b0000000000000000;
	sram_mem[79624] = 16'b0000000000000000;
	sram_mem[79625] = 16'b0000000000000000;
	sram_mem[79626] = 16'b0000000000000000;
	sram_mem[79627] = 16'b0000000000000000;
	sram_mem[79628] = 16'b0000000000000000;
	sram_mem[79629] = 16'b0000000000000000;
	sram_mem[79630] = 16'b0000000000000000;
	sram_mem[79631] = 16'b0000000000000000;
	sram_mem[79632] = 16'b0000000000000000;
	sram_mem[79633] = 16'b0000000000000000;
	sram_mem[79634] = 16'b0000000000000000;
	sram_mem[79635] = 16'b0000000000000000;
	sram_mem[79636] = 16'b0000000000000000;
	sram_mem[79637] = 16'b0000000000000000;
	sram_mem[79638] = 16'b0000000000000000;
	sram_mem[79639] = 16'b0000000000000000;
	sram_mem[79640] = 16'b0000000000000000;
	sram_mem[79641] = 16'b0000000000000000;
	sram_mem[79642] = 16'b0000000000000000;
	sram_mem[79643] = 16'b0000000000000000;
	sram_mem[79644] = 16'b0000000000000000;
	sram_mem[79645] = 16'b0000000000000000;
	sram_mem[79646] = 16'b0000000000000000;
	sram_mem[79647] = 16'b0000000000000000;
	sram_mem[79648] = 16'b0000000000000000;
	sram_mem[79649] = 16'b0000000000000000;
	sram_mem[79650] = 16'b0000000000000000;
	sram_mem[79651] = 16'b0000000000000000;
	sram_mem[79652] = 16'b0000000000000000;
	sram_mem[79653] = 16'b0000000000000000;
	sram_mem[79654] = 16'b0000000000000000;
	sram_mem[79655] = 16'b0000000000000000;
	sram_mem[79656] = 16'b0000000000000000;
	sram_mem[79657] = 16'b0000000000000000;
	sram_mem[79658] = 16'b0000000000000000;
	sram_mem[79659] = 16'b0000000000000000;
	sram_mem[79660] = 16'b0000000000000000;
	sram_mem[79661] = 16'b0000000000000000;
	sram_mem[79662] = 16'b0000000000000000;
	sram_mem[79663] = 16'b0000000000000000;
	sram_mem[79664] = 16'b0000000000000000;
	sram_mem[79665] = 16'b0000000000000000;
	sram_mem[79666] = 16'b0000000000000000;
	sram_mem[79667] = 16'b0000000000000000;
	sram_mem[79668] = 16'b0000000000000000;
	sram_mem[79669] = 16'b0000000000000000;
	sram_mem[79670] = 16'b0000000000000000;
	sram_mem[79671] = 16'b0000000000000000;
	sram_mem[79672] = 16'b0000000000000000;
	sram_mem[79673] = 16'b0000000000000000;
	sram_mem[79674] = 16'b0000000000000000;
	sram_mem[79675] = 16'b0000000000000000;
	sram_mem[79676] = 16'b0000000000000000;
	sram_mem[79677] = 16'b0000000000000000;
	sram_mem[79678] = 16'b0000000000000000;
	sram_mem[79679] = 16'b0000000000000000;
	sram_mem[79680] = 16'b0000000000000000;
	sram_mem[79681] = 16'b0000000000000000;
	sram_mem[79682] = 16'b0000000000000000;
	sram_mem[79683] = 16'b0000000000000000;
	sram_mem[79684] = 16'b0000000000000000;
	sram_mem[79685] = 16'b0000000000000000;
	sram_mem[79686] = 16'b0000000000000000;
	sram_mem[79687] = 16'b0000000000000000;
	sram_mem[79688] = 16'b0000000000000000;
	sram_mem[79689] = 16'b0000000000000000;
	sram_mem[79690] = 16'b0000000000000000;
	sram_mem[79691] = 16'b0000000000000000;
	sram_mem[79692] = 16'b0000000000000000;
	sram_mem[79693] = 16'b0000000000000000;
	sram_mem[79694] = 16'b0000000000000000;
	sram_mem[79695] = 16'b0000000000000000;
	sram_mem[79696] = 16'b0000000000000000;
	sram_mem[79697] = 16'b0000000000000000;
	sram_mem[79698] = 16'b0000000000000000;
	sram_mem[79699] = 16'b0000000000000000;
	sram_mem[79700] = 16'b0000000000000000;
	sram_mem[79701] = 16'b0000000000000000;
	sram_mem[79702] = 16'b0000000000000000;
	sram_mem[79703] = 16'b0000000000000000;
	sram_mem[79704] = 16'b0000000000000000;
	sram_mem[79705] = 16'b0000000000000000;
	sram_mem[79706] = 16'b0000000000000000;
	sram_mem[79707] = 16'b0000000000000000;
	sram_mem[79708] = 16'b0000000000000000;
	sram_mem[79709] = 16'b0000000000000000;
	sram_mem[79710] = 16'b0000000000000000;
	sram_mem[79711] = 16'b0000000000000000;
	sram_mem[79712] = 16'b0000000000000000;
	sram_mem[79713] = 16'b0000000000000000;
	sram_mem[79714] = 16'b0000000000000000;
	sram_mem[79715] = 16'b0000000000000000;
	sram_mem[79716] = 16'b0000000000000000;
	sram_mem[79717] = 16'b0000000000000000;
	sram_mem[79718] = 16'b0000000000000000;
	sram_mem[79719] = 16'b0000000000000000;
	sram_mem[79720] = 16'b0000000000000000;
	sram_mem[79721] = 16'b0000000000000000;
	sram_mem[79722] = 16'b0000000000000000;
	sram_mem[79723] = 16'b0000000000000000;
	sram_mem[79724] = 16'b0000000000000000;
	sram_mem[79725] = 16'b0000000000000000;
	sram_mem[79726] = 16'b0000000000000000;
	sram_mem[79727] = 16'b0000000000000000;
	sram_mem[79728] = 16'b0000000000000000;
	sram_mem[79729] = 16'b0000000000000000;
	sram_mem[79730] = 16'b0000000000000000;
	sram_mem[79731] = 16'b0000000000000000;
	sram_mem[79732] = 16'b0000000000000000;
	sram_mem[79733] = 16'b0000000000000000;
	sram_mem[79734] = 16'b0000000000000000;
	sram_mem[79735] = 16'b0000000000000000;
	sram_mem[79736] = 16'b0000000000000000;
	sram_mem[79737] = 16'b0000000000000000;
	sram_mem[79738] = 16'b0000000000000000;
	sram_mem[79739] = 16'b0000000000000000;
	sram_mem[79740] = 16'b0000000000000000;
	sram_mem[79741] = 16'b0000000000000000;
	sram_mem[79742] = 16'b0000000000000000;
	sram_mem[79743] = 16'b0000000000000000;
	sram_mem[79744] = 16'b0000000000000000;
	sram_mem[79745] = 16'b0000000000000000;
	sram_mem[79746] = 16'b0000000000000000;
	sram_mem[79747] = 16'b0000000000000000;
	sram_mem[79748] = 16'b0000000000000000;
	sram_mem[79749] = 16'b0000000000000000;
	sram_mem[79750] = 16'b0000000000000000;
	sram_mem[79751] = 16'b0000000000000000;
	sram_mem[79752] = 16'b0000000000000000;
	sram_mem[79753] = 16'b0000000000000000;
	sram_mem[79754] = 16'b0000000000000000;
	sram_mem[79755] = 16'b0000000000000000;
	sram_mem[79756] = 16'b0000000000000000;
	sram_mem[79757] = 16'b0000000000000000;
	sram_mem[79758] = 16'b0000000000000000;
	sram_mem[79759] = 16'b0000000000000000;
	sram_mem[79760] = 16'b0000000000000000;
	sram_mem[79761] = 16'b0000000000000000;
	sram_mem[79762] = 16'b0000000000000000;
	sram_mem[79763] = 16'b0000000000000000;
	sram_mem[79764] = 16'b0000000000000000;
	sram_mem[79765] = 16'b0000000000000000;
	sram_mem[79766] = 16'b0000000000000000;
	sram_mem[79767] = 16'b0000000000000000;
	sram_mem[79768] = 16'b0000000000000000;
	sram_mem[79769] = 16'b0000000000000000;
	sram_mem[79770] = 16'b0000000000000000;
	sram_mem[79771] = 16'b0000000000000000;
	sram_mem[79772] = 16'b0000000000000000;
	sram_mem[79773] = 16'b0000000000000000;
	sram_mem[79774] = 16'b0000000000000000;
	sram_mem[79775] = 16'b0000000000000000;
	sram_mem[79776] = 16'b0000000000000000;
	sram_mem[79777] = 16'b0000000000000000;
	sram_mem[79778] = 16'b0000000000000000;
	sram_mem[79779] = 16'b0000000000000000;
	sram_mem[79780] = 16'b0000000000000000;
	sram_mem[79781] = 16'b0000000000000000;
	sram_mem[79782] = 16'b0000000000000000;
	sram_mem[79783] = 16'b0000000000000000;
	sram_mem[79784] = 16'b0000000000000000;
	sram_mem[79785] = 16'b0000000000000000;
	sram_mem[79786] = 16'b0000000000000000;
	sram_mem[79787] = 16'b0000000000000000;
	sram_mem[79788] = 16'b0000000000000000;
	sram_mem[79789] = 16'b0000000000000000;
	sram_mem[79790] = 16'b0000000000000000;
	sram_mem[79791] = 16'b0000000000000000;
	sram_mem[79792] = 16'b0000000000000000;
	sram_mem[79793] = 16'b0000000000000000;
	sram_mem[79794] = 16'b0000000000000000;
	sram_mem[79795] = 16'b0000000000000000;
	sram_mem[79796] = 16'b0000000000000000;
	sram_mem[79797] = 16'b0000000000000000;
	sram_mem[79798] = 16'b0000000000000000;
	sram_mem[79799] = 16'b0000000000000000;
	sram_mem[79800] = 16'b0000000000000000;
	sram_mem[79801] = 16'b0000000000000000;
	sram_mem[79802] = 16'b0000000000000000;
	sram_mem[79803] = 16'b0000000000000000;
	sram_mem[79804] = 16'b0000000000000000;
	sram_mem[79805] = 16'b0000000000000000;
	sram_mem[79806] = 16'b0000000000000000;
	sram_mem[79807] = 16'b0000000000000000;
	sram_mem[79808] = 16'b0000000000000000;
	sram_mem[79809] = 16'b0000000000000000;
	sram_mem[79810] = 16'b0000000000000000;
	sram_mem[79811] = 16'b0000000000000000;
	sram_mem[79812] = 16'b0000000000000000;
	sram_mem[79813] = 16'b0000000000000000;
	sram_mem[79814] = 16'b0000000000000000;
	sram_mem[79815] = 16'b0000000000000000;
	sram_mem[79816] = 16'b0000000000000000;
	sram_mem[79817] = 16'b0000000000000000;
	sram_mem[79818] = 16'b0000000000000000;
	sram_mem[79819] = 16'b0000000000000000;
	sram_mem[79820] = 16'b0000000000000000;
	sram_mem[79821] = 16'b0000000000000000;
	sram_mem[79822] = 16'b0000000000000000;
	sram_mem[79823] = 16'b0000000000000000;
	sram_mem[79824] = 16'b0000000000000000;
	sram_mem[79825] = 16'b0000000000000000;
	sram_mem[79826] = 16'b0000000000000000;
	sram_mem[79827] = 16'b0000000000000000;
	sram_mem[79828] = 16'b0000000000000000;
	sram_mem[79829] = 16'b0000000000000000;
	sram_mem[79830] = 16'b0000000000000000;
	sram_mem[79831] = 16'b0000000000000000;
	sram_mem[79832] = 16'b0000000000000000;
	sram_mem[79833] = 16'b0000000000000000;
	sram_mem[79834] = 16'b0000000000000000;
	sram_mem[79835] = 16'b0000000000000000;
	sram_mem[79836] = 16'b0000000000000000;
	sram_mem[79837] = 16'b0000000000000000;
	sram_mem[79838] = 16'b0000000000000000;
	sram_mem[79839] = 16'b0000000000000000;
	sram_mem[79840] = 16'b0000000000000000;
	sram_mem[79841] = 16'b0000000000000000;
	sram_mem[79842] = 16'b0000000000000000;
	sram_mem[79843] = 16'b0000000000000000;
	sram_mem[79844] = 16'b0000000000000000;
	sram_mem[79845] = 16'b0000000000000000;
	sram_mem[79846] = 16'b0000000000000000;
	sram_mem[79847] = 16'b0000000000000000;
	sram_mem[79848] = 16'b0000000000000000;
	sram_mem[79849] = 16'b0000000000000000;
	sram_mem[79850] = 16'b0000000000000000;
	sram_mem[79851] = 16'b0000000000000000;
	sram_mem[79852] = 16'b0000000000000000;
	sram_mem[79853] = 16'b0000000000000000;
	sram_mem[79854] = 16'b0000000000000000;
	sram_mem[79855] = 16'b0000000000000000;
	sram_mem[79856] = 16'b0000000000000000;
	sram_mem[79857] = 16'b0000000000000000;
	sram_mem[79858] = 16'b0000000000000000;
	sram_mem[79859] = 16'b0000000000000000;
	sram_mem[79860] = 16'b0000000000000000;
	sram_mem[79861] = 16'b0000000000000000;
	sram_mem[79862] = 16'b0000000000000000;
	sram_mem[79863] = 16'b0000000000000000;
	sram_mem[79864] = 16'b0000000000000000;
	sram_mem[79865] = 16'b0000000000000000;
	sram_mem[79866] = 16'b0000000000000000;
	sram_mem[79867] = 16'b0000000000000000;
	sram_mem[79868] = 16'b0000000000000000;
	sram_mem[79869] = 16'b0000000000000000;
	sram_mem[79870] = 16'b0000000000000000;
	sram_mem[79871] = 16'b0000000000000000;
	sram_mem[79872] = 16'b0000000000000000;
	sram_mem[79873] = 16'b0000000000000000;
	sram_mem[79874] = 16'b0000000000000000;
	sram_mem[79875] = 16'b0000000000000000;
	sram_mem[79876] = 16'b0000000000000000;
	sram_mem[79877] = 16'b0000000000000000;
	sram_mem[79878] = 16'b0000000000000000;
	sram_mem[79879] = 16'b0000000000000000;
	sram_mem[79880] = 16'b0000000000000000;
	sram_mem[79881] = 16'b0000000000000000;
	sram_mem[79882] = 16'b0000000000000000;
	sram_mem[79883] = 16'b0000000000000000;
	sram_mem[79884] = 16'b0000000000000000;
	sram_mem[79885] = 16'b0000000000000000;
	sram_mem[79886] = 16'b0000000000000000;
	sram_mem[79887] = 16'b0000000000000000;
	sram_mem[79888] = 16'b0000000000000000;
	sram_mem[79889] = 16'b0000000000000000;
	sram_mem[79890] = 16'b0000000000000000;
	sram_mem[79891] = 16'b0000000000000000;
	sram_mem[79892] = 16'b0000000000000000;
	sram_mem[79893] = 16'b0000000000000000;
	sram_mem[79894] = 16'b0000000000000000;
	sram_mem[79895] = 16'b0000000000000000;
	sram_mem[79896] = 16'b0000000000000000;
	sram_mem[79897] = 16'b0000000000000000;
	sram_mem[79898] = 16'b0000000000000000;
	sram_mem[79899] = 16'b0000000000000000;
	sram_mem[79900] = 16'b0000000000000000;
	sram_mem[79901] = 16'b0000000000000000;
	sram_mem[79902] = 16'b0000000000000000;
	sram_mem[79903] = 16'b0000000000000000;
	sram_mem[79904] = 16'b0000000000000000;
	sram_mem[79905] = 16'b0000000000000000;
	sram_mem[79906] = 16'b0000000000000000;
	sram_mem[79907] = 16'b0000000000000000;
	sram_mem[79908] = 16'b0000000000000000;
	sram_mem[79909] = 16'b0000000000000000;
	sram_mem[79910] = 16'b0000000000000000;
	sram_mem[79911] = 16'b0000000000000000;
	sram_mem[79912] = 16'b0000000000000000;
	sram_mem[79913] = 16'b0000000000000000;
	sram_mem[79914] = 16'b0000000000000000;
	sram_mem[79915] = 16'b0000000000000000;
	sram_mem[79916] = 16'b0000000000000000;
	sram_mem[79917] = 16'b0000000000000000;
	sram_mem[79918] = 16'b0000000000000000;
	sram_mem[79919] = 16'b0000000000000000;
	sram_mem[79920] = 16'b0000000000000000;
	sram_mem[79921] = 16'b0000000000000000;
	sram_mem[79922] = 16'b0000000000000000;
	sram_mem[79923] = 16'b0000000000000000;
	sram_mem[79924] = 16'b0000000000000000;
	sram_mem[79925] = 16'b0000000000000000;
	sram_mem[79926] = 16'b0000000000000000;
	sram_mem[79927] = 16'b0000000000000000;
	sram_mem[79928] = 16'b0000000000000000;
	sram_mem[79929] = 16'b0000000000000000;
	sram_mem[79930] = 16'b0000000000000000;
	sram_mem[79931] = 16'b0000000000000000;
	sram_mem[79932] = 16'b0000000000000000;
	sram_mem[79933] = 16'b0000000000000000;
	sram_mem[79934] = 16'b0000000000000000;
	sram_mem[79935] = 16'b0000000000000000;
	sram_mem[79936] = 16'b0000000000000000;
	sram_mem[79937] = 16'b0000000000000000;
	sram_mem[79938] = 16'b0000000000000000;
	sram_mem[79939] = 16'b0000000000000000;
	sram_mem[79940] = 16'b0000000000000000;
	sram_mem[79941] = 16'b0000000000000000;
	sram_mem[79942] = 16'b0000000000000000;
	sram_mem[79943] = 16'b0000000000000000;
	sram_mem[79944] = 16'b0000000000000000;
	sram_mem[79945] = 16'b0000000000000000;
	sram_mem[79946] = 16'b0000000000000000;
	sram_mem[79947] = 16'b0000000000000000;
	sram_mem[79948] = 16'b0000000000000000;
	sram_mem[79949] = 16'b0000000000000000;
	sram_mem[79950] = 16'b0000000000000000;
	sram_mem[79951] = 16'b0000000000000000;
	sram_mem[79952] = 16'b0000000000000000;
	sram_mem[79953] = 16'b0000000000000000;
	sram_mem[79954] = 16'b0000000000000000;
	sram_mem[79955] = 16'b0000000000000000;
	sram_mem[79956] = 16'b0000000000000000;
	sram_mem[79957] = 16'b0000000000000000;
	sram_mem[79958] = 16'b0000000000000000;
	sram_mem[79959] = 16'b0000000000000000;
	sram_mem[79960] = 16'b0000000000000000;
	sram_mem[79961] = 16'b0000000000000000;
	sram_mem[79962] = 16'b0000000000000000;
	sram_mem[79963] = 16'b0000000000000000;
	sram_mem[79964] = 16'b0000000000000000;
	sram_mem[79965] = 16'b0000000000000000;
	sram_mem[79966] = 16'b0000000000000000;
	sram_mem[79967] = 16'b0000000000000000;
	sram_mem[79968] = 16'b0000000000000000;
	sram_mem[79969] = 16'b0000000000000000;
	sram_mem[79970] = 16'b0000000000000000;
	sram_mem[79971] = 16'b0000000000000000;
	sram_mem[79972] = 16'b0000000000000000;
	sram_mem[79973] = 16'b0000000000000000;
	sram_mem[79974] = 16'b0000000000000000;
	sram_mem[79975] = 16'b0000000000000000;
	sram_mem[79976] = 16'b0000000000000000;
	sram_mem[79977] = 16'b0000000000000000;
	sram_mem[79978] = 16'b0000000000000000;
	sram_mem[79979] = 16'b0000000000000000;
	sram_mem[79980] = 16'b0000000000000000;
	sram_mem[79981] = 16'b0000000000000000;
	sram_mem[79982] = 16'b0000000000000000;
	sram_mem[79983] = 16'b0000000000000000;
	sram_mem[79984] = 16'b0000000000000000;
	sram_mem[79985] = 16'b0000000000000000;
	sram_mem[79986] = 16'b0000000000000000;
	sram_mem[79987] = 16'b0000000000000000;
	sram_mem[79988] = 16'b0000000000000000;
	sram_mem[79989] = 16'b0000000000000000;
	sram_mem[79990] = 16'b0000000000000000;
	sram_mem[79991] = 16'b0000000000000000;
	sram_mem[79992] = 16'b0000000000000000;
	sram_mem[79993] = 16'b0000000000000000;
	sram_mem[79994] = 16'b0000000000000000;
	sram_mem[79995] = 16'b0000000000000000;
	sram_mem[79996] = 16'b0000000000000000;
	sram_mem[79997] = 16'b0000000000000000;
	sram_mem[79998] = 16'b0000000000000000;
	sram_mem[79999] = 16'b0000000000000000;
	sram_mem[80000] = 16'b0000000000000000;
	sram_mem[80001] = 16'b0000000000000000;
	sram_mem[80002] = 16'b0000000000000000;
	sram_mem[80003] = 16'b0000000000000000;
	sram_mem[80004] = 16'b0000000000000000;
	sram_mem[80005] = 16'b0000000000000000;
	sram_mem[80006] = 16'b0000000000000000;
	sram_mem[80007] = 16'b0000000000000000;
	sram_mem[80008] = 16'b0000000000000000;
	sram_mem[80009] = 16'b0000000000000000;
	sram_mem[80010] = 16'b0000000000000000;
	sram_mem[80011] = 16'b0000000000000000;
	sram_mem[80012] = 16'b0000000000000000;
	sram_mem[80013] = 16'b0000000000000000;
	sram_mem[80014] = 16'b0000000000000000;
	sram_mem[80015] = 16'b0000000000000000;
	sram_mem[80016] = 16'b0000000000000000;
	sram_mem[80017] = 16'b0000000000000000;
	sram_mem[80018] = 16'b0000000000000000;
	sram_mem[80019] = 16'b0000000000000000;
	sram_mem[80020] = 16'b0000000000000000;
	sram_mem[80021] = 16'b0000000000000000;
	sram_mem[80022] = 16'b0000000000000000;
	sram_mem[80023] = 16'b0000000000000000;
	sram_mem[80024] = 16'b0000000000000000;
	sram_mem[80025] = 16'b0000000000000000;
	sram_mem[80026] = 16'b0000000000000000;
	sram_mem[80027] = 16'b0000000000000000;
	sram_mem[80028] = 16'b0000000000000000;
	sram_mem[80029] = 16'b0000000000000000;
	sram_mem[80030] = 16'b0000000000000000;
	sram_mem[80031] = 16'b0000000000000000;
	sram_mem[80032] = 16'b0000000000000000;
	sram_mem[80033] = 16'b0000000000000000;
	sram_mem[80034] = 16'b0000000000000000;
	sram_mem[80035] = 16'b0000000000000000;
	sram_mem[80036] = 16'b0000000000000000;
	sram_mem[80037] = 16'b0000000000000000;
	sram_mem[80038] = 16'b0000000000000000;
	sram_mem[80039] = 16'b0000000000000000;
	sram_mem[80040] = 16'b0000000000000000;
	sram_mem[80041] = 16'b0000000000000000;
	sram_mem[80042] = 16'b0000000000000000;
	sram_mem[80043] = 16'b0000000000000000;
	sram_mem[80044] = 16'b0000000000000000;
	sram_mem[80045] = 16'b0000000000000000;
	sram_mem[80046] = 16'b0000000000000000;
	sram_mem[80047] = 16'b0000000000000000;
	sram_mem[80048] = 16'b0000000000000000;
	sram_mem[80049] = 16'b0000000000000000;
	sram_mem[80050] = 16'b0000000000000000;
	sram_mem[80051] = 16'b0000000000000000;
	sram_mem[80052] = 16'b0000000000000000;
	sram_mem[80053] = 16'b0000000000000000;
	sram_mem[80054] = 16'b0000000000000000;
	sram_mem[80055] = 16'b0000000000000000;
	sram_mem[80056] = 16'b0000000000000000;
	sram_mem[80057] = 16'b0000000000000000;
	sram_mem[80058] = 16'b0000000000000000;
	sram_mem[80059] = 16'b0000000000000000;
	sram_mem[80060] = 16'b0000000000000000;
	sram_mem[80061] = 16'b0000000000000000;
	sram_mem[80062] = 16'b0000000000000000;
	sram_mem[80063] = 16'b0000000000000000;
	sram_mem[80064] = 16'b0000000000000000;
	sram_mem[80065] = 16'b0000000000000000;
	sram_mem[80066] = 16'b0000000000000000;
	sram_mem[80067] = 16'b0000000000000000;
	sram_mem[80068] = 16'b0000000000000000;
	sram_mem[80069] = 16'b0000000000000000;
	sram_mem[80070] = 16'b0000000000000000;
	sram_mem[80071] = 16'b0000000000000000;
	sram_mem[80072] = 16'b0000000000000000;
	sram_mem[80073] = 16'b0000000000000000;
	sram_mem[80074] = 16'b0000000000000000;
	sram_mem[80075] = 16'b0000000000000000;
	sram_mem[80076] = 16'b0000000000000000;
	sram_mem[80077] = 16'b0000000000000000;
	sram_mem[80078] = 16'b0000000000000000;
	sram_mem[80079] = 16'b0000000000000000;
	sram_mem[80080] = 16'b0000000000000000;
	sram_mem[80081] = 16'b0000000000000000;
	sram_mem[80082] = 16'b0000000000000000;
	sram_mem[80083] = 16'b0000000000000000;
	sram_mem[80084] = 16'b0000000000000000;
	sram_mem[80085] = 16'b0000000000000000;
	sram_mem[80086] = 16'b0000000000000000;
	sram_mem[80087] = 16'b0000000000000000;
	sram_mem[80088] = 16'b0000000000000000;
	sram_mem[80089] = 16'b0000000000000000;
	sram_mem[80090] = 16'b0000000000000000;
	sram_mem[80091] = 16'b0000000000000000;
	sram_mem[80092] = 16'b0000000000000000;
	sram_mem[80093] = 16'b0000000000000000;
	sram_mem[80094] = 16'b0000000000000000;
	sram_mem[80095] = 16'b0000000000000000;
	sram_mem[80096] = 16'b0000000000000000;
	sram_mem[80097] = 16'b0000000000000000;
	sram_mem[80098] = 16'b0000000000000000;
	sram_mem[80099] = 16'b0000000000000000;
	sram_mem[80100] = 16'b0000000000000000;
	sram_mem[80101] = 16'b0000000000000000;
	sram_mem[80102] = 16'b0000000000000000;
	sram_mem[80103] = 16'b0000000000000000;
	sram_mem[80104] = 16'b0000000000000000;
	sram_mem[80105] = 16'b0000000000000000;
	sram_mem[80106] = 16'b0000000000000000;
	sram_mem[80107] = 16'b0000000000000000;
	sram_mem[80108] = 16'b0000000000000000;
	sram_mem[80109] = 16'b0000000000000000;
	sram_mem[80110] = 16'b0000000000000000;
	sram_mem[80111] = 16'b0000000000000000;
	sram_mem[80112] = 16'b0000000000000000;
	sram_mem[80113] = 16'b0000000000000000;
	sram_mem[80114] = 16'b0000000000000000;
	sram_mem[80115] = 16'b0000000000000000;
	sram_mem[80116] = 16'b0000000000000000;
	sram_mem[80117] = 16'b0000000000000000;
	sram_mem[80118] = 16'b0000000000000000;
	sram_mem[80119] = 16'b0000000000000000;
	sram_mem[80120] = 16'b0000000000000000;
	sram_mem[80121] = 16'b0000000000000000;
	sram_mem[80122] = 16'b0000000000000000;
	sram_mem[80123] = 16'b0000000000000000;
	sram_mem[80124] = 16'b0000000000000000;
	sram_mem[80125] = 16'b0000000000000000;
	sram_mem[80126] = 16'b0000000000000000;
	sram_mem[80127] = 16'b0000000000000000;
	sram_mem[80128] = 16'b0000000000000000;
	sram_mem[80129] = 16'b0000000000000000;
	sram_mem[80130] = 16'b0000000000000000;
	sram_mem[80131] = 16'b0000000000000000;
	sram_mem[80132] = 16'b0000000000000000;
	sram_mem[80133] = 16'b0000000000000000;
	sram_mem[80134] = 16'b0000000000000000;
	sram_mem[80135] = 16'b0000000000000000;
	sram_mem[80136] = 16'b0000000000000000;
	sram_mem[80137] = 16'b0000000000000000;
	sram_mem[80138] = 16'b0000000000000000;
	sram_mem[80139] = 16'b0000000000000000;
	sram_mem[80140] = 16'b0000000000000000;
	sram_mem[80141] = 16'b0000000000000000;
	sram_mem[80142] = 16'b0000000000000000;
	sram_mem[80143] = 16'b0000000000000000;
	sram_mem[80144] = 16'b0000000000000000;
	sram_mem[80145] = 16'b0000000000000000;
	sram_mem[80146] = 16'b0000000000000000;
	sram_mem[80147] = 16'b0000000000000000;
	sram_mem[80148] = 16'b0000000000000000;
	sram_mem[80149] = 16'b0000000000000000;
	sram_mem[80150] = 16'b0000000000000000;
	sram_mem[80151] = 16'b0000000000000000;
	sram_mem[80152] = 16'b0000000000000000;
	sram_mem[80153] = 16'b0000000000000000;
	sram_mem[80154] = 16'b0000000000000000;
	sram_mem[80155] = 16'b0000000000000000;
	sram_mem[80156] = 16'b0000000000000000;
	sram_mem[80157] = 16'b0000000000000000;
	sram_mem[80158] = 16'b0000000000000000;
	sram_mem[80159] = 16'b0000000000000000;
	sram_mem[80160] = 16'b0000000000000000;
	sram_mem[80161] = 16'b0000000000000000;
	sram_mem[80162] = 16'b0000000000000000;
	sram_mem[80163] = 16'b0000000000000000;
	sram_mem[80164] = 16'b0000000000000000;
	sram_mem[80165] = 16'b0000000000000000;
	sram_mem[80166] = 16'b0000000000000000;
	sram_mem[80167] = 16'b0000000000000000;
	sram_mem[80168] = 16'b0000000000000000;
	sram_mem[80169] = 16'b0000000000000000;
	sram_mem[80170] = 16'b0000000000000000;
	sram_mem[80171] = 16'b0000000000000000;
	sram_mem[80172] = 16'b0000000000000000;
	sram_mem[80173] = 16'b0000000000000000;
	sram_mem[80174] = 16'b0000000000000000;
	sram_mem[80175] = 16'b0000000000000000;
	sram_mem[80176] = 16'b0000000000000000;
	sram_mem[80177] = 16'b0000000000000000;
	sram_mem[80178] = 16'b0000000000000000;
	sram_mem[80179] = 16'b0000000000000000;
	sram_mem[80180] = 16'b0000000000000000;
	sram_mem[80181] = 16'b0000000000000000;
	sram_mem[80182] = 16'b0000000000000000;
	sram_mem[80183] = 16'b0000000000000000;
	sram_mem[80184] = 16'b0000000000000000;
	sram_mem[80185] = 16'b0000000000000000;
	sram_mem[80186] = 16'b0000000000000000;
	sram_mem[80187] = 16'b0000000000000000;
	sram_mem[80188] = 16'b0000000000000000;
	sram_mem[80189] = 16'b0000000000000000;
	sram_mem[80190] = 16'b0000000000000000;
	sram_mem[80191] = 16'b0000000000000000;
	sram_mem[80192] = 16'b0000000000000000;
	sram_mem[80193] = 16'b0000000000000000;
	sram_mem[80194] = 16'b0000000000000000;
	sram_mem[80195] = 16'b0000000000000000;
	sram_mem[80196] = 16'b0000000000000000;
	sram_mem[80197] = 16'b0000000000000000;
	sram_mem[80198] = 16'b0000000000000000;
	sram_mem[80199] = 16'b0000000000000000;
	sram_mem[80200] = 16'b0000000000000000;
	sram_mem[80201] = 16'b0000000000000000;
	sram_mem[80202] = 16'b0000000000000000;
	sram_mem[80203] = 16'b0000000000000000;
	sram_mem[80204] = 16'b0000000000000000;
	sram_mem[80205] = 16'b0000000000000000;
	sram_mem[80206] = 16'b0000000000000000;
	sram_mem[80207] = 16'b0000000000000000;
	sram_mem[80208] = 16'b0000000000000000;
	sram_mem[80209] = 16'b0000000000000000;
	sram_mem[80210] = 16'b0000000000000000;
	sram_mem[80211] = 16'b0000000000000000;
	sram_mem[80212] = 16'b0000000000000000;
	sram_mem[80213] = 16'b0000000000000000;
	sram_mem[80214] = 16'b0000000000000000;
	sram_mem[80215] = 16'b0000000000000000;
	sram_mem[80216] = 16'b0000000000000000;
	sram_mem[80217] = 16'b0000000000000000;
	sram_mem[80218] = 16'b0000000000000000;
	sram_mem[80219] = 16'b0000000000000000;
	sram_mem[80220] = 16'b0000000000000000;
	sram_mem[80221] = 16'b0000000000000000;
	sram_mem[80222] = 16'b0000000000000000;
	sram_mem[80223] = 16'b0000000000000000;
	sram_mem[80224] = 16'b0000000000000000;
	sram_mem[80225] = 16'b0000000000000000;
	sram_mem[80226] = 16'b0000000000000000;
	sram_mem[80227] = 16'b0000000000000000;
	sram_mem[80228] = 16'b0000000000000000;
	sram_mem[80229] = 16'b0000000000000000;
	sram_mem[80230] = 16'b0000000000000000;
	sram_mem[80231] = 16'b0000000000000000;
	sram_mem[80232] = 16'b0000000000000000;
	sram_mem[80233] = 16'b0000000000000000;
	sram_mem[80234] = 16'b0000000000000000;
	sram_mem[80235] = 16'b0000000000000000;
	sram_mem[80236] = 16'b0000000000000000;
	sram_mem[80237] = 16'b0000000000000000;
	sram_mem[80238] = 16'b0000000000000000;
	sram_mem[80239] = 16'b0000000000000000;
	sram_mem[80240] = 16'b0000000000000000;
	sram_mem[80241] = 16'b0000000000000000;
	sram_mem[80242] = 16'b0000000000000000;
	sram_mem[80243] = 16'b0000000000000000;
	sram_mem[80244] = 16'b0000000000000000;
	sram_mem[80245] = 16'b0000000000000000;
	sram_mem[80246] = 16'b0000000000000000;
	sram_mem[80247] = 16'b0000000000000000;
	sram_mem[80248] = 16'b0000000000000000;
	sram_mem[80249] = 16'b0000000000000000;
	sram_mem[80250] = 16'b0000000000000000;
	sram_mem[80251] = 16'b0000000000000000;
	sram_mem[80252] = 16'b0000000000000000;
	sram_mem[80253] = 16'b0000000000000000;
	sram_mem[80254] = 16'b0000000000000000;
	sram_mem[80255] = 16'b0000000000000000;
	sram_mem[80256] = 16'b0000000000000000;
	sram_mem[80257] = 16'b0000000000000000;
	sram_mem[80258] = 16'b0000000000000000;
	sram_mem[80259] = 16'b0000000000000000;
	sram_mem[80260] = 16'b0000000000000000;
	sram_mem[80261] = 16'b0000000000000000;
	sram_mem[80262] = 16'b0000000000000000;
	sram_mem[80263] = 16'b0000000000000000;
	sram_mem[80264] = 16'b0000000000000000;
	sram_mem[80265] = 16'b0000000000000000;
	sram_mem[80266] = 16'b0000000000000000;
	sram_mem[80267] = 16'b0000000000000000;
	sram_mem[80268] = 16'b0000000000000000;
	sram_mem[80269] = 16'b0000000000000000;
	sram_mem[80270] = 16'b0000000000000000;
	sram_mem[80271] = 16'b0000000000000000;
	sram_mem[80272] = 16'b0000000000000000;
	sram_mem[80273] = 16'b0000000000000000;
	sram_mem[80274] = 16'b0000000000000000;
	sram_mem[80275] = 16'b0000000000000000;
	sram_mem[80276] = 16'b0000000000000000;
	sram_mem[80277] = 16'b0000000000000000;
	sram_mem[80278] = 16'b0000000000000000;
	sram_mem[80279] = 16'b0000000000000000;
	sram_mem[80280] = 16'b0000000000000000;
	sram_mem[80281] = 16'b0000000000000000;
	sram_mem[80282] = 16'b0000000000000000;
	sram_mem[80283] = 16'b0000000000000000;
	sram_mem[80284] = 16'b0000000000000000;
	sram_mem[80285] = 16'b0000000000000000;
	sram_mem[80286] = 16'b0000000000000000;
	sram_mem[80287] = 16'b0000000000000000;
	sram_mem[80288] = 16'b0000000000000000;
	sram_mem[80289] = 16'b0000000000000000;
	sram_mem[80290] = 16'b0000000000000000;
	sram_mem[80291] = 16'b0000000000000000;
	sram_mem[80292] = 16'b0000000000000000;
	sram_mem[80293] = 16'b0000000000000000;
	sram_mem[80294] = 16'b0000000000000000;
	sram_mem[80295] = 16'b0000000000000000;
	sram_mem[80296] = 16'b0000000000000000;
	sram_mem[80297] = 16'b0000000000000000;
	sram_mem[80298] = 16'b0000000000000000;
	sram_mem[80299] = 16'b0000000000000000;
	sram_mem[80300] = 16'b0000000000000000;
	sram_mem[80301] = 16'b0000000000000000;
	sram_mem[80302] = 16'b0000000000000000;
	sram_mem[80303] = 16'b0000000000000000;
	sram_mem[80304] = 16'b0000000000000000;
	sram_mem[80305] = 16'b0000000000000000;
	sram_mem[80306] = 16'b0000000000000000;
	sram_mem[80307] = 16'b0000000000000000;
	sram_mem[80308] = 16'b0000000000000000;
	sram_mem[80309] = 16'b0000000000000000;
	sram_mem[80310] = 16'b0000000000000000;
	sram_mem[80311] = 16'b0000000000000000;
	sram_mem[80312] = 16'b0000000000000000;
	sram_mem[80313] = 16'b0000000000000000;
	sram_mem[80314] = 16'b0000000000000000;
	sram_mem[80315] = 16'b0000000000000000;
	sram_mem[80316] = 16'b0000000000000000;
	sram_mem[80317] = 16'b0000000000000000;
	sram_mem[80318] = 16'b0000000000000000;
	sram_mem[80319] = 16'b0000000000000000;
	sram_mem[80320] = 16'b0000000000000000;
	sram_mem[80321] = 16'b0000000000000000;
	sram_mem[80322] = 16'b0000000000000000;
	sram_mem[80323] = 16'b0000000000000000;
	sram_mem[80324] = 16'b0000000000000000;
	sram_mem[80325] = 16'b0000000000000000;
	sram_mem[80326] = 16'b0000000000000000;
	sram_mem[80327] = 16'b0000000000000000;
	sram_mem[80328] = 16'b0000000000000000;
	sram_mem[80329] = 16'b0000000000000000;
	sram_mem[80330] = 16'b0000000000000000;
	sram_mem[80331] = 16'b0000000000000000;
	sram_mem[80332] = 16'b0000000000000000;
	sram_mem[80333] = 16'b0000000000000000;
	sram_mem[80334] = 16'b0000000000000000;
	sram_mem[80335] = 16'b0000000000000000;
	sram_mem[80336] = 16'b0000000000000000;
	sram_mem[80337] = 16'b0000000000000000;
	sram_mem[80338] = 16'b0000000000000000;
	sram_mem[80339] = 16'b0000000000000000;
	sram_mem[80340] = 16'b0000000000000000;
	sram_mem[80341] = 16'b0000000000000000;
	sram_mem[80342] = 16'b0000000000000000;
	sram_mem[80343] = 16'b0000000000000000;
	sram_mem[80344] = 16'b0000000000000000;
	sram_mem[80345] = 16'b0000000000000000;
	sram_mem[80346] = 16'b0000000000000000;
	sram_mem[80347] = 16'b0000000000000000;
	sram_mem[80348] = 16'b0000000000000000;
	sram_mem[80349] = 16'b0000000000000000;
	sram_mem[80350] = 16'b0000000000000000;
	sram_mem[80351] = 16'b0000000000000000;
	sram_mem[80352] = 16'b0000000000000000;
	sram_mem[80353] = 16'b0000000000000000;
	sram_mem[80354] = 16'b0000000000000000;
	sram_mem[80355] = 16'b0000000000000000;
	sram_mem[80356] = 16'b0000000000000000;
	sram_mem[80357] = 16'b0000000000000000;
	sram_mem[80358] = 16'b0000000000000000;
	sram_mem[80359] = 16'b0000000000000000;
	sram_mem[80360] = 16'b0000000000000000;
	sram_mem[80361] = 16'b0000000000000000;
	sram_mem[80362] = 16'b0000000000000000;
	sram_mem[80363] = 16'b0000000000000000;
	sram_mem[80364] = 16'b0000000000000000;
	sram_mem[80365] = 16'b0000000000000000;
	sram_mem[80366] = 16'b0000000000000000;
	sram_mem[80367] = 16'b0000000000000000;
	sram_mem[80368] = 16'b0000000000000000;
	sram_mem[80369] = 16'b0000000000000000;
	sram_mem[80370] = 16'b0000000000000000;
	sram_mem[80371] = 16'b0000000000000000;
	sram_mem[80372] = 16'b0000000000000000;
	sram_mem[80373] = 16'b0000000000000000;
	sram_mem[80374] = 16'b0000000000000000;
	sram_mem[80375] = 16'b0000000000000000;
	sram_mem[80376] = 16'b0000000000000000;
	sram_mem[80377] = 16'b0000000000000000;
	sram_mem[80378] = 16'b0000000000000000;
	sram_mem[80379] = 16'b0000000000000000;
	sram_mem[80380] = 16'b0000000000000000;
	sram_mem[80381] = 16'b0000000000000000;
	sram_mem[80382] = 16'b0000000000000000;
	sram_mem[80383] = 16'b0000000000000000;
	sram_mem[80384] = 16'b0000000000000000;
	sram_mem[80385] = 16'b0000000000000000;
	sram_mem[80386] = 16'b0000000000000000;
	sram_mem[80387] = 16'b0000000000000000;
	sram_mem[80388] = 16'b0000000000000000;
	sram_mem[80389] = 16'b0000000000000000;
	sram_mem[80390] = 16'b0000000000000000;
	sram_mem[80391] = 16'b0000000000000000;
	sram_mem[80392] = 16'b0000000000000000;
	sram_mem[80393] = 16'b0000000000000000;
	sram_mem[80394] = 16'b0000000000000000;
	sram_mem[80395] = 16'b0000000000000000;
	sram_mem[80396] = 16'b0000000000000000;
	sram_mem[80397] = 16'b0000000000000000;
	sram_mem[80398] = 16'b0000000000000000;
	sram_mem[80399] = 16'b0000000000000000;
	sram_mem[80400] = 16'b0000000000000000;
	sram_mem[80401] = 16'b0000000000000000;
	sram_mem[80402] = 16'b0000000000000000;
	sram_mem[80403] = 16'b0000000000000000;
	sram_mem[80404] = 16'b0000000000000000;
	sram_mem[80405] = 16'b0000000000000000;
	sram_mem[80406] = 16'b0000000000000000;
	sram_mem[80407] = 16'b0000000000000000;
	sram_mem[80408] = 16'b0000000000000000;
	sram_mem[80409] = 16'b0000000000000000;
	sram_mem[80410] = 16'b0000000000000000;
	sram_mem[80411] = 16'b0000000000000000;
	sram_mem[80412] = 16'b0000000000000000;
	sram_mem[80413] = 16'b0000000000000000;
	sram_mem[80414] = 16'b0000000000000000;
	sram_mem[80415] = 16'b0000000000000000;
	sram_mem[80416] = 16'b0000000000000000;
	sram_mem[80417] = 16'b0000000000000000;
	sram_mem[80418] = 16'b0000000000000000;
	sram_mem[80419] = 16'b0000000000000000;
	sram_mem[80420] = 16'b0000000000000000;
	sram_mem[80421] = 16'b0000000000000000;
	sram_mem[80422] = 16'b0000000000000000;
	sram_mem[80423] = 16'b0000000000000000;
	sram_mem[80424] = 16'b0000000000000000;
	sram_mem[80425] = 16'b0000000000000000;
	sram_mem[80426] = 16'b0000000000000000;
	sram_mem[80427] = 16'b0000000000000000;
	sram_mem[80428] = 16'b0000000000000000;
	sram_mem[80429] = 16'b0000000000000000;
	sram_mem[80430] = 16'b0000000000000000;
	sram_mem[80431] = 16'b0000000000000000;
	sram_mem[80432] = 16'b0000000000000000;
	sram_mem[80433] = 16'b0000000000000000;
	sram_mem[80434] = 16'b0000000000000000;
	sram_mem[80435] = 16'b0000000000000000;
	sram_mem[80436] = 16'b0000000000000000;
	sram_mem[80437] = 16'b0000000000000000;
	sram_mem[80438] = 16'b0000000000000000;
	sram_mem[80439] = 16'b0000000000000000;
	sram_mem[80440] = 16'b0000000000000000;
	sram_mem[80441] = 16'b0000000000000000;
	sram_mem[80442] = 16'b0000000000000000;
	sram_mem[80443] = 16'b0000000000000000;
	sram_mem[80444] = 16'b0000000000000000;
	sram_mem[80445] = 16'b0000000000000000;
	sram_mem[80446] = 16'b0000000000000000;
	sram_mem[80447] = 16'b0000000000000000;
	sram_mem[80448] = 16'b0000000000000000;
	sram_mem[80449] = 16'b0000000000000000;
	sram_mem[80450] = 16'b0000000000000000;
	sram_mem[80451] = 16'b0000000000000000;
	sram_mem[80452] = 16'b0000000000000000;
	sram_mem[80453] = 16'b0000000000000000;
	sram_mem[80454] = 16'b0000000000000000;
	sram_mem[80455] = 16'b0000000000000000;
	sram_mem[80456] = 16'b0000000000000000;
	sram_mem[80457] = 16'b0000000000000000;
	sram_mem[80458] = 16'b0000000000000000;
	sram_mem[80459] = 16'b0000000000000000;
	sram_mem[80460] = 16'b0000000000000000;
	sram_mem[80461] = 16'b0000000000000000;
	sram_mem[80462] = 16'b0000000000000000;
	sram_mem[80463] = 16'b0000000000000000;
	sram_mem[80464] = 16'b0000000000000000;
	sram_mem[80465] = 16'b0000000000000000;
	sram_mem[80466] = 16'b0000000000000000;
	sram_mem[80467] = 16'b0000000000000000;
	sram_mem[80468] = 16'b0000000000000000;
	sram_mem[80469] = 16'b0000000000000000;
	sram_mem[80470] = 16'b0000000000000000;
	sram_mem[80471] = 16'b0000000000000000;
	sram_mem[80472] = 16'b0000000000000000;
	sram_mem[80473] = 16'b0000000000000000;
	sram_mem[80474] = 16'b0000000000000000;
	sram_mem[80475] = 16'b0000000000000000;
	sram_mem[80476] = 16'b0000000000000000;
	sram_mem[80477] = 16'b0000000000000000;
	sram_mem[80478] = 16'b0000000000000000;
	sram_mem[80479] = 16'b0000000000000000;
	sram_mem[80480] = 16'b0000000000000000;
	sram_mem[80481] = 16'b0000000000000000;
	sram_mem[80482] = 16'b0000000000000000;
	sram_mem[80483] = 16'b0000000000000000;
	sram_mem[80484] = 16'b0000000000000000;
	sram_mem[80485] = 16'b0000000000000000;
	sram_mem[80486] = 16'b0000000000000000;
	sram_mem[80487] = 16'b0000000000000000;
	sram_mem[80488] = 16'b0000000000000000;
	sram_mem[80489] = 16'b0000000000000000;
	sram_mem[80490] = 16'b0000000000000000;
	sram_mem[80491] = 16'b0000000000000000;
	sram_mem[80492] = 16'b0000000000000000;
	sram_mem[80493] = 16'b0000000000000000;
	sram_mem[80494] = 16'b0000000000000000;
	sram_mem[80495] = 16'b0000000000000000;
	sram_mem[80496] = 16'b0000000000000000;
	sram_mem[80497] = 16'b0000000000000000;
	sram_mem[80498] = 16'b0000000000000000;
	sram_mem[80499] = 16'b0000000000000000;
	sram_mem[80500] = 16'b0000000000000000;
	sram_mem[80501] = 16'b0000000000000000;
	sram_mem[80502] = 16'b0000000000000000;
	sram_mem[80503] = 16'b0000000000000000;
	sram_mem[80504] = 16'b0000000000000000;
	sram_mem[80505] = 16'b0000000000000000;
	sram_mem[80506] = 16'b0000000000000000;
	sram_mem[80507] = 16'b0000000000000000;
	sram_mem[80508] = 16'b0000000000000000;
	sram_mem[80509] = 16'b0000000000000000;
	sram_mem[80510] = 16'b0000000000000000;
	sram_mem[80511] = 16'b0000000000000000;
	sram_mem[80512] = 16'b0000000000000000;
	sram_mem[80513] = 16'b0000000000000000;
	sram_mem[80514] = 16'b0000000000000000;
	sram_mem[80515] = 16'b0000000000000000;
	sram_mem[80516] = 16'b0000000000000000;
	sram_mem[80517] = 16'b0000000000000000;
	sram_mem[80518] = 16'b0000000000000000;
	sram_mem[80519] = 16'b0000000000000000;
	sram_mem[80520] = 16'b0000000000000000;
	sram_mem[80521] = 16'b0000000000000000;
	sram_mem[80522] = 16'b0000000000000000;
	sram_mem[80523] = 16'b0000000000000000;
	sram_mem[80524] = 16'b0000000000000000;
	sram_mem[80525] = 16'b0000000000000000;
	sram_mem[80526] = 16'b0000000000000000;
	sram_mem[80527] = 16'b0000000000000000;
	sram_mem[80528] = 16'b0000000000000000;
	sram_mem[80529] = 16'b0000000000000000;
	sram_mem[80530] = 16'b0000000000000000;
	sram_mem[80531] = 16'b0000000000000000;
	sram_mem[80532] = 16'b0000000000000000;
	sram_mem[80533] = 16'b0000000000000000;
	sram_mem[80534] = 16'b0000000000000000;
	sram_mem[80535] = 16'b0000000000000000;
	sram_mem[80536] = 16'b0000000000000000;
	sram_mem[80537] = 16'b0000000000000000;
	sram_mem[80538] = 16'b0000000000000000;
	sram_mem[80539] = 16'b0000000000000000;
	sram_mem[80540] = 16'b0000000000000000;
	sram_mem[80541] = 16'b0000000000000000;
	sram_mem[80542] = 16'b0000000000000000;
	sram_mem[80543] = 16'b0000000000000000;
	sram_mem[80544] = 16'b0000000000000000;
	sram_mem[80545] = 16'b0000000000000000;
	sram_mem[80546] = 16'b0000000000000000;
	sram_mem[80547] = 16'b0000000000000000;
	sram_mem[80548] = 16'b0000000000000000;
	sram_mem[80549] = 16'b0000000000000000;
	sram_mem[80550] = 16'b0000000000000000;
	sram_mem[80551] = 16'b0000000000000000;
	sram_mem[80552] = 16'b0000000000000000;
	sram_mem[80553] = 16'b0000000000000000;
	sram_mem[80554] = 16'b0000000000000000;
	sram_mem[80555] = 16'b0000000000000000;
	sram_mem[80556] = 16'b0000000000000000;
	sram_mem[80557] = 16'b0000000000000000;
	sram_mem[80558] = 16'b0000000000000000;
	sram_mem[80559] = 16'b0000000000000000;
	sram_mem[80560] = 16'b0000000000000000;
	sram_mem[80561] = 16'b0000000000000000;
	sram_mem[80562] = 16'b0000000000000000;
	sram_mem[80563] = 16'b0000000000000000;
	sram_mem[80564] = 16'b0000000000000000;
	sram_mem[80565] = 16'b0000000000000000;
	sram_mem[80566] = 16'b0000000000000000;
	sram_mem[80567] = 16'b0000000000000000;
	sram_mem[80568] = 16'b0000000000000000;
	sram_mem[80569] = 16'b0000000000000000;
	sram_mem[80570] = 16'b0000000000000000;
	sram_mem[80571] = 16'b0000000000000000;
	sram_mem[80572] = 16'b0000000000000000;
	sram_mem[80573] = 16'b0000000000000000;
	sram_mem[80574] = 16'b0000000000000000;
	sram_mem[80575] = 16'b0000000000000000;
	sram_mem[80576] = 16'b0000000000000000;
	sram_mem[80577] = 16'b0000000000000000;
	sram_mem[80578] = 16'b0000000000000000;
	sram_mem[80579] = 16'b0000000000000000;
	sram_mem[80580] = 16'b0000000000000000;
	sram_mem[80581] = 16'b0000000000000000;
	sram_mem[80582] = 16'b0000000000000000;
	sram_mem[80583] = 16'b0000000000000000;
	sram_mem[80584] = 16'b0000000000000000;
	sram_mem[80585] = 16'b0000000000000000;
	sram_mem[80586] = 16'b0000000000000000;
	sram_mem[80587] = 16'b0000000000000000;
	sram_mem[80588] = 16'b0000000000000000;
	sram_mem[80589] = 16'b0000000000000000;
	sram_mem[80590] = 16'b0000000000000000;
	sram_mem[80591] = 16'b0000000000000000;
	sram_mem[80592] = 16'b0000000000000000;
	sram_mem[80593] = 16'b0000000000000000;
	sram_mem[80594] = 16'b0000000000000000;
	sram_mem[80595] = 16'b0000000000000000;
	sram_mem[80596] = 16'b0000000000000000;
	sram_mem[80597] = 16'b0000000000000000;
	sram_mem[80598] = 16'b0000000000000000;
	sram_mem[80599] = 16'b0000000000000000;
	sram_mem[80600] = 16'b0000000000000000;
	sram_mem[80601] = 16'b0000000000000000;
	sram_mem[80602] = 16'b0000000000000000;
	sram_mem[80603] = 16'b0000000000000000;
	sram_mem[80604] = 16'b0000000000000000;
	sram_mem[80605] = 16'b0000000000000000;
	sram_mem[80606] = 16'b0000000000000000;
	sram_mem[80607] = 16'b0000000000000000;
	sram_mem[80608] = 16'b0000000000000000;
	sram_mem[80609] = 16'b0000000000000000;
	sram_mem[80610] = 16'b0000000000000000;
	sram_mem[80611] = 16'b0000000000000000;
	sram_mem[80612] = 16'b0000000000000000;
	sram_mem[80613] = 16'b0000000000000000;
	sram_mem[80614] = 16'b0000000000000000;
	sram_mem[80615] = 16'b0000000000000000;
	sram_mem[80616] = 16'b0000000000000000;
	sram_mem[80617] = 16'b0000000000000000;
	sram_mem[80618] = 16'b0000000000000000;
	sram_mem[80619] = 16'b0000000000000000;
	sram_mem[80620] = 16'b0000000000000000;
	sram_mem[80621] = 16'b0000000000000000;
	sram_mem[80622] = 16'b0000000000000000;
	sram_mem[80623] = 16'b0000000000000000;
	sram_mem[80624] = 16'b0000000000000000;
	sram_mem[80625] = 16'b0000000000000000;
	sram_mem[80626] = 16'b0000000000000000;
	sram_mem[80627] = 16'b0000000000000000;
	sram_mem[80628] = 16'b0000000000000000;
	sram_mem[80629] = 16'b0000000000000000;
	sram_mem[80630] = 16'b0000000000000000;
	sram_mem[80631] = 16'b0000000000000000;
	sram_mem[80632] = 16'b0000000000000000;
	sram_mem[80633] = 16'b0000000000000000;
	sram_mem[80634] = 16'b0000000000000000;
	sram_mem[80635] = 16'b0000000000000000;
	sram_mem[80636] = 16'b0000000000000000;
	sram_mem[80637] = 16'b0000000000000000;
	sram_mem[80638] = 16'b0000000000000000;
	sram_mem[80639] = 16'b0000000000000000;
	sram_mem[80640] = 16'b0000000000000000;
	sram_mem[80641] = 16'b0000000000000000;
	sram_mem[80642] = 16'b0000000000000000;
	sram_mem[80643] = 16'b0000000000000000;
	sram_mem[80644] = 16'b0000000000000000;
	sram_mem[80645] = 16'b0000000000000000;
	sram_mem[80646] = 16'b0000000000000000;
	sram_mem[80647] = 16'b0000000000000000;
	sram_mem[80648] = 16'b0000000000000000;
	sram_mem[80649] = 16'b0000000000000000;
	sram_mem[80650] = 16'b0000000000000000;
	sram_mem[80651] = 16'b0000000000000000;
	sram_mem[80652] = 16'b0000000000000000;
	sram_mem[80653] = 16'b0000000000000000;
	sram_mem[80654] = 16'b0000000000000000;
	sram_mem[80655] = 16'b0000000000000000;
	sram_mem[80656] = 16'b0000000000000000;
	sram_mem[80657] = 16'b0000000000000000;
	sram_mem[80658] = 16'b0000000000000000;
	sram_mem[80659] = 16'b0000000000000000;
	sram_mem[80660] = 16'b0000000000000000;
	sram_mem[80661] = 16'b0000000000000000;
	sram_mem[80662] = 16'b0000000000000000;
	sram_mem[80663] = 16'b0000000000000000;
	sram_mem[80664] = 16'b0000000000000000;
	sram_mem[80665] = 16'b0000000000000000;
	sram_mem[80666] = 16'b0000000000000000;
	sram_mem[80667] = 16'b0000000000000000;
	sram_mem[80668] = 16'b0000000000000000;
	sram_mem[80669] = 16'b0000000000000000;
	sram_mem[80670] = 16'b0000000000000000;
	sram_mem[80671] = 16'b0000000000000000;
	sram_mem[80672] = 16'b0000000000000000;
	sram_mem[80673] = 16'b0000000000000000;
	sram_mem[80674] = 16'b0000000000000000;
	sram_mem[80675] = 16'b0000000000000000;
	sram_mem[80676] = 16'b0000000000000000;
	sram_mem[80677] = 16'b0000000000000000;
	sram_mem[80678] = 16'b0000000000000000;
	sram_mem[80679] = 16'b0000000000000000;
	sram_mem[80680] = 16'b0000000000000000;
	sram_mem[80681] = 16'b0000000000000000;
	sram_mem[80682] = 16'b0000000000000000;
	sram_mem[80683] = 16'b0000000000000000;
	sram_mem[80684] = 16'b0000000000000000;
	sram_mem[80685] = 16'b0000000000000000;
	sram_mem[80686] = 16'b0000000000000000;
	sram_mem[80687] = 16'b0000000000000000;
	sram_mem[80688] = 16'b0000000000000000;
	sram_mem[80689] = 16'b0000000000000000;
	sram_mem[80690] = 16'b0000000000000000;
	sram_mem[80691] = 16'b0000000000000000;
	sram_mem[80692] = 16'b0000000000000000;
	sram_mem[80693] = 16'b0000000000000000;
	sram_mem[80694] = 16'b0000000000000000;
	sram_mem[80695] = 16'b0000000000000000;
	sram_mem[80696] = 16'b0000000000000000;
	sram_mem[80697] = 16'b0000000000000000;
	sram_mem[80698] = 16'b0000000000000000;
	sram_mem[80699] = 16'b0000000000000000;
	sram_mem[80700] = 16'b0000000000000000;
	sram_mem[80701] = 16'b0000000000000000;
	sram_mem[80702] = 16'b0000000000000000;
	sram_mem[80703] = 16'b0000000000000000;
	sram_mem[80704] = 16'b0000000000000000;
	sram_mem[80705] = 16'b0000000000000000;
	sram_mem[80706] = 16'b0000000000000000;
	sram_mem[80707] = 16'b0000000000000000;
	sram_mem[80708] = 16'b0000000000000000;
	sram_mem[80709] = 16'b0000000000000000;
	sram_mem[80710] = 16'b0000000000000000;
	sram_mem[80711] = 16'b0000000000000000;
	sram_mem[80712] = 16'b0000000000000000;
	sram_mem[80713] = 16'b0000000000000000;
	sram_mem[80714] = 16'b0000000000000000;
	sram_mem[80715] = 16'b0000000000000000;
	sram_mem[80716] = 16'b0000000000000000;
	sram_mem[80717] = 16'b0000000000000000;
	sram_mem[80718] = 16'b0000000000000000;
	sram_mem[80719] = 16'b0000000000000000;
	sram_mem[80720] = 16'b0000000000000000;
	sram_mem[80721] = 16'b0000000000000000;
	sram_mem[80722] = 16'b0000000000000000;
	sram_mem[80723] = 16'b0000000000000000;
	sram_mem[80724] = 16'b0000000000000000;
	sram_mem[80725] = 16'b0000000000000000;
	sram_mem[80726] = 16'b0000000000000000;
	sram_mem[80727] = 16'b0000000000000000;
	sram_mem[80728] = 16'b0000000000000000;
	sram_mem[80729] = 16'b0000000000000000;
	sram_mem[80730] = 16'b0000000000000000;
	sram_mem[80731] = 16'b0000000000000000;
	sram_mem[80732] = 16'b0000000000000000;
	sram_mem[80733] = 16'b0000000000000000;
	sram_mem[80734] = 16'b0000000000000000;
	sram_mem[80735] = 16'b0000000000000000;
	sram_mem[80736] = 16'b0000000000000000;
	sram_mem[80737] = 16'b0000000000000000;
	sram_mem[80738] = 16'b0000000000000000;
	sram_mem[80739] = 16'b0000000000000000;
	sram_mem[80740] = 16'b0000000000000000;
	sram_mem[80741] = 16'b0000000000000000;
	sram_mem[80742] = 16'b0000000000000000;
	sram_mem[80743] = 16'b0000000000000000;
	sram_mem[80744] = 16'b0000000000000000;
	sram_mem[80745] = 16'b0000000000000000;
	sram_mem[80746] = 16'b0000000000000000;
	sram_mem[80747] = 16'b0000000000000000;
	sram_mem[80748] = 16'b0000000000000000;
	sram_mem[80749] = 16'b0000000000000000;
	sram_mem[80750] = 16'b0000000000000000;
	sram_mem[80751] = 16'b0000000000000000;
	sram_mem[80752] = 16'b0000000000000000;
	sram_mem[80753] = 16'b0000000000000000;
	sram_mem[80754] = 16'b0000000000000000;
	sram_mem[80755] = 16'b0000000000000000;
	sram_mem[80756] = 16'b0000000000000000;
	sram_mem[80757] = 16'b0000000000000000;
	sram_mem[80758] = 16'b0000000000000000;
	sram_mem[80759] = 16'b0000000000000000;
	sram_mem[80760] = 16'b0000000000000000;
	sram_mem[80761] = 16'b0000000000000000;
	sram_mem[80762] = 16'b0000000000000000;
	sram_mem[80763] = 16'b0000000000000000;
	sram_mem[80764] = 16'b0000000000000000;
	sram_mem[80765] = 16'b0000000000000000;
	sram_mem[80766] = 16'b0000000000000000;
	sram_mem[80767] = 16'b0000000000000000;
	sram_mem[80768] = 16'b0000000000000000;
	sram_mem[80769] = 16'b0000000000000000;
	sram_mem[80770] = 16'b0000000000000000;
	sram_mem[80771] = 16'b0000000000000000;
	sram_mem[80772] = 16'b0000000000000000;
	sram_mem[80773] = 16'b0000000000000000;
	sram_mem[80774] = 16'b0000000000000000;
	sram_mem[80775] = 16'b0000000000000000;
	sram_mem[80776] = 16'b0000000000000000;
	sram_mem[80777] = 16'b0000000000000000;
	sram_mem[80778] = 16'b0000000000000000;
	sram_mem[80779] = 16'b0000000000000000;
	sram_mem[80780] = 16'b0000000000000000;
	sram_mem[80781] = 16'b0000000000000000;
	sram_mem[80782] = 16'b0000000000000000;
	sram_mem[80783] = 16'b0000000000000000;
	sram_mem[80784] = 16'b0000000000000000;
	sram_mem[80785] = 16'b0000000000000000;
	sram_mem[80786] = 16'b0000000000000000;
	sram_mem[80787] = 16'b0000000000000000;
	sram_mem[80788] = 16'b0000000000000000;
	sram_mem[80789] = 16'b0000000000000000;
	sram_mem[80790] = 16'b0000000000000000;
	sram_mem[80791] = 16'b0000000000000000;
	sram_mem[80792] = 16'b0000000000000000;
	sram_mem[80793] = 16'b0000000000000000;
	sram_mem[80794] = 16'b0000000000000000;
	sram_mem[80795] = 16'b0000000000000000;
	sram_mem[80796] = 16'b0000000000000000;
	sram_mem[80797] = 16'b0000000000000000;
	sram_mem[80798] = 16'b0000000000000000;
	sram_mem[80799] = 16'b0000000000000000;
	sram_mem[80800] = 16'b0000000000000000;
	sram_mem[80801] = 16'b0000000000000000;
	sram_mem[80802] = 16'b0000000000000000;
	sram_mem[80803] = 16'b0000000000000000;
	sram_mem[80804] = 16'b0000000000000000;
	sram_mem[80805] = 16'b0000000000000000;
	sram_mem[80806] = 16'b0000000000000000;
	sram_mem[80807] = 16'b0000000000000000;
	sram_mem[80808] = 16'b0000000000000000;
	sram_mem[80809] = 16'b0000000000000000;
	sram_mem[80810] = 16'b0000000000000000;
	sram_mem[80811] = 16'b0000000000000000;
	sram_mem[80812] = 16'b0000000000000000;
	sram_mem[80813] = 16'b0000000000000000;
	sram_mem[80814] = 16'b0000000000000000;
	sram_mem[80815] = 16'b0000000000000000;
	sram_mem[80816] = 16'b0000000000000000;
	sram_mem[80817] = 16'b0000000000000000;
	sram_mem[80818] = 16'b0000000000000000;
	sram_mem[80819] = 16'b0000000000000000;
	sram_mem[80820] = 16'b0000000000000000;
	sram_mem[80821] = 16'b0000000000000000;
	sram_mem[80822] = 16'b0000000000000000;
	sram_mem[80823] = 16'b0000000000000000;
	sram_mem[80824] = 16'b0000000000000000;
	sram_mem[80825] = 16'b0000000000000000;
	sram_mem[80826] = 16'b0000000000000000;
	sram_mem[80827] = 16'b0000000000000000;
	sram_mem[80828] = 16'b0000000000000000;
	sram_mem[80829] = 16'b0000000000000000;
	sram_mem[80830] = 16'b0000000000000000;
	sram_mem[80831] = 16'b0000000000000000;
	sram_mem[80832] = 16'b0000000000000000;
	sram_mem[80833] = 16'b0000000000000000;
	sram_mem[80834] = 16'b0000000000000000;
	sram_mem[80835] = 16'b0000000000000000;
	sram_mem[80836] = 16'b0000000000000000;
	sram_mem[80837] = 16'b0000000000000000;
	sram_mem[80838] = 16'b0000000000000000;
	sram_mem[80839] = 16'b0000000000000000;
	sram_mem[80840] = 16'b0000000000000000;
	sram_mem[80841] = 16'b0000000000000000;
	sram_mem[80842] = 16'b0000000000000000;
	sram_mem[80843] = 16'b0000000000000000;
	sram_mem[80844] = 16'b0000000000000000;
	sram_mem[80845] = 16'b0000000000000000;
	sram_mem[80846] = 16'b0000000000000000;
	sram_mem[80847] = 16'b0000000000000000;
	sram_mem[80848] = 16'b0000000000000000;
	sram_mem[80849] = 16'b0000000000000000;
	sram_mem[80850] = 16'b0000000000000000;
	sram_mem[80851] = 16'b0000000000000000;
	sram_mem[80852] = 16'b0000000000000000;
	sram_mem[80853] = 16'b0000000000000000;
	sram_mem[80854] = 16'b0000000000000000;
	sram_mem[80855] = 16'b0000000000000000;
	sram_mem[80856] = 16'b0000000000000000;
	sram_mem[80857] = 16'b0000000000000000;
	sram_mem[80858] = 16'b0000000000000000;
	sram_mem[80859] = 16'b0000000000000000;
	sram_mem[80860] = 16'b0000000000000000;
	sram_mem[80861] = 16'b0000000000000000;
	sram_mem[80862] = 16'b0000000000000000;
	sram_mem[80863] = 16'b0000000000000000;
	sram_mem[80864] = 16'b0000000000000000;
	sram_mem[80865] = 16'b0000000000000000;
	sram_mem[80866] = 16'b0000000000000000;
	sram_mem[80867] = 16'b0000000000000000;
	sram_mem[80868] = 16'b0000000000000000;
	sram_mem[80869] = 16'b0000000000000000;
	sram_mem[80870] = 16'b0000000000000000;
	sram_mem[80871] = 16'b0000000000000000;
	sram_mem[80872] = 16'b0000000000000000;
	sram_mem[80873] = 16'b0000000000000000;
	sram_mem[80874] = 16'b0000000000000000;
	sram_mem[80875] = 16'b0000000000000000;
	sram_mem[80876] = 16'b0000000000000000;
	sram_mem[80877] = 16'b0000000000000000;
	sram_mem[80878] = 16'b0000000000000000;
	sram_mem[80879] = 16'b0000000000000000;
	sram_mem[80880] = 16'b0000000000000000;
	sram_mem[80881] = 16'b0000000000000000;
	sram_mem[80882] = 16'b0000000000000000;
	sram_mem[80883] = 16'b0000000000000000;
	sram_mem[80884] = 16'b0000000000000000;
	sram_mem[80885] = 16'b0000000000000000;
	sram_mem[80886] = 16'b0000000000000000;
	sram_mem[80887] = 16'b0000000000000000;
	sram_mem[80888] = 16'b0000000000000000;
	sram_mem[80889] = 16'b0000000000000000;
	sram_mem[80890] = 16'b0000000000000000;
	sram_mem[80891] = 16'b0000000000000000;
	sram_mem[80892] = 16'b0000000000000000;
	sram_mem[80893] = 16'b0000000000000000;
	sram_mem[80894] = 16'b0000000000000000;
	sram_mem[80895] = 16'b0000000000000000;
	sram_mem[80896] = 16'b0000000000000000;
	sram_mem[80897] = 16'b0000000000000000;
	sram_mem[80898] = 16'b0000000000000000;
	sram_mem[80899] = 16'b0000000000000000;
	sram_mem[80900] = 16'b0000000000000000;
	sram_mem[80901] = 16'b0000000000000000;
	sram_mem[80902] = 16'b0000000000000000;
	sram_mem[80903] = 16'b0000000000000000;
	sram_mem[80904] = 16'b0000000000000000;
	sram_mem[80905] = 16'b0000000000000000;
	sram_mem[80906] = 16'b0000000000000000;
	sram_mem[80907] = 16'b0000000000000000;
	sram_mem[80908] = 16'b0000000000000000;
	sram_mem[80909] = 16'b0000000000000000;
	sram_mem[80910] = 16'b0000000000000000;
	sram_mem[80911] = 16'b0000000000000000;
	sram_mem[80912] = 16'b0000000000000000;
	sram_mem[80913] = 16'b0000000000000000;
	sram_mem[80914] = 16'b0000000000000000;
	sram_mem[80915] = 16'b0000000000000000;
	sram_mem[80916] = 16'b0000000000000000;
	sram_mem[80917] = 16'b0000000000000000;
	sram_mem[80918] = 16'b0000000000000000;
	sram_mem[80919] = 16'b0000000000000000;
	sram_mem[80920] = 16'b0000000000000000;
	sram_mem[80921] = 16'b0000000000000000;
	sram_mem[80922] = 16'b0000000000000000;
	sram_mem[80923] = 16'b0000000000000000;
	sram_mem[80924] = 16'b0000000000000000;
	sram_mem[80925] = 16'b0000000000000000;
	sram_mem[80926] = 16'b0000000000000000;
	sram_mem[80927] = 16'b0000000000000000;
	sram_mem[80928] = 16'b0000000000000000;
	sram_mem[80929] = 16'b0000000000000000;
	sram_mem[80930] = 16'b0000000000000000;
	sram_mem[80931] = 16'b0000000000000000;
	sram_mem[80932] = 16'b0000000000000000;
	sram_mem[80933] = 16'b0000000000000000;
	sram_mem[80934] = 16'b0000000000000000;
	sram_mem[80935] = 16'b0000000000000000;
	sram_mem[80936] = 16'b0000000000000000;
	sram_mem[80937] = 16'b0000000000000000;
	sram_mem[80938] = 16'b0000000000000000;
	sram_mem[80939] = 16'b0000000000000000;
	sram_mem[80940] = 16'b0000000000000000;
	sram_mem[80941] = 16'b0000000000000000;
	sram_mem[80942] = 16'b0000000000000000;
	sram_mem[80943] = 16'b0000000000000000;
	sram_mem[80944] = 16'b0000000000000000;
	sram_mem[80945] = 16'b0000000000000000;
	sram_mem[80946] = 16'b0000000000000000;
	sram_mem[80947] = 16'b0000000000000000;
	sram_mem[80948] = 16'b0000000000000000;
	sram_mem[80949] = 16'b0000000000000000;
	sram_mem[80950] = 16'b0000000000000000;
	sram_mem[80951] = 16'b0000000000000000;
	sram_mem[80952] = 16'b0000000000000000;
	sram_mem[80953] = 16'b0000000000000000;
	sram_mem[80954] = 16'b0000000000000000;
	sram_mem[80955] = 16'b0000000000000000;
	sram_mem[80956] = 16'b0000000000000000;
	sram_mem[80957] = 16'b0000000000000000;
	sram_mem[80958] = 16'b0000000000000000;
	sram_mem[80959] = 16'b0000000000000000;
	sram_mem[80960] = 16'b0000000000000000;
	sram_mem[80961] = 16'b0000000000000000;
	sram_mem[80962] = 16'b0000000000000000;
	sram_mem[80963] = 16'b0000000000000000;
	sram_mem[80964] = 16'b0000000000000000;
	sram_mem[80965] = 16'b0000000000000000;
	sram_mem[80966] = 16'b0000000000000000;
	sram_mem[80967] = 16'b0000000000000000;
	sram_mem[80968] = 16'b0000000000000000;
	sram_mem[80969] = 16'b0000000000000000;
	sram_mem[80970] = 16'b0000000000000000;
	sram_mem[80971] = 16'b0000000000000000;
	sram_mem[80972] = 16'b0000000000000000;
	sram_mem[80973] = 16'b0000000000000000;
	sram_mem[80974] = 16'b0000000000000000;
	sram_mem[80975] = 16'b0000000000000000;
	sram_mem[80976] = 16'b0000000000000000;
	sram_mem[80977] = 16'b0000000000000000;
	sram_mem[80978] = 16'b0000000000000000;
	sram_mem[80979] = 16'b0000000000000000;
	sram_mem[80980] = 16'b0000000000000000;
	sram_mem[80981] = 16'b0000000000000000;
	sram_mem[80982] = 16'b0000000000000000;
	sram_mem[80983] = 16'b0000000000000000;
	sram_mem[80984] = 16'b0000000000000000;
	sram_mem[80985] = 16'b0000000000000000;
	sram_mem[80986] = 16'b0000000000000000;
	sram_mem[80987] = 16'b0000000000000000;
	sram_mem[80988] = 16'b0000000000000000;
	sram_mem[80989] = 16'b0000000000000000;
	sram_mem[80990] = 16'b0000000000000000;
	sram_mem[80991] = 16'b0000000000000000;
	sram_mem[80992] = 16'b0000000000000000;
	sram_mem[80993] = 16'b0000000000000000;
	sram_mem[80994] = 16'b0000000000000000;
	sram_mem[80995] = 16'b0000000000000000;
	sram_mem[80996] = 16'b0000000000000000;
	sram_mem[80997] = 16'b0000000000000000;
	sram_mem[80998] = 16'b0000000000000000;
	sram_mem[80999] = 16'b0000000000000000;
	sram_mem[81000] = 16'b0000000000000000;
	sram_mem[81001] = 16'b0000000000000000;
	sram_mem[81002] = 16'b0000000000000000;
	sram_mem[81003] = 16'b0000000000000000;
	sram_mem[81004] = 16'b0000000000000000;
	sram_mem[81005] = 16'b0000000000000000;
	sram_mem[81006] = 16'b0000000000000000;
	sram_mem[81007] = 16'b0000000000000000;
	sram_mem[81008] = 16'b0000000000000000;
	sram_mem[81009] = 16'b0000000000000000;
	sram_mem[81010] = 16'b0000000000000000;
	sram_mem[81011] = 16'b0000000000000000;
	sram_mem[81012] = 16'b0000000000000000;
	sram_mem[81013] = 16'b0000000000000000;
	sram_mem[81014] = 16'b0000000000000000;
	sram_mem[81015] = 16'b0000000000000000;
	sram_mem[81016] = 16'b0000000000000000;
	sram_mem[81017] = 16'b0000000000000000;
	sram_mem[81018] = 16'b0000000000000000;
	sram_mem[81019] = 16'b0000000000000000;
	sram_mem[81020] = 16'b0000000000000000;
	sram_mem[81021] = 16'b0000000000000000;
	sram_mem[81022] = 16'b0000000000000000;
	sram_mem[81023] = 16'b0000000000000000;
	sram_mem[81024] = 16'b0000000000000000;
	sram_mem[81025] = 16'b0000000000000000;
	sram_mem[81026] = 16'b0000000000000000;
	sram_mem[81027] = 16'b0000000000000000;
	sram_mem[81028] = 16'b0000000000000000;
	sram_mem[81029] = 16'b0000000000000000;
	sram_mem[81030] = 16'b0000000000000000;
	sram_mem[81031] = 16'b0000000000000000;
	sram_mem[81032] = 16'b0000000000000000;
	sram_mem[81033] = 16'b0000000000000000;
	sram_mem[81034] = 16'b0000000000000000;
	sram_mem[81035] = 16'b0000000000000000;
	sram_mem[81036] = 16'b0000000000000000;
	sram_mem[81037] = 16'b0000000000000000;
	sram_mem[81038] = 16'b0000000000000000;
	sram_mem[81039] = 16'b0000000000000000;
	sram_mem[81040] = 16'b0000000000000000;
	sram_mem[81041] = 16'b0000000000000000;
	sram_mem[81042] = 16'b0000000000000000;
	sram_mem[81043] = 16'b0000000000000000;
	sram_mem[81044] = 16'b0000000000000000;
	sram_mem[81045] = 16'b0000000000000000;
	sram_mem[81046] = 16'b0000000000000000;
	sram_mem[81047] = 16'b0000000000000000;
	sram_mem[81048] = 16'b0000000000000000;
	sram_mem[81049] = 16'b0000000000000000;
	sram_mem[81050] = 16'b0000000000000000;
	sram_mem[81051] = 16'b0000000000000000;
	sram_mem[81052] = 16'b0000000000000000;
	sram_mem[81053] = 16'b0000000000000000;
	sram_mem[81054] = 16'b0000000000000000;
	sram_mem[81055] = 16'b0000000000000000;
	sram_mem[81056] = 16'b0000000000000000;
	sram_mem[81057] = 16'b0000000000000000;
	sram_mem[81058] = 16'b0000000000000000;
	sram_mem[81059] = 16'b0000000000000000;
	sram_mem[81060] = 16'b0000000000000000;
	sram_mem[81061] = 16'b0000000000000000;
	sram_mem[81062] = 16'b0000000000000000;
	sram_mem[81063] = 16'b0000000000000000;
	sram_mem[81064] = 16'b0000000000000000;
	sram_mem[81065] = 16'b0000000000000000;
	sram_mem[81066] = 16'b0000000000000000;
	sram_mem[81067] = 16'b0000000000000000;
	sram_mem[81068] = 16'b0000000000000000;
	sram_mem[81069] = 16'b0000000000000000;
	sram_mem[81070] = 16'b0000000000000000;
	sram_mem[81071] = 16'b0000000000000000;
	sram_mem[81072] = 16'b0000000000000000;
	sram_mem[81073] = 16'b0000000000000000;
	sram_mem[81074] = 16'b0000000000000000;
	sram_mem[81075] = 16'b0000000000000000;
	sram_mem[81076] = 16'b0000000000000000;
	sram_mem[81077] = 16'b0000000000000000;
	sram_mem[81078] = 16'b0000000000000000;
	sram_mem[81079] = 16'b0000000000000000;
	sram_mem[81080] = 16'b0000000000000000;
	sram_mem[81081] = 16'b0000000000000000;
	sram_mem[81082] = 16'b0000000000000000;
	sram_mem[81083] = 16'b0000000000000000;
	sram_mem[81084] = 16'b0000000000000000;
	sram_mem[81085] = 16'b0000000000000000;
	sram_mem[81086] = 16'b0000000000000000;
	sram_mem[81087] = 16'b0000000000000000;
	sram_mem[81088] = 16'b0000000000000000;
	sram_mem[81089] = 16'b0000000000000000;
	sram_mem[81090] = 16'b0000000000000000;
	sram_mem[81091] = 16'b0000000000000000;
	sram_mem[81092] = 16'b0000000000000000;
	sram_mem[81093] = 16'b0000000000000000;
	sram_mem[81094] = 16'b0000000000000000;
	sram_mem[81095] = 16'b0000000000000000;
	sram_mem[81096] = 16'b0000000000000000;
	sram_mem[81097] = 16'b0000000000000000;
	sram_mem[81098] = 16'b0000000000000000;
	sram_mem[81099] = 16'b0000000000000000;
	sram_mem[81100] = 16'b0000000000000000;
	sram_mem[81101] = 16'b0000000000000000;
	sram_mem[81102] = 16'b0000000000000000;
	sram_mem[81103] = 16'b0000000000000000;
	sram_mem[81104] = 16'b0000000000000000;
	sram_mem[81105] = 16'b0000000000000000;
	sram_mem[81106] = 16'b0000000000000000;
	sram_mem[81107] = 16'b0000000000000000;
	sram_mem[81108] = 16'b0000000000000000;
	sram_mem[81109] = 16'b0000000000000000;
	sram_mem[81110] = 16'b0000000000000000;
	sram_mem[81111] = 16'b0000000000000000;
	sram_mem[81112] = 16'b0000000000000000;
	sram_mem[81113] = 16'b0000000000000000;
	sram_mem[81114] = 16'b0000000000000000;
	sram_mem[81115] = 16'b0000000000000000;
	sram_mem[81116] = 16'b0000000000000000;
	sram_mem[81117] = 16'b0000000000000000;
	sram_mem[81118] = 16'b0000000000000000;
	sram_mem[81119] = 16'b0000000000000000;
	sram_mem[81120] = 16'b0000000000000000;
	sram_mem[81121] = 16'b0000000000000000;
	sram_mem[81122] = 16'b0000000000000000;
	sram_mem[81123] = 16'b0000000000000000;
	sram_mem[81124] = 16'b0000000000000000;
	sram_mem[81125] = 16'b0000000000000000;
	sram_mem[81126] = 16'b0000000000000000;
	sram_mem[81127] = 16'b0000000000000000;
	sram_mem[81128] = 16'b0000000000000000;
	sram_mem[81129] = 16'b0000000000000000;
	sram_mem[81130] = 16'b0000000000000000;
	sram_mem[81131] = 16'b0000000000000000;
	sram_mem[81132] = 16'b0000000000000000;
	sram_mem[81133] = 16'b0000000000000000;
	sram_mem[81134] = 16'b0000000000000000;
	sram_mem[81135] = 16'b0000000000000000;
	sram_mem[81136] = 16'b0000000000000000;
	sram_mem[81137] = 16'b0000000000000000;
	sram_mem[81138] = 16'b0000000000000000;
	sram_mem[81139] = 16'b0000000000000000;
	sram_mem[81140] = 16'b0000000000000000;
	sram_mem[81141] = 16'b0000000000000000;
	sram_mem[81142] = 16'b0000000000000000;
	sram_mem[81143] = 16'b0000000000000000;
	sram_mem[81144] = 16'b0000000000000000;
	sram_mem[81145] = 16'b0000000000000000;
	sram_mem[81146] = 16'b0000000000000000;
	sram_mem[81147] = 16'b0000000000000000;
	sram_mem[81148] = 16'b0000000000000000;
	sram_mem[81149] = 16'b0000000000000000;
	sram_mem[81150] = 16'b0000000000000000;
	sram_mem[81151] = 16'b0000000000000000;
	sram_mem[81152] = 16'b0000000000000000;
	sram_mem[81153] = 16'b0000000000000000;
	sram_mem[81154] = 16'b0000000000000000;
	sram_mem[81155] = 16'b0000000000000000;
	sram_mem[81156] = 16'b0000000000000000;
	sram_mem[81157] = 16'b0000000000000000;
	sram_mem[81158] = 16'b0000000000000000;
	sram_mem[81159] = 16'b0000000000000000;
	sram_mem[81160] = 16'b0000000000000000;
	sram_mem[81161] = 16'b0000000000000000;
	sram_mem[81162] = 16'b0000000000000000;
	sram_mem[81163] = 16'b0000000000000000;
	sram_mem[81164] = 16'b0000000000000000;
	sram_mem[81165] = 16'b0000000000000000;
	sram_mem[81166] = 16'b0000000000000000;
	sram_mem[81167] = 16'b0000000000000000;
	sram_mem[81168] = 16'b0000000000000000;
	sram_mem[81169] = 16'b0000000000000000;
	sram_mem[81170] = 16'b0000000000000000;
	sram_mem[81171] = 16'b0000000000000000;
	sram_mem[81172] = 16'b0000000000000000;
	sram_mem[81173] = 16'b0000000000000000;
	sram_mem[81174] = 16'b0000000000000000;
	sram_mem[81175] = 16'b0000000000000000;
	sram_mem[81176] = 16'b0000000000000000;
	sram_mem[81177] = 16'b0000000000000000;
	sram_mem[81178] = 16'b0000000000000000;
	sram_mem[81179] = 16'b0000000000000000;
	sram_mem[81180] = 16'b0000000000000000;
	sram_mem[81181] = 16'b0000000000000000;
	sram_mem[81182] = 16'b0000000000000000;
	sram_mem[81183] = 16'b0000000000000000;
	sram_mem[81184] = 16'b0000000000000000;
	sram_mem[81185] = 16'b0000000000000000;
	sram_mem[81186] = 16'b0000000000000000;
	sram_mem[81187] = 16'b0000000000000000;
	sram_mem[81188] = 16'b0000000000000000;
	sram_mem[81189] = 16'b0000000000000000;
	sram_mem[81190] = 16'b0000000000000000;
	sram_mem[81191] = 16'b0000000000000000;
	sram_mem[81192] = 16'b0000000000000000;
	sram_mem[81193] = 16'b0000000000000000;
	sram_mem[81194] = 16'b0000000000000000;
	sram_mem[81195] = 16'b0000000000000000;
	sram_mem[81196] = 16'b0000000000000000;
	sram_mem[81197] = 16'b0000000000000000;
	sram_mem[81198] = 16'b0000000000000000;
	sram_mem[81199] = 16'b0000000000000000;
	sram_mem[81200] = 16'b0000000000000000;
	sram_mem[81201] = 16'b0000000000000000;
	sram_mem[81202] = 16'b0000000000000000;
	sram_mem[81203] = 16'b0000000000000000;
	sram_mem[81204] = 16'b0000000000000000;
	sram_mem[81205] = 16'b0000000000000000;
	sram_mem[81206] = 16'b0000000000000000;
	sram_mem[81207] = 16'b0000000000000000;
	sram_mem[81208] = 16'b0000000000000000;
	sram_mem[81209] = 16'b0000000000000000;
	sram_mem[81210] = 16'b0000000000000000;
	sram_mem[81211] = 16'b0000000000000000;
	sram_mem[81212] = 16'b0000000000000000;
	sram_mem[81213] = 16'b0000000000000000;
	sram_mem[81214] = 16'b0000000000000000;
	sram_mem[81215] = 16'b0000000000000000;
	sram_mem[81216] = 16'b0000000000000000;
	sram_mem[81217] = 16'b0000000000000000;
	sram_mem[81218] = 16'b0000000000000000;
	sram_mem[81219] = 16'b0000000000000000;
	sram_mem[81220] = 16'b0000000000000000;
	sram_mem[81221] = 16'b0000000000000000;
	sram_mem[81222] = 16'b0000000000000000;
	sram_mem[81223] = 16'b0000000000000000;
	sram_mem[81224] = 16'b0000000000000000;
	sram_mem[81225] = 16'b0000000000000000;
	sram_mem[81226] = 16'b0000000000000000;
	sram_mem[81227] = 16'b0000000000000000;
	sram_mem[81228] = 16'b0000000000000000;
	sram_mem[81229] = 16'b0000000000000000;
	sram_mem[81230] = 16'b0000000000000000;
	sram_mem[81231] = 16'b0000000000000000;
	sram_mem[81232] = 16'b0000000000000000;
	sram_mem[81233] = 16'b0000000000000000;
	sram_mem[81234] = 16'b0000000000000000;
	sram_mem[81235] = 16'b0000000000000000;
	sram_mem[81236] = 16'b0000000000000000;
	sram_mem[81237] = 16'b0000000000000000;
	sram_mem[81238] = 16'b0000000000000000;
	sram_mem[81239] = 16'b0000000000000000;
	sram_mem[81240] = 16'b0000000000000000;
	sram_mem[81241] = 16'b0000000000000000;
	sram_mem[81242] = 16'b0000000000000000;
	sram_mem[81243] = 16'b0000000000000000;
	sram_mem[81244] = 16'b0000000000000000;
	sram_mem[81245] = 16'b0000000000000000;
	sram_mem[81246] = 16'b0000000000000000;
	sram_mem[81247] = 16'b0000000000000000;
	sram_mem[81248] = 16'b0000000000000000;
	sram_mem[81249] = 16'b0000000000000000;
	sram_mem[81250] = 16'b0000000000000000;
	sram_mem[81251] = 16'b0000000000000000;
	sram_mem[81252] = 16'b0000000000000000;
	sram_mem[81253] = 16'b0000000000000000;
	sram_mem[81254] = 16'b0000000000000000;
	sram_mem[81255] = 16'b0000000000000000;
	sram_mem[81256] = 16'b0000000000000000;
	sram_mem[81257] = 16'b0000000000000000;
	sram_mem[81258] = 16'b0000000000000000;
	sram_mem[81259] = 16'b0000000000000000;
	sram_mem[81260] = 16'b0000000000000000;
	sram_mem[81261] = 16'b0000000000000000;
	sram_mem[81262] = 16'b0000000000000000;
	sram_mem[81263] = 16'b0000000000000000;
	sram_mem[81264] = 16'b0000000000000000;
	sram_mem[81265] = 16'b0000000000000000;
	sram_mem[81266] = 16'b0000000000000000;
	sram_mem[81267] = 16'b0000000000000000;
	sram_mem[81268] = 16'b0000000000000000;
	sram_mem[81269] = 16'b0000000000000000;
	sram_mem[81270] = 16'b0000000000000000;
	sram_mem[81271] = 16'b0000000000000000;
	sram_mem[81272] = 16'b0000000000000000;
	sram_mem[81273] = 16'b0000000000000000;
	sram_mem[81274] = 16'b0000000000000000;
	sram_mem[81275] = 16'b0000000000000000;
	sram_mem[81276] = 16'b0000000000000000;
	sram_mem[81277] = 16'b0000000000000000;
	sram_mem[81278] = 16'b0000000000000000;
	sram_mem[81279] = 16'b0000000000000000;
	sram_mem[81280] = 16'b0000000000000000;
	sram_mem[81281] = 16'b0000000000000000;
	sram_mem[81282] = 16'b0000000000000000;
	sram_mem[81283] = 16'b0000000000000000;
	sram_mem[81284] = 16'b0000000000000000;
	sram_mem[81285] = 16'b0000000000000000;
	sram_mem[81286] = 16'b0000000000000000;
	sram_mem[81287] = 16'b0000000000000000;
	sram_mem[81288] = 16'b0000000000000000;
	sram_mem[81289] = 16'b0000000000000000;
	sram_mem[81290] = 16'b0000000000000000;
	sram_mem[81291] = 16'b0000000000000000;
	sram_mem[81292] = 16'b0000000000000000;
	sram_mem[81293] = 16'b0000000000000000;
	sram_mem[81294] = 16'b0000000000000000;
	sram_mem[81295] = 16'b0000000000000000;
	sram_mem[81296] = 16'b0000000000000000;
	sram_mem[81297] = 16'b0000000000000000;
	sram_mem[81298] = 16'b0000000000000000;
	sram_mem[81299] = 16'b0000000000000000;
	sram_mem[81300] = 16'b0000000000000000;
	sram_mem[81301] = 16'b0000000000000000;
	sram_mem[81302] = 16'b0000000000000000;
	sram_mem[81303] = 16'b0000000000000000;
	sram_mem[81304] = 16'b0000000000000000;
	sram_mem[81305] = 16'b0000000000000000;
	sram_mem[81306] = 16'b0000000000000000;
	sram_mem[81307] = 16'b0000000000000000;
	sram_mem[81308] = 16'b0000000000000000;
	sram_mem[81309] = 16'b0000000000000000;
	sram_mem[81310] = 16'b0000000000000000;
	sram_mem[81311] = 16'b0000000000000000;
	sram_mem[81312] = 16'b0000000000000000;
	sram_mem[81313] = 16'b0000000000000000;
	sram_mem[81314] = 16'b0000000000000000;
	sram_mem[81315] = 16'b0000000000000000;
	sram_mem[81316] = 16'b0000000000000000;
	sram_mem[81317] = 16'b0000000000000000;
	sram_mem[81318] = 16'b0000000000000000;
	sram_mem[81319] = 16'b0000000000000000;
	sram_mem[81320] = 16'b0000000000000000;
	sram_mem[81321] = 16'b0000000000000000;
	sram_mem[81322] = 16'b0000000000000000;
	sram_mem[81323] = 16'b0000000000000000;
	sram_mem[81324] = 16'b0000000000000000;
	sram_mem[81325] = 16'b0000000000000000;
	sram_mem[81326] = 16'b0000000000000000;
	sram_mem[81327] = 16'b0000000000000000;
	sram_mem[81328] = 16'b0000000000000000;
	sram_mem[81329] = 16'b0000000000000000;
	sram_mem[81330] = 16'b0000000000000000;
	sram_mem[81331] = 16'b0000000000000000;
	sram_mem[81332] = 16'b0000000000000000;
	sram_mem[81333] = 16'b0000000000000000;
	sram_mem[81334] = 16'b0000000000000000;
	sram_mem[81335] = 16'b0000000000000000;
	sram_mem[81336] = 16'b0000000000000000;
	sram_mem[81337] = 16'b0000000000000000;
	sram_mem[81338] = 16'b0000000000000000;
	sram_mem[81339] = 16'b0000000000000000;
	sram_mem[81340] = 16'b0000000000000000;
	sram_mem[81341] = 16'b0000000000000000;
	sram_mem[81342] = 16'b0000000000000000;
	sram_mem[81343] = 16'b0000000000000000;
	sram_mem[81344] = 16'b0000000000000000;
	sram_mem[81345] = 16'b0000000000000000;
	sram_mem[81346] = 16'b0000000000000000;
	sram_mem[81347] = 16'b0000000000000000;
	sram_mem[81348] = 16'b0000000000000000;
	sram_mem[81349] = 16'b0000000000000000;
	sram_mem[81350] = 16'b0000000000000000;
	sram_mem[81351] = 16'b0000000000000000;
	sram_mem[81352] = 16'b0000000000000000;
	sram_mem[81353] = 16'b0000000000000000;
	sram_mem[81354] = 16'b0000000000000000;
	sram_mem[81355] = 16'b0000000000000000;
	sram_mem[81356] = 16'b0000000000000000;
	sram_mem[81357] = 16'b0000000000000000;
	sram_mem[81358] = 16'b0000000000000000;
	sram_mem[81359] = 16'b0000000000000000;
	sram_mem[81360] = 16'b0000000000000000;
	sram_mem[81361] = 16'b0000000000000000;
	sram_mem[81362] = 16'b0000000000000000;
	sram_mem[81363] = 16'b0000000000000000;
	sram_mem[81364] = 16'b0000000000000000;
	sram_mem[81365] = 16'b0000000000000000;
	sram_mem[81366] = 16'b0000000000000000;
	sram_mem[81367] = 16'b0000000000000000;
	sram_mem[81368] = 16'b0000000000000000;
	sram_mem[81369] = 16'b0000000000000000;
	sram_mem[81370] = 16'b0000000000000000;
	sram_mem[81371] = 16'b0000000000000000;
	sram_mem[81372] = 16'b0000000000000000;
	sram_mem[81373] = 16'b0000000000000000;
	sram_mem[81374] = 16'b0000000000000000;
	sram_mem[81375] = 16'b0000000000000000;
	sram_mem[81376] = 16'b0000000000000000;
	sram_mem[81377] = 16'b0000000000000000;
	sram_mem[81378] = 16'b0000000000000000;
	sram_mem[81379] = 16'b0000000000000000;
	sram_mem[81380] = 16'b0000000000000000;
	sram_mem[81381] = 16'b0000000000000000;
	sram_mem[81382] = 16'b0000000000000000;
	sram_mem[81383] = 16'b0000000000000000;
	sram_mem[81384] = 16'b0000000000000000;
	sram_mem[81385] = 16'b0000000000000000;
	sram_mem[81386] = 16'b0000000000000000;
	sram_mem[81387] = 16'b0000000000000000;
	sram_mem[81388] = 16'b0000000000000000;
	sram_mem[81389] = 16'b0000000000000000;
	sram_mem[81390] = 16'b0000000000000000;
	sram_mem[81391] = 16'b0000000000000000;
	sram_mem[81392] = 16'b0000000000000000;
	sram_mem[81393] = 16'b0000000000000000;
	sram_mem[81394] = 16'b0000000000000000;
	sram_mem[81395] = 16'b0000000000000000;
	sram_mem[81396] = 16'b0000000000000000;
	sram_mem[81397] = 16'b0000000000000000;
	sram_mem[81398] = 16'b0000000000000000;
	sram_mem[81399] = 16'b0000000000000000;
	sram_mem[81400] = 16'b0000000000000000;
	sram_mem[81401] = 16'b0000000000000000;
	sram_mem[81402] = 16'b0000000000000000;
	sram_mem[81403] = 16'b0000000000000000;
	sram_mem[81404] = 16'b0000000000000000;
	sram_mem[81405] = 16'b0000000000000000;
	sram_mem[81406] = 16'b0000000000000000;
	sram_mem[81407] = 16'b0000000000000000;
	sram_mem[81408] = 16'b0000000000000000;
	sram_mem[81409] = 16'b0000000000000000;
	sram_mem[81410] = 16'b0000000000000000;
	sram_mem[81411] = 16'b0000000000000000;
	sram_mem[81412] = 16'b0000000000000000;
	sram_mem[81413] = 16'b0000000000000000;
	sram_mem[81414] = 16'b0000000000000000;
	sram_mem[81415] = 16'b0000000000000000;
	sram_mem[81416] = 16'b0000000000000000;
	sram_mem[81417] = 16'b0000000000000000;
	sram_mem[81418] = 16'b0000000000000000;
	sram_mem[81419] = 16'b0000000000000000;
	sram_mem[81420] = 16'b0000000000000000;
	sram_mem[81421] = 16'b0000000000000000;
	sram_mem[81422] = 16'b0000000000000000;
	sram_mem[81423] = 16'b0000000000000000;
	sram_mem[81424] = 16'b0000000000000000;
	sram_mem[81425] = 16'b0000000000000000;
	sram_mem[81426] = 16'b0000000000000000;
	sram_mem[81427] = 16'b0000000000000000;
	sram_mem[81428] = 16'b0000000000000000;
	sram_mem[81429] = 16'b0000000000000000;
	sram_mem[81430] = 16'b0000000000000000;
	sram_mem[81431] = 16'b0000000000000000;
	sram_mem[81432] = 16'b0000000000000000;
	sram_mem[81433] = 16'b0000000000000000;
	sram_mem[81434] = 16'b0000000000000000;
	sram_mem[81435] = 16'b0000000000000000;
	sram_mem[81436] = 16'b0000000000000000;
	sram_mem[81437] = 16'b0000000000000000;
	sram_mem[81438] = 16'b0000000000000000;
	sram_mem[81439] = 16'b0000000000000000;
	sram_mem[81440] = 16'b0000000000000000;
	sram_mem[81441] = 16'b0000000000000000;
	sram_mem[81442] = 16'b0000000000000000;
	sram_mem[81443] = 16'b0000000000000000;
	sram_mem[81444] = 16'b0000000000000000;
	sram_mem[81445] = 16'b0000000000000000;
	sram_mem[81446] = 16'b0000000000000000;
	sram_mem[81447] = 16'b0000000000000000;
	sram_mem[81448] = 16'b0000000000000000;
	sram_mem[81449] = 16'b0000000000000000;
	sram_mem[81450] = 16'b0000000000000000;
	sram_mem[81451] = 16'b0000000000000000;
	sram_mem[81452] = 16'b0000000000000000;
	sram_mem[81453] = 16'b0000000000000000;
	sram_mem[81454] = 16'b0000000000000000;
	sram_mem[81455] = 16'b0000000000000000;
	sram_mem[81456] = 16'b0000000000000000;
	sram_mem[81457] = 16'b0000000000000000;
	sram_mem[81458] = 16'b0000000000000000;
	sram_mem[81459] = 16'b0000000000000000;
	sram_mem[81460] = 16'b0000000000000000;
	sram_mem[81461] = 16'b0000000000000000;
	sram_mem[81462] = 16'b0000000000000000;
	sram_mem[81463] = 16'b0000000000000000;
	sram_mem[81464] = 16'b0000000000000000;
	sram_mem[81465] = 16'b0000000000000000;
	sram_mem[81466] = 16'b0000000000000000;
	sram_mem[81467] = 16'b0000000000000000;
	sram_mem[81468] = 16'b0000000000000000;
	sram_mem[81469] = 16'b0000000000000000;
	sram_mem[81470] = 16'b0000000000000000;
	sram_mem[81471] = 16'b0000000000000000;
	sram_mem[81472] = 16'b0000000000000000;
	sram_mem[81473] = 16'b0000000000000000;
	sram_mem[81474] = 16'b0000000000000000;
	sram_mem[81475] = 16'b0000000000000000;
	sram_mem[81476] = 16'b0000000000000000;
	sram_mem[81477] = 16'b0000000000000000;
	sram_mem[81478] = 16'b0000000000000000;
	sram_mem[81479] = 16'b0000000000000000;
	sram_mem[81480] = 16'b0000000000000000;
	sram_mem[81481] = 16'b0000000000000000;
	sram_mem[81482] = 16'b0000000000000000;
	sram_mem[81483] = 16'b0000000000000000;
	sram_mem[81484] = 16'b0000000000000000;
	sram_mem[81485] = 16'b0000000000000000;
	sram_mem[81486] = 16'b0000000000000000;
	sram_mem[81487] = 16'b0000000000000000;
	sram_mem[81488] = 16'b0000000000000000;
	sram_mem[81489] = 16'b0000000000000000;
	sram_mem[81490] = 16'b0000000000000000;
	sram_mem[81491] = 16'b0000000000000000;
	sram_mem[81492] = 16'b0000000000000000;
	sram_mem[81493] = 16'b0000000000000000;
	sram_mem[81494] = 16'b0000000000000000;
	sram_mem[81495] = 16'b0000000000000000;
	sram_mem[81496] = 16'b0000000000000000;
	sram_mem[81497] = 16'b0000000000000000;
	sram_mem[81498] = 16'b0000000000000000;
	sram_mem[81499] = 16'b0000000000000000;
	sram_mem[81500] = 16'b0000000000000000;
	sram_mem[81501] = 16'b0000000000000000;
	sram_mem[81502] = 16'b0000000000000000;
	sram_mem[81503] = 16'b0000000000000000;
	sram_mem[81504] = 16'b0000000000000000;
	sram_mem[81505] = 16'b0000000000000000;
	sram_mem[81506] = 16'b0000000000000000;
	sram_mem[81507] = 16'b0000000000000000;
	sram_mem[81508] = 16'b0000000000000000;
	sram_mem[81509] = 16'b0000000000000000;
	sram_mem[81510] = 16'b0000000000000000;
	sram_mem[81511] = 16'b0000000000000000;
	sram_mem[81512] = 16'b0000000000000000;
	sram_mem[81513] = 16'b0000000000000000;
	sram_mem[81514] = 16'b0000000000000000;
	sram_mem[81515] = 16'b0000000000000000;
	sram_mem[81516] = 16'b0000000000000000;
	sram_mem[81517] = 16'b0000000000000000;
	sram_mem[81518] = 16'b0000000000000000;
	sram_mem[81519] = 16'b0000000000000000;
	sram_mem[81520] = 16'b0000000000000000;
	sram_mem[81521] = 16'b0000000000000000;
	sram_mem[81522] = 16'b0000000000000000;
	sram_mem[81523] = 16'b0000000000000000;
	sram_mem[81524] = 16'b0000000000000000;
	sram_mem[81525] = 16'b0000000000000000;
	sram_mem[81526] = 16'b0000000000000000;
	sram_mem[81527] = 16'b0000000000000000;
	sram_mem[81528] = 16'b0000000000000000;
	sram_mem[81529] = 16'b0000000000000000;
	sram_mem[81530] = 16'b0000000000000000;
	sram_mem[81531] = 16'b0000000000000000;
	sram_mem[81532] = 16'b0000000000000000;
	sram_mem[81533] = 16'b0000000000000000;
	sram_mem[81534] = 16'b0000000000000000;
	sram_mem[81535] = 16'b0000000000000000;
	sram_mem[81536] = 16'b0000000000000000;
	sram_mem[81537] = 16'b0000000000000000;
	sram_mem[81538] = 16'b0000000000000000;
	sram_mem[81539] = 16'b0000000000000000;
	sram_mem[81540] = 16'b0000000000000000;
	sram_mem[81541] = 16'b0000000000000000;
	sram_mem[81542] = 16'b0000000000000000;
	sram_mem[81543] = 16'b0000000000000000;
	sram_mem[81544] = 16'b0000000000000000;
	sram_mem[81545] = 16'b0000000000000000;
	sram_mem[81546] = 16'b0000000000000000;
	sram_mem[81547] = 16'b0000000000000000;
	sram_mem[81548] = 16'b0000000000000000;
	sram_mem[81549] = 16'b0000000000000000;
	sram_mem[81550] = 16'b0000000000000000;
	sram_mem[81551] = 16'b0000000000000000;
	sram_mem[81552] = 16'b0000000000000000;
	sram_mem[81553] = 16'b0000000000000000;
	sram_mem[81554] = 16'b0000000000000000;
	sram_mem[81555] = 16'b0000000000000000;
	sram_mem[81556] = 16'b0000000000000000;
	sram_mem[81557] = 16'b0000000000000000;
	sram_mem[81558] = 16'b0000000000000000;
	sram_mem[81559] = 16'b0000000000000000;
	sram_mem[81560] = 16'b0000000000000000;
	sram_mem[81561] = 16'b0000000000000000;
	sram_mem[81562] = 16'b0000000000000000;
	sram_mem[81563] = 16'b0000000000000000;
	sram_mem[81564] = 16'b0000000000000000;
	sram_mem[81565] = 16'b0000000000000000;
	sram_mem[81566] = 16'b0000000000000000;
	sram_mem[81567] = 16'b0000000000000000;
	sram_mem[81568] = 16'b0000000000000000;
	sram_mem[81569] = 16'b0000000000000000;
	sram_mem[81570] = 16'b0000000000000000;
	sram_mem[81571] = 16'b0000000000000000;
	sram_mem[81572] = 16'b0000000000000000;
	sram_mem[81573] = 16'b0000000000000000;
	sram_mem[81574] = 16'b0000000000000000;
	sram_mem[81575] = 16'b0000000000000000;
	sram_mem[81576] = 16'b0000000000000000;
	sram_mem[81577] = 16'b0000000000000000;
	sram_mem[81578] = 16'b0000000000000000;
	sram_mem[81579] = 16'b0000000000000000;
	sram_mem[81580] = 16'b0000000000000000;
	sram_mem[81581] = 16'b0000000000000000;
	sram_mem[81582] = 16'b0000000000000000;
	sram_mem[81583] = 16'b0000000000000000;
	sram_mem[81584] = 16'b0000000000000000;
	sram_mem[81585] = 16'b0000000000000000;
	sram_mem[81586] = 16'b0000000000000000;
	sram_mem[81587] = 16'b0000000000000000;
	sram_mem[81588] = 16'b0000000000000000;
	sram_mem[81589] = 16'b0000000000000000;
	sram_mem[81590] = 16'b0000000000000000;
	sram_mem[81591] = 16'b0000000000000000;
	sram_mem[81592] = 16'b0000000000000000;
	sram_mem[81593] = 16'b0000000000000000;
	sram_mem[81594] = 16'b0000000000000000;
	sram_mem[81595] = 16'b0000000000000000;
	sram_mem[81596] = 16'b0000000000000000;
	sram_mem[81597] = 16'b0000000000000000;
	sram_mem[81598] = 16'b0000000000000000;
	sram_mem[81599] = 16'b0000000000000000;
	sram_mem[81600] = 16'b0000000000000000;
	sram_mem[81601] = 16'b0000000000000000;
	sram_mem[81602] = 16'b0000000000000000;
	sram_mem[81603] = 16'b0000000000000000;
	sram_mem[81604] = 16'b0000000000000000;
	sram_mem[81605] = 16'b0000000000000000;
	sram_mem[81606] = 16'b0000000000000000;
	sram_mem[81607] = 16'b0000000000000000;
	sram_mem[81608] = 16'b0000000000000000;
	sram_mem[81609] = 16'b0000000000000000;
	sram_mem[81610] = 16'b0000000000000000;
	sram_mem[81611] = 16'b0000000000000000;
	sram_mem[81612] = 16'b0000000000000000;
	sram_mem[81613] = 16'b0000000000000000;
	sram_mem[81614] = 16'b0000000000000000;
	sram_mem[81615] = 16'b0000000000000000;
	sram_mem[81616] = 16'b0000000000000000;
	sram_mem[81617] = 16'b0000000000000000;
	sram_mem[81618] = 16'b0000000000000000;
	sram_mem[81619] = 16'b0000000000000000;
	sram_mem[81620] = 16'b0000000000000000;
	sram_mem[81621] = 16'b0000000000000000;
	sram_mem[81622] = 16'b0000000000000000;
	sram_mem[81623] = 16'b0000000000000000;
	sram_mem[81624] = 16'b0000000000000000;
	sram_mem[81625] = 16'b0000000000000000;
	sram_mem[81626] = 16'b0000000000000000;
	sram_mem[81627] = 16'b0000000000000000;
	sram_mem[81628] = 16'b0000000000000000;
	sram_mem[81629] = 16'b0000000000000000;
	sram_mem[81630] = 16'b0000000000000000;
	sram_mem[81631] = 16'b0000000000000000;
	sram_mem[81632] = 16'b0000000000000000;
	sram_mem[81633] = 16'b0000000000000000;
	sram_mem[81634] = 16'b0000000000000000;
	sram_mem[81635] = 16'b0000000000000000;
	sram_mem[81636] = 16'b0000000000000000;
	sram_mem[81637] = 16'b0000000000000000;
	sram_mem[81638] = 16'b0000000000000000;
	sram_mem[81639] = 16'b0000000000000000;
	sram_mem[81640] = 16'b0000000000000000;
	sram_mem[81641] = 16'b0000000000000000;
	sram_mem[81642] = 16'b0000000000000000;
	sram_mem[81643] = 16'b0000000000000000;
	sram_mem[81644] = 16'b0000000000000000;
	sram_mem[81645] = 16'b0000000000000000;
	sram_mem[81646] = 16'b0000000000000000;
	sram_mem[81647] = 16'b0000000000000000;
	sram_mem[81648] = 16'b0000000000000000;
	sram_mem[81649] = 16'b0000000000000000;
	sram_mem[81650] = 16'b0000000000000000;
	sram_mem[81651] = 16'b0000000000000000;
	sram_mem[81652] = 16'b0000000000000000;
	sram_mem[81653] = 16'b0000000000000000;
	sram_mem[81654] = 16'b0000000000000000;
	sram_mem[81655] = 16'b0000000000000000;
	sram_mem[81656] = 16'b0000000000000000;
	sram_mem[81657] = 16'b0000000000000000;
	sram_mem[81658] = 16'b0000000000000000;
	sram_mem[81659] = 16'b0000000000000000;
	sram_mem[81660] = 16'b0000000000000000;
	sram_mem[81661] = 16'b0000000000000000;
	sram_mem[81662] = 16'b0000000000000000;
	sram_mem[81663] = 16'b0000000000000000;
	sram_mem[81664] = 16'b0000000000000000;
	sram_mem[81665] = 16'b0000000000000000;
	sram_mem[81666] = 16'b0000000000000000;
	sram_mem[81667] = 16'b0000000000000000;
	sram_mem[81668] = 16'b0000000000000000;
	sram_mem[81669] = 16'b0000000000000000;
	sram_mem[81670] = 16'b0000000000000000;
	sram_mem[81671] = 16'b0000000000000000;
	sram_mem[81672] = 16'b0000000000000000;
	sram_mem[81673] = 16'b0000000000000000;
	sram_mem[81674] = 16'b0000000000000000;
	sram_mem[81675] = 16'b0000000000000000;
	sram_mem[81676] = 16'b0000000000000000;
	sram_mem[81677] = 16'b0000000000000000;
	sram_mem[81678] = 16'b0000000000000000;
	sram_mem[81679] = 16'b0000000000000000;
	sram_mem[81680] = 16'b0000000000000000;
	sram_mem[81681] = 16'b0000000000000000;
	sram_mem[81682] = 16'b0000000000000000;
	sram_mem[81683] = 16'b0000000000000000;
	sram_mem[81684] = 16'b0000000000000000;
	sram_mem[81685] = 16'b0000000000000000;
	sram_mem[81686] = 16'b0000000000000000;
	sram_mem[81687] = 16'b0000000000000000;
	sram_mem[81688] = 16'b0000000000000000;
	sram_mem[81689] = 16'b0000000000000000;
	sram_mem[81690] = 16'b0000000000000000;
	sram_mem[81691] = 16'b0000000000000000;
	sram_mem[81692] = 16'b0000000000000000;
	sram_mem[81693] = 16'b0000000000000000;
	sram_mem[81694] = 16'b0000000000000000;
	sram_mem[81695] = 16'b0000000000000000;
	sram_mem[81696] = 16'b0000000000000000;
	sram_mem[81697] = 16'b0000000000000000;
	sram_mem[81698] = 16'b0000000000000000;
	sram_mem[81699] = 16'b0000000000000000;
	sram_mem[81700] = 16'b0000000000000000;
	sram_mem[81701] = 16'b0000000000000000;
	sram_mem[81702] = 16'b0000000000000000;
	sram_mem[81703] = 16'b0000000000000000;
	sram_mem[81704] = 16'b0000000000000000;
	sram_mem[81705] = 16'b0000000000000000;
	sram_mem[81706] = 16'b0000000000000000;
	sram_mem[81707] = 16'b0000000000000000;
	sram_mem[81708] = 16'b0000000000000000;
	sram_mem[81709] = 16'b0000000000000000;
	sram_mem[81710] = 16'b0000000000000000;
	sram_mem[81711] = 16'b0000000000000000;
	sram_mem[81712] = 16'b0000000000000000;
	sram_mem[81713] = 16'b0000000000000000;
	sram_mem[81714] = 16'b0000000000000000;
	sram_mem[81715] = 16'b0000000000000000;
	sram_mem[81716] = 16'b0000000000000000;
	sram_mem[81717] = 16'b0000000000000000;
	sram_mem[81718] = 16'b0000000000000000;
	sram_mem[81719] = 16'b0000000000000000;
	sram_mem[81720] = 16'b0000000000000000;
	sram_mem[81721] = 16'b0000000000000000;
	sram_mem[81722] = 16'b0000000000000000;
	sram_mem[81723] = 16'b0000000000000000;
	sram_mem[81724] = 16'b0000000000000000;
	sram_mem[81725] = 16'b0000000000000000;
	sram_mem[81726] = 16'b0000000000000000;
	sram_mem[81727] = 16'b0000000000000000;
	sram_mem[81728] = 16'b0000000000000000;
	sram_mem[81729] = 16'b0000000000000000;
	sram_mem[81730] = 16'b0000000000000000;
	sram_mem[81731] = 16'b0000000000000000;
	sram_mem[81732] = 16'b0000000000000000;
	sram_mem[81733] = 16'b0000000000000000;
	sram_mem[81734] = 16'b0000000000000000;
	sram_mem[81735] = 16'b0000000000000000;
	sram_mem[81736] = 16'b0000000000000000;
	sram_mem[81737] = 16'b0000000000000000;
	sram_mem[81738] = 16'b0000000000000000;
	sram_mem[81739] = 16'b0000000000000000;
	sram_mem[81740] = 16'b0000000000000000;
	sram_mem[81741] = 16'b0000000000000000;
	sram_mem[81742] = 16'b0000000000000000;
	sram_mem[81743] = 16'b0000000000000000;
	sram_mem[81744] = 16'b0000000000000000;
	sram_mem[81745] = 16'b0000000000000000;
	sram_mem[81746] = 16'b0000000000000000;
	sram_mem[81747] = 16'b0000000000000000;
	sram_mem[81748] = 16'b0000000000000000;
	sram_mem[81749] = 16'b0000000000000000;
	sram_mem[81750] = 16'b0000000000000000;
	sram_mem[81751] = 16'b0000000000000000;
	sram_mem[81752] = 16'b0000000000000000;
	sram_mem[81753] = 16'b0000000000000000;
	sram_mem[81754] = 16'b0000000000000000;
	sram_mem[81755] = 16'b0000000000000000;
	sram_mem[81756] = 16'b0000000000000000;
	sram_mem[81757] = 16'b0000000000000000;
	sram_mem[81758] = 16'b0000000000000000;
	sram_mem[81759] = 16'b0000000000000000;
	sram_mem[81760] = 16'b0000000000000000;
	sram_mem[81761] = 16'b0000000000000000;
	sram_mem[81762] = 16'b0000000000000000;
	sram_mem[81763] = 16'b0000000000000000;
	sram_mem[81764] = 16'b0000000000000000;
	sram_mem[81765] = 16'b0000000000000000;
	sram_mem[81766] = 16'b0000000000000000;
	sram_mem[81767] = 16'b0000000000000000;
	sram_mem[81768] = 16'b0000000000000000;
	sram_mem[81769] = 16'b0000000000000000;
	sram_mem[81770] = 16'b0000000000000000;
	sram_mem[81771] = 16'b0000000000000000;
	sram_mem[81772] = 16'b0000000000000000;
	sram_mem[81773] = 16'b0000000000000000;
	sram_mem[81774] = 16'b0000000000000000;
	sram_mem[81775] = 16'b0000000000000000;
	sram_mem[81776] = 16'b0000000000000000;
	sram_mem[81777] = 16'b0000000000000000;
	sram_mem[81778] = 16'b0000000000000000;
	sram_mem[81779] = 16'b0000000000000000;
	sram_mem[81780] = 16'b0000000000000000;
	sram_mem[81781] = 16'b0000000000000000;
	sram_mem[81782] = 16'b0000000000000000;
	sram_mem[81783] = 16'b0000000000000000;
	sram_mem[81784] = 16'b0000000000000000;
	sram_mem[81785] = 16'b0000000000000000;
	sram_mem[81786] = 16'b0000000000000000;
	sram_mem[81787] = 16'b0000000000000000;
	sram_mem[81788] = 16'b0000000000000000;
	sram_mem[81789] = 16'b0000000000000000;
	sram_mem[81790] = 16'b0000000000000000;
	sram_mem[81791] = 16'b0000000000000000;
	sram_mem[81792] = 16'b0000000000000000;
	sram_mem[81793] = 16'b0000000000000000;
	sram_mem[81794] = 16'b0000000000000000;
	sram_mem[81795] = 16'b0000000000000000;
	sram_mem[81796] = 16'b0000000000000000;
	sram_mem[81797] = 16'b0000000000000000;
	sram_mem[81798] = 16'b0000000000000000;
	sram_mem[81799] = 16'b0000000000000000;
	sram_mem[81800] = 16'b0000000000000000;
	sram_mem[81801] = 16'b0000000000000000;
	sram_mem[81802] = 16'b0000000000000000;
	sram_mem[81803] = 16'b0000000000000000;
	sram_mem[81804] = 16'b0000000000000000;
	sram_mem[81805] = 16'b0000000000000000;
	sram_mem[81806] = 16'b0000000000000000;
	sram_mem[81807] = 16'b0000000000000000;
	sram_mem[81808] = 16'b0000000000000000;
	sram_mem[81809] = 16'b0000000000000000;
	sram_mem[81810] = 16'b0000000000000000;
	sram_mem[81811] = 16'b0000000000000000;
	sram_mem[81812] = 16'b0000000000000000;
	sram_mem[81813] = 16'b0000000000000000;
	sram_mem[81814] = 16'b0000000000000000;
	sram_mem[81815] = 16'b0000000000000000;
	sram_mem[81816] = 16'b0000000000000000;
	sram_mem[81817] = 16'b0000000000000000;
	sram_mem[81818] = 16'b0000000000000000;
	sram_mem[81819] = 16'b0000000000000000;
	sram_mem[81820] = 16'b0000000000000000;
	sram_mem[81821] = 16'b0000000000000000;
	sram_mem[81822] = 16'b0000000000000000;
	sram_mem[81823] = 16'b0000000000000000;
	sram_mem[81824] = 16'b0000000000000000;
	sram_mem[81825] = 16'b0000000000000000;
	sram_mem[81826] = 16'b0000000000000000;
	sram_mem[81827] = 16'b0000000000000000;
	sram_mem[81828] = 16'b0000000000000000;
	sram_mem[81829] = 16'b0000000000000000;
	sram_mem[81830] = 16'b0000000000000000;
	sram_mem[81831] = 16'b0000000000000000;
	sram_mem[81832] = 16'b0000000000000000;
	sram_mem[81833] = 16'b0000000000000000;
	sram_mem[81834] = 16'b0000000000000000;
	sram_mem[81835] = 16'b0000000000000000;
	sram_mem[81836] = 16'b0000000000000000;
	sram_mem[81837] = 16'b0000000000000000;
	sram_mem[81838] = 16'b0000000000000000;
	sram_mem[81839] = 16'b0000000000000000;
	sram_mem[81840] = 16'b0000000000000000;
	sram_mem[81841] = 16'b0000000000000000;
	sram_mem[81842] = 16'b0000000000000000;
	sram_mem[81843] = 16'b0000000000000000;
	sram_mem[81844] = 16'b0000000000000000;
	sram_mem[81845] = 16'b0000000000000000;
	sram_mem[81846] = 16'b0000000000000000;
	sram_mem[81847] = 16'b0000000000000000;
	sram_mem[81848] = 16'b0000000000000000;
	sram_mem[81849] = 16'b0000000000000000;
	sram_mem[81850] = 16'b0000000000000000;
	sram_mem[81851] = 16'b0000000000000000;
	sram_mem[81852] = 16'b0000000000000000;
	sram_mem[81853] = 16'b0000000000000000;
	sram_mem[81854] = 16'b0000000000000000;
	sram_mem[81855] = 16'b0000000000000000;
	sram_mem[81856] = 16'b0000000000000000;
	sram_mem[81857] = 16'b0000000000000000;
	sram_mem[81858] = 16'b0000000000000000;
	sram_mem[81859] = 16'b0000000000000000;
	sram_mem[81860] = 16'b0000000000000000;
	sram_mem[81861] = 16'b0000000000000000;
	sram_mem[81862] = 16'b0000000000000000;
	sram_mem[81863] = 16'b0000000000000000;
	sram_mem[81864] = 16'b0000000000000000;
	sram_mem[81865] = 16'b0000000000000000;
	sram_mem[81866] = 16'b0000000000000000;
	sram_mem[81867] = 16'b0000000000000000;
	sram_mem[81868] = 16'b0000000000000000;
	sram_mem[81869] = 16'b0000000000000000;
	sram_mem[81870] = 16'b0000000000000000;
	sram_mem[81871] = 16'b0000000000000000;
	sram_mem[81872] = 16'b0000000000000000;
	sram_mem[81873] = 16'b0000000000000000;
	sram_mem[81874] = 16'b0000000000000000;
	sram_mem[81875] = 16'b0000000000000000;
	sram_mem[81876] = 16'b0000000000000000;
	sram_mem[81877] = 16'b0000000000000000;
	sram_mem[81878] = 16'b0000000000000000;
	sram_mem[81879] = 16'b0000000000000000;
	sram_mem[81880] = 16'b0000000000000000;
	sram_mem[81881] = 16'b0000000000000000;
	sram_mem[81882] = 16'b0000000000000000;
	sram_mem[81883] = 16'b0000000000000000;
	sram_mem[81884] = 16'b0000000000000000;
	sram_mem[81885] = 16'b0000000000000000;
	sram_mem[81886] = 16'b0000000000000000;
	sram_mem[81887] = 16'b0000000000000000;
	sram_mem[81888] = 16'b0000000000000000;
	sram_mem[81889] = 16'b0000000000000000;
	sram_mem[81890] = 16'b0000000000000000;
	sram_mem[81891] = 16'b0000000000000000;
	sram_mem[81892] = 16'b0000000000000000;
	sram_mem[81893] = 16'b0000000000000000;
	sram_mem[81894] = 16'b0000000000000000;
	sram_mem[81895] = 16'b0000000000000000;
	sram_mem[81896] = 16'b0000000000000000;
	sram_mem[81897] = 16'b0000000000000000;
	sram_mem[81898] = 16'b0000000000000000;
	sram_mem[81899] = 16'b0000000000000000;
	sram_mem[81900] = 16'b0000000000000000;
	sram_mem[81901] = 16'b0000000000000000;
	sram_mem[81902] = 16'b0000000000000000;
	sram_mem[81903] = 16'b0000000000000000;
	sram_mem[81904] = 16'b0000000000000000;
	sram_mem[81905] = 16'b0000000000000000;
	sram_mem[81906] = 16'b0000000000000000;
	sram_mem[81907] = 16'b0000000000000000;
	sram_mem[81908] = 16'b0000000000000000;
	sram_mem[81909] = 16'b0000000000000000;
	sram_mem[81910] = 16'b0000000000000000;
	sram_mem[81911] = 16'b0000000000000000;
	sram_mem[81912] = 16'b0000000000000000;
	sram_mem[81913] = 16'b0000000000000000;
	sram_mem[81914] = 16'b0000000000000000;
	sram_mem[81915] = 16'b0000000000000000;
	sram_mem[81916] = 16'b0000000000000000;
	sram_mem[81917] = 16'b0000000000000000;
	sram_mem[81918] = 16'b0000000000000000;
	sram_mem[81919] = 16'b0000000000000000;
	sram_mem[81920] = 16'b0000000000000000;
	sram_mem[81921] = 16'b0000000000000000;
	sram_mem[81922] = 16'b0000000000000000;
	sram_mem[81923] = 16'b0000000000000000;
	sram_mem[81924] = 16'b0000000000000000;
	sram_mem[81925] = 16'b0000000000000000;
	sram_mem[81926] = 16'b0000000000000000;
	sram_mem[81927] = 16'b0000000000000000;
	sram_mem[81928] = 16'b0000000000000000;
	sram_mem[81929] = 16'b0000000000000000;
	sram_mem[81930] = 16'b0000000000000000;
	sram_mem[81931] = 16'b0000000000000000;
	sram_mem[81932] = 16'b0000000000000000;
	sram_mem[81933] = 16'b0000000000000000;
	sram_mem[81934] = 16'b0000000000000000;
	sram_mem[81935] = 16'b0000000000000000;
	sram_mem[81936] = 16'b0000000000000000;
	sram_mem[81937] = 16'b0000000000000000;
	sram_mem[81938] = 16'b0000000000000000;
	sram_mem[81939] = 16'b0000000000000000;
	sram_mem[81940] = 16'b0000000000000000;
	sram_mem[81941] = 16'b0000000000000000;
	sram_mem[81942] = 16'b0000000000000000;
	sram_mem[81943] = 16'b0000000000000000;
	sram_mem[81944] = 16'b0000000000000000;
	sram_mem[81945] = 16'b0000000000000000;
	sram_mem[81946] = 16'b0000000000000000;
	sram_mem[81947] = 16'b0000000000000000;
	sram_mem[81948] = 16'b0000000000000000;
	sram_mem[81949] = 16'b0000000000000000;
	sram_mem[81950] = 16'b0000000000000000;
	sram_mem[81951] = 16'b0000000000000000;
	sram_mem[81952] = 16'b0000000000000000;
	sram_mem[81953] = 16'b0000000000000000;
	sram_mem[81954] = 16'b0000000000000000;
	sram_mem[81955] = 16'b0000000000000000;
	sram_mem[81956] = 16'b0000000000000000;
	sram_mem[81957] = 16'b0000000000000000;
	sram_mem[81958] = 16'b0000000000000000;
	sram_mem[81959] = 16'b0000000000000000;
	sram_mem[81960] = 16'b0000000000000000;
	sram_mem[81961] = 16'b0000000000000000;
	sram_mem[81962] = 16'b0000000000000000;
	sram_mem[81963] = 16'b0000000000000000;
	sram_mem[81964] = 16'b0000000000000000;
	sram_mem[81965] = 16'b0000000000000000;
	sram_mem[81966] = 16'b0000000000000000;
	sram_mem[81967] = 16'b0000000000000000;
	sram_mem[81968] = 16'b0000000000000000;
	sram_mem[81969] = 16'b0000000000000000;
	sram_mem[81970] = 16'b0000000000000000;
	sram_mem[81971] = 16'b0000000000000000;
	sram_mem[81972] = 16'b0000000000000000;
	sram_mem[81973] = 16'b0000000000000000;
	sram_mem[81974] = 16'b0000000000000000;
	sram_mem[81975] = 16'b0000000000000000;
	sram_mem[81976] = 16'b0000000000000000;
	sram_mem[81977] = 16'b0000000000000000;
	sram_mem[81978] = 16'b0000000000000000;
	sram_mem[81979] = 16'b0000000000000000;
	sram_mem[81980] = 16'b0000000000000000;
	sram_mem[81981] = 16'b0000000000000000;
	sram_mem[81982] = 16'b0000000000000000;
	sram_mem[81983] = 16'b0000000000000000;
	sram_mem[81984] = 16'b0000000000000000;
	sram_mem[81985] = 16'b0000000000000000;
	sram_mem[81986] = 16'b0000000000000000;
	sram_mem[81987] = 16'b0000000000000000;
	sram_mem[81988] = 16'b0000000000000000;
	sram_mem[81989] = 16'b0000000000000000;
	sram_mem[81990] = 16'b0000000000000000;
	sram_mem[81991] = 16'b0000000000000000;
	sram_mem[81992] = 16'b0000000000000000;
	sram_mem[81993] = 16'b0000000000000000;
	sram_mem[81994] = 16'b0000000000000000;
	sram_mem[81995] = 16'b0000000000000000;
	sram_mem[81996] = 16'b0000000000000000;
	sram_mem[81997] = 16'b0000000000000000;
	sram_mem[81998] = 16'b0000000000000000;
	sram_mem[81999] = 16'b0000000000000000;
	sram_mem[82000] = 16'b0000000000000000;
	sram_mem[82001] = 16'b0000000000000000;
	sram_mem[82002] = 16'b0000000000000000;
	sram_mem[82003] = 16'b0000000000000000;
	sram_mem[82004] = 16'b0000000000000000;
	sram_mem[82005] = 16'b0000000000000000;
	sram_mem[82006] = 16'b0000000000000000;
	sram_mem[82007] = 16'b0000000000000000;
	sram_mem[82008] = 16'b0000000000000000;
	sram_mem[82009] = 16'b0000000000000000;
	sram_mem[82010] = 16'b0000000000000000;
	sram_mem[82011] = 16'b0000000000000000;
	sram_mem[82012] = 16'b0000000000000000;
	sram_mem[82013] = 16'b0000000000000000;
	sram_mem[82014] = 16'b0000000000000000;
	sram_mem[82015] = 16'b0000000000000000;
	sram_mem[82016] = 16'b0000000000000000;
	sram_mem[82017] = 16'b0000000000000000;
	sram_mem[82018] = 16'b0000000000000000;
	sram_mem[82019] = 16'b0000000000000000;
	sram_mem[82020] = 16'b0000000000000000;
	sram_mem[82021] = 16'b0000000000000000;
	sram_mem[82022] = 16'b0000000000000000;
	sram_mem[82023] = 16'b0000000000000000;
	sram_mem[82024] = 16'b0000000000000000;
	sram_mem[82025] = 16'b0000000000000000;
	sram_mem[82026] = 16'b0000000000000000;
	sram_mem[82027] = 16'b0000000000000000;
	sram_mem[82028] = 16'b0000000000000000;
	sram_mem[82029] = 16'b0000000000000000;
	sram_mem[82030] = 16'b0000000000000000;
	sram_mem[82031] = 16'b0000000000000000;
	sram_mem[82032] = 16'b0000000000000000;
	sram_mem[82033] = 16'b0000000000000000;
	sram_mem[82034] = 16'b0000000000000000;
	sram_mem[82035] = 16'b0000000000000000;
	sram_mem[82036] = 16'b0000000000000000;
	sram_mem[82037] = 16'b0000000000000000;
	sram_mem[82038] = 16'b0000000000000000;
	sram_mem[82039] = 16'b0000000000000000;
	sram_mem[82040] = 16'b0000000000000000;
	sram_mem[82041] = 16'b0000000000000000;
	sram_mem[82042] = 16'b0000000000000000;
	sram_mem[82043] = 16'b0000000000000000;
	sram_mem[82044] = 16'b0000000000000000;
	sram_mem[82045] = 16'b0000000000000000;
	sram_mem[82046] = 16'b0000000000000000;
	sram_mem[82047] = 16'b0000000000000000;
	sram_mem[82048] = 16'b0000000000000000;
	sram_mem[82049] = 16'b0000000000000000;
	sram_mem[82050] = 16'b0000000000000000;
	sram_mem[82051] = 16'b0000000000000000;
	sram_mem[82052] = 16'b0000000000000000;
	sram_mem[82053] = 16'b0000000000000000;
	sram_mem[82054] = 16'b0000000000000000;
	sram_mem[82055] = 16'b0000000000000000;
	sram_mem[82056] = 16'b0000000000000000;
	sram_mem[82057] = 16'b0000000000000000;
	sram_mem[82058] = 16'b0000000000000000;
	sram_mem[82059] = 16'b0000000000000000;
	sram_mem[82060] = 16'b0000000000000000;
	sram_mem[82061] = 16'b0000000000000000;
	sram_mem[82062] = 16'b0000000000000000;
	sram_mem[82063] = 16'b0000000000000000;
	sram_mem[82064] = 16'b0000000000000000;
	sram_mem[82065] = 16'b0000000000000000;
	sram_mem[82066] = 16'b0000000000000000;
	sram_mem[82067] = 16'b0000000000000000;
	sram_mem[82068] = 16'b0000000000000000;
	sram_mem[82069] = 16'b0000000000000000;
	sram_mem[82070] = 16'b0000000000000000;
	sram_mem[82071] = 16'b0000000000000000;
	sram_mem[82072] = 16'b0000000000000000;
	sram_mem[82073] = 16'b0000000000000000;
	sram_mem[82074] = 16'b0000000000000000;
	sram_mem[82075] = 16'b0000000000000000;
	sram_mem[82076] = 16'b0000000000000000;
	sram_mem[82077] = 16'b0000000000000000;
	sram_mem[82078] = 16'b0000000000000000;
	sram_mem[82079] = 16'b0000000000000000;
	sram_mem[82080] = 16'b0000000000000000;
	sram_mem[82081] = 16'b0000000000000000;
	sram_mem[82082] = 16'b0000000000000000;
	sram_mem[82083] = 16'b0000000000000000;
	sram_mem[82084] = 16'b0000000000000000;
	sram_mem[82085] = 16'b0000000000000000;
	sram_mem[82086] = 16'b0000000000000000;
	sram_mem[82087] = 16'b0000000000000000;
	sram_mem[82088] = 16'b0000000000000000;
	sram_mem[82089] = 16'b0000000000000000;
	sram_mem[82090] = 16'b0000000000000000;
	sram_mem[82091] = 16'b0000000000000000;
	sram_mem[82092] = 16'b0000000000000000;
	sram_mem[82093] = 16'b0000000000000000;
	sram_mem[82094] = 16'b0000000000000000;
	sram_mem[82095] = 16'b0000000000000000;
	sram_mem[82096] = 16'b0000000000000000;
	sram_mem[82097] = 16'b0000000000000000;
	sram_mem[82098] = 16'b0000000000000000;
	sram_mem[82099] = 16'b0000000000000000;
	sram_mem[82100] = 16'b0000000000000000;
	sram_mem[82101] = 16'b0000000000000000;
	sram_mem[82102] = 16'b0000000000000000;
	sram_mem[82103] = 16'b0000000000000000;
	sram_mem[82104] = 16'b0000000000000000;
	sram_mem[82105] = 16'b0000000000000000;
	sram_mem[82106] = 16'b0000000000000000;
	sram_mem[82107] = 16'b0000000000000000;
	sram_mem[82108] = 16'b0000000000000000;
	sram_mem[82109] = 16'b0000000000000000;
	sram_mem[82110] = 16'b0000000000000000;
	sram_mem[82111] = 16'b0000000000000000;
	sram_mem[82112] = 16'b0000000000000000;
	sram_mem[82113] = 16'b0000000000000000;
	sram_mem[82114] = 16'b0000000000000000;
	sram_mem[82115] = 16'b0000000000000000;
	sram_mem[82116] = 16'b0000000000000000;
	sram_mem[82117] = 16'b0000000000000000;
	sram_mem[82118] = 16'b0000000000000000;
	sram_mem[82119] = 16'b0000000000000000;
	sram_mem[82120] = 16'b0000000000000000;
	sram_mem[82121] = 16'b0000000000000000;
	sram_mem[82122] = 16'b0000000000000000;
	sram_mem[82123] = 16'b0000000000000000;
	sram_mem[82124] = 16'b0000000000000000;
	sram_mem[82125] = 16'b0000000000000000;
	sram_mem[82126] = 16'b0000000000000000;
	sram_mem[82127] = 16'b0000000000000000;
	sram_mem[82128] = 16'b0000000000000000;
	sram_mem[82129] = 16'b0000000000000000;
	sram_mem[82130] = 16'b0000000000000000;
	sram_mem[82131] = 16'b0000000000000000;
	sram_mem[82132] = 16'b0000000000000000;
	sram_mem[82133] = 16'b0000000000000000;
	sram_mem[82134] = 16'b0000000000000000;
	sram_mem[82135] = 16'b0000000000000000;
	sram_mem[82136] = 16'b0000000000000000;
	sram_mem[82137] = 16'b0000000000000000;
	sram_mem[82138] = 16'b0000000000000000;
	sram_mem[82139] = 16'b0000000000000000;
	sram_mem[82140] = 16'b0000000000000000;
	sram_mem[82141] = 16'b0000000000000000;
	sram_mem[82142] = 16'b0000000000000000;
	sram_mem[82143] = 16'b0000000000000000;
	sram_mem[82144] = 16'b0000000000000000;
	sram_mem[82145] = 16'b0000000000000000;
	sram_mem[82146] = 16'b0000000000000000;
	sram_mem[82147] = 16'b0000000000000000;
	sram_mem[82148] = 16'b0000000000000000;
	sram_mem[82149] = 16'b0000000000000000;
	sram_mem[82150] = 16'b0000000000000000;
	sram_mem[82151] = 16'b0000000000000000;
	sram_mem[82152] = 16'b0000000000000000;
	sram_mem[82153] = 16'b0000000000000000;
	sram_mem[82154] = 16'b0000000000000000;
	sram_mem[82155] = 16'b0000000000000000;
	sram_mem[82156] = 16'b0000000000000000;
	sram_mem[82157] = 16'b0000000000000000;
	sram_mem[82158] = 16'b0000000000000000;
	sram_mem[82159] = 16'b0000000000000000;
	sram_mem[82160] = 16'b0000000000000000;
	sram_mem[82161] = 16'b0000000000000000;
	sram_mem[82162] = 16'b0000000000000000;
	sram_mem[82163] = 16'b0000000000000000;
	sram_mem[82164] = 16'b0000000000000000;
	sram_mem[82165] = 16'b0000000000000000;
	sram_mem[82166] = 16'b0000000000000000;
	sram_mem[82167] = 16'b0000000000000000;
	sram_mem[82168] = 16'b0000000000000000;
	sram_mem[82169] = 16'b0000000000000000;
	sram_mem[82170] = 16'b0000000000000000;
	sram_mem[82171] = 16'b0000000000000000;
	sram_mem[82172] = 16'b0000000000000000;
	sram_mem[82173] = 16'b0000000000000000;
	sram_mem[82174] = 16'b0000000000000000;
	sram_mem[82175] = 16'b0000000000000000;
	sram_mem[82176] = 16'b0000000000000000;
	sram_mem[82177] = 16'b0000000000000000;
	sram_mem[82178] = 16'b0000000000000000;
	sram_mem[82179] = 16'b0000000000000000;
	sram_mem[82180] = 16'b0000000000000000;
	sram_mem[82181] = 16'b0000000000000000;
	sram_mem[82182] = 16'b0000000000000000;
	sram_mem[82183] = 16'b0000000000000000;
	sram_mem[82184] = 16'b0000000000000000;
	sram_mem[82185] = 16'b0000000000000000;
	sram_mem[82186] = 16'b0000000000000000;
	sram_mem[82187] = 16'b0000000000000000;
	sram_mem[82188] = 16'b0000000000000000;
	sram_mem[82189] = 16'b0000000000000000;
	sram_mem[82190] = 16'b0000000000000000;
	sram_mem[82191] = 16'b0000000000000000;
	sram_mem[82192] = 16'b0000000000000000;
	sram_mem[82193] = 16'b0000000000000000;
	sram_mem[82194] = 16'b0000000000000000;
	sram_mem[82195] = 16'b0000000000000000;
	sram_mem[82196] = 16'b0000000000000000;
	sram_mem[82197] = 16'b0000000000000000;
	sram_mem[82198] = 16'b0000000000000000;
	sram_mem[82199] = 16'b0000000000000000;
	sram_mem[82200] = 16'b0000000000000000;
	sram_mem[82201] = 16'b0000000000000000;
	sram_mem[82202] = 16'b0000000000000000;
	sram_mem[82203] = 16'b0000000000000000;
	sram_mem[82204] = 16'b0000000000000000;
	sram_mem[82205] = 16'b0000000000000000;
	sram_mem[82206] = 16'b0000000000000000;
	sram_mem[82207] = 16'b0000000000000000;
	sram_mem[82208] = 16'b0000000000000000;
	sram_mem[82209] = 16'b0000000000000000;
	sram_mem[82210] = 16'b0000000000000000;
	sram_mem[82211] = 16'b0000000000000000;
	sram_mem[82212] = 16'b0000000000000000;
	sram_mem[82213] = 16'b0000000000000000;
	sram_mem[82214] = 16'b0000000000000000;
	sram_mem[82215] = 16'b0000000000000000;
	sram_mem[82216] = 16'b0000000000000000;
	sram_mem[82217] = 16'b0000000000000000;
	sram_mem[82218] = 16'b0000000000000000;
	sram_mem[82219] = 16'b0000000000000000;
	sram_mem[82220] = 16'b0000000000000000;
	sram_mem[82221] = 16'b0000000000000000;
	sram_mem[82222] = 16'b0000000000000000;
	sram_mem[82223] = 16'b0000000000000000;
	sram_mem[82224] = 16'b0000000000000000;
	sram_mem[82225] = 16'b0000000000000000;
	sram_mem[82226] = 16'b0000000000000000;
	sram_mem[82227] = 16'b0000000000000000;
	sram_mem[82228] = 16'b0000000000000000;
	sram_mem[82229] = 16'b0000000000000000;
	sram_mem[82230] = 16'b0000000000000000;
	sram_mem[82231] = 16'b0000000000000000;
	sram_mem[82232] = 16'b0000000000000000;
	sram_mem[82233] = 16'b0000000000000000;
	sram_mem[82234] = 16'b0000000000000000;
	sram_mem[82235] = 16'b0000000000000000;
	sram_mem[82236] = 16'b0000000000000000;
	sram_mem[82237] = 16'b0000000000000000;
	sram_mem[82238] = 16'b0000000000000000;
	sram_mem[82239] = 16'b0000000000000000;
	sram_mem[82240] = 16'b0000000000000000;
	sram_mem[82241] = 16'b0000000000000000;
	sram_mem[82242] = 16'b0000000000000000;
	sram_mem[82243] = 16'b0000000000000000;
	sram_mem[82244] = 16'b0000000000000000;
	sram_mem[82245] = 16'b0000000000000000;
	sram_mem[82246] = 16'b0000000000000000;
	sram_mem[82247] = 16'b0000000000000000;
	sram_mem[82248] = 16'b0000000000000000;
	sram_mem[82249] = 16'b0000000000000000;
	sram_mem[82250] = 16'b0000000000000000;
	sram_mem[82251] = 16'b0000000000000000;
	sram_mem[82252] = 16'b0000000000000000;
	sram_mem[82253] = 16'b0000000000000000;
	sram_mem[82254] = 16'b0000000000000000;
	sram_mem[82255] = 16'b0000000000000000;
	sram_mem[82256] = 16'b0000000000000000;
	sram_mem[82257] = 16'b0000000000000000;
	sram_mem[82258] = 16'b0000000000000000;
	sram_mem[82259] = 16'b0000000000000000;
	sram_mem[82260] = 16'b0000000000000000;
	sram_mem[82261] = 16'b0000000000000000;
	sram_mem[82262] = 16'b0000000000000000;
	sram_mem[82263] = 16'b0000000000000000;
	sram_mem[82264] = 16'b0000000000000000;
	sram_mem[82265] = 16'b0000000000000000;
	sram_mem[82266] = 16'b0000000000000000;
	sram_mem[82267] = 16'b0000000000000000;
	sram_mem[82268] = 16'b0000000000000000;
	sram_mem[82269] = 16'b0000000000000000;
	sram_mem[82270] = 16'b0000000000000000;
	sram_mem[82271] = 16'b0000000000000000;
	sram_mem[82272] = 16'b0000000000000000;
	sram_mem[82273] = 16'b0000000000000000;
	sram_mem[82274] = 16'b0000000000000000;
	sram_mem[82275] = 16'b0000000000000000;
	sram_mem[82276] = 16'b0000000000000000;
	sram_mem[82277] = 16'b0000000000000000;
	sram_mem[82278] = 16'b0000000000000000;
	sram_mem[82279] = 16'b0000000000000000;
	sram_mem[82280] = 16'b0000000000000000;
	sram_mem[82281] = 16'b0000000000000000;
	sram_mem[82282] = 16'b0000000000000000;
	sram_mem[82283] = 16'b0000000000000000;
	sram_mem[82284] = 16'b0000000000000000;
	sram_mem[82285] = 16'b0000000000000000;
	sram_mem[82286] = 16'b0000000000000000;
	sram_mem[82287] = 16'b0000000000000000;
	sram_mem[82288] = 16'b0000000000000000;
	sram_mem[82289] = 16'b0000000000000000;
	sram_mem[82290] = 16'b0000000000000000;
	sram_mem[82291] = 16'b0000000000000000;
	sram_mem[82292] = 16'b0000000000000000;
	sram_mem[82293] = 16'b0000000000000000;
	sram_mem[82294] = 16'b0000000000000000;
	sram_mem[82295] = 16'b0000000000000000;
	sram_mem[82296] = 16'b0000000000000000;
	sram_mem[82297] = 16'b0000000000000000;
	sram_mem[82298] = 16'b0000000000000000;
	sram_mem[82299] = 16'b0000000000000000;
	sram_mem[82300] = 16'b0000000000000000;
	sram_mem[82301] = 16'b0000000000000000;
	sram_mem[82302] = 16'b0000000000000000;
	sram_mem[82303] = 16'b0000000000000000;
	sram_mem[82304] = 16'b0000000000000000;
	sram_mem[82305] = 16'b0000000000000000;
	sram_mem[82306] = 16'b0000000000000000;
	sram_mem[82307] = 16'b0000000000000000;
	sram_mem[82308] = 16'b0000000000000000;
	sram_mem[82309] = 16'b0000000000000000;
	sram_mem[82310] = 16'b0000000000000000;
	sram_mem[82311] = 16'b0000000000000000;
	sram_mem[82312] = 16'b0000000000000000;
	sram_mem[82313] = 16'b0000000000000000;
	sram_mem[82314] = 16'b0000000000000000;
	sram_mem[82315] = 16'b0000000000000000;
	sram_mem[82316] = 16'b0000000000000000;
	sram_mem[82317] = 16'b0000000000000000;
	sram_mem[82318] = 16'b0000000000000000;
	sram_mem[82319] = 16'b0000000000000000;
	sram_mem[82320] = 16'b0000000000000000;
	sram_mem[82321] = 16'b0000000000000000;
	sram_mem[82322] = 16'b0000000000000000;
	sram_mem[82323] = 16'b0000000000000000;
	sram_mem[82324] = 16'b0000000000000000;
	sram_mem[82325] = 16'b0000000000000000;
	sram_mem[82326] = 16'b0000000000000000;
	sram_mem[82327] = 16'b0000000000000000;
	sram_mem[82328] = 16'b0000000000000000;
	sram_mem[82329] = 16'b0000000000000000;
	sram_mem[82330] = 16'b0000000000000000;
	sram_mem[82331] = 16'b0000000000000000;
	sram_mem[82332] = 16'b0000000000000000;
	sram_mem[82333] = 16'b0000000000000000;
	sram_mem[82334] = 16'b0000000000000000;
	sram_mem[82335] = 16'b0000000000000000;
	sram_mem[82336] = 16'b0000000000000000;
	sram_mem[82337] = 16'b0000000000000000;
	sram_mem[82338] = 16'b0000000000000000;
	sram_mem[82339] = 16'b0000000000000000;
	sram_mem[82340] = 16'b0000000000000000;
	sram_mem[82341] = 16'b0000000000000000;
	sram_mem[82342] = 16'b0000000000000000;
	sram_mem[82343] = 16'b0000000000000000;
	sram_mem[82344] = 16'b0000000000000000;
	sram_mem[82345] = 16'b0000000000000000;
	sram_mem[82346] = 16'b0000000000000000;
	sram_mem[82347] = 16'b0000000000000000;
	sram_mem[82348] = 16'b0000000000000000;
	sram_mem[82349] = 16'b0000000000000000;
	sram_mem[82350] = 16'b0000000000000000;
	sram_mem[82351] = 16'b0000000000000000;
	sram_mem[82352] = 16'b0000000000000000;
	sram_mem[82353] = 16'b0000000000000000;
	sram_mem[82354] = 16'b0000000000000000;
	sram_mem[82355] = 16'b0000000000000000;
	sram_mem[82356] = 16'b0000000000000000;
	sram_mem[82357] = 16'b0000000000000000;
	sram_mem[82358] = 16'b0000000000000000;
	sram_mem[82359] = 16'b0000000000000000;
	sram_mem[82360] = 16'b0000000000000000;
	sram_mem[82361] = 16'b0000000000000000;
	sram_mem[82362] = 16'b0000000000000000;
	sram_mem[82363] = 16'b0000000000000000;
	sram_mem[82364] = 16'b0000000000000000;
	sram_mem[82365] = 16'b0000000000000000;
	sram_mem[82366] = 16'b0000000000000000;
	sram_mem[82367] = 16'b0000000000000000;
	sram_mem[82368] = 16'b0000000000000000;
	sram_mem[82369] = 16'b0000000000000000;
	sram_mem[82370] = 16'b0000000000000000;
	sram_mem[82371] = 16'b0000000000000000;
	sram_mem[82372] = 16'b0000000000000000;
	sram_mem[82373] = 16'b0000000000000000;
	sram_mem[82374] = 16'b0000000000000000;
	sram_mem[82375] = 16'b0000000000000000;
	sram_mem[82376] = 16'b0000000000000000;
	sram_mem[82377] = 16'b0000000000000000;
	sram_mem[82378] = 16'b0000000000000000;
	sram_mem[82379] = 16'b0000000000000000;
	sram_mem[82380] = 16'b0000000000000000;
	sram_mem[82381] = 16'b0000000000000000;
	sram_mem[82382] = 16'b0000000000000000;
	sram_mem[82383] = 16'b0000000000000000;
	sram_mem[82384] = 16'b0000000000000000;
	sram_mem[82385] = 16'b0000000000000000;
	sram_mem[82386] = 16'b0000000000000000;
	sram_mem[82387] = 16'b0000000000000000;
	sram_mem[82388] = 16'b0000000000000000;
	sram_mem[82389] = 16'b0000000000000000;
	sram_mem[82390] = 16'b0000000000000000;
	sram_mem[82391] = 16'b0000000000000000;
	sram_mem[82392] = 16'b0000000000000000;
	sram_mem[82393] = 16'b0000000000000000;
	sram_mem[82394] = 16'b0000000000000000;
	sram_mem[82395] = 16'b0000000000000000;
	sram_mem[82396] = 16'b0000000000000000;
	sram_mem[82397] = 16'b0000000000000000;
	sram_mem[82398] = 16'b0000000000000000;
	sram_mem[82399] = 16'b0000000000000000;
	sram_mem[82400] = 16'b0000000000000000;
	sram_mem[82401] = 16'b0000000000000000;
	sram_mem[82402] = 16'b0000000000000000;
	sram_mem[82403] = 16'b0000000000000000;
	sram_mem[82404] = 16'b0000000000000000;
	sram_mem[82405] = 16'b0000000000000000;
	sram_mem[82406] = 16'b0000000000000000;
	sram_mem[82407] = 16'b0000000000000000;
	sram_mem[82408] = 16'b0000000000000000;
	sram_mem[82409] = 16'b0000000000000000;
	sram_mem[82410] = 16'b0000000000000000;
	sram_mem[82411] = 16'b0000000000000000;
	sram_mem[82412] = 16'b0000000000000000;
	sram_mem[82413] = 16'b0000000000000000;
	sram_mem[82414] = 16'b0000000000000000;
	sram_mem[82415] = 16'b0000000000000000;
	sram_mem[82416] = 16'b0000000000000000;
	sram_mem[82417] = 16'b0000000000000000;
	sram_mem[82418] = 16'b0000000000000000;
	sram_mem[82419] = 16'b0000000000000000;
	sram_mem[82420] = 16'b0000000000000000;
	sram_mem[82421] = 16'b0000000000000000;
	sram_mem[82422] = 16'b0000000000000000;
	sram_mem[82423] = 16'b0000000000000000;
	sram_mem[82424] = 16'b0000000000000000;
	sram_mem[82425] = 16'b0000000000000000;
	sram_mem[82426] = 16'b0000000000000000;
	sram_mem[82427] = 16'b0000000000000000;
	sram_mem[82428] = 16'b0000000000000000;
	sram_mem[82429] = 16'b0000000000000000;
	sram_mem[82430] = 16'b0000000000000000;
	sram_mem[82431] = 16'b0000000000000000;
	sram_mem[82432] = 16'b0000000000000000;
	sram_mem[82433] = 16'b0000000000000000;
	sram_mem[82434] = 16'b0000000000000000;
	sram_mem[82435] = 16'b0000000000000000;
	sram_mem[82436] = 16'b0000000000000000;
	sram_mem[82437] = 16'b0000000000000000;
	sram_mem[82438] = 16'b0000000000000000;
	sram_mem[82439] = 16'b0000000000000000;
	sram_mem[82440] = 16'b0000000000000000;
	sram_mem[82441] = 16'b0000000000000000;
	sram_mem[82442] = 16'b0000000000000000;
	sram_mem[82443] = 16'b0000000000000000;
	sram_mem[82444] = 16'b0000000000000000;
	sram_mem[82445] = 16'b0000000000000000;
	sram_mem[82446] = 16'b0000000000000000;
	sram_mem[82447] = 16'b0000000000000000;
	sram_mem[82448] = 16'b0000000000000000;
	sram_mem[82449] = 16'b0000000000000000;
	sram_mem[82450] = 16'b0000000000000000;
	sram_mem[82451] = 16'b0000000000000000;
	sram_mem[82452] = 16'b0000000000000000;
	sram_mem[82453] = 16'b0000000000000000;
	sram_mem[82454] = 16'b0000000000000000;
	sram_mem[82455] = 16'b0000000000000000;
	sram_mem[82456] = 16'b0000000000000000;
	sram_mem[82457] = 16'b0000000000000000;
	sram_mem[82458] = 16'b0000000000000000;
	sram_mem[82459] = 16'b0000000000000000;
	sram_mem[82460] = 16'b0000000000000000;
	sram_mem[82461] = 16'b0000000000000000;
	sram_mem[82462] = 16'b0000000000000000;
	sram_mem[82463] = 16'b0000000000000000;
	sram_mem[82464] = 16'b0000000000000000;
	sram_mem[82465] = 16'b0000000000000000;
	sram_mem[82466] = 16'b0000000000000000;
	sram_mem[82467] = 16'b0000000000000000;
	sram_mem[82468] = 16'b0000000000000000;
	sram_mem[82469] = 16'b0000000000000000;
	sram_mem[82470] = 16'b0000000000000000;
	sram_mem[82471] = 16'b0000000000000000;
	sram_mem[82472] = 16'b0000000000000000;
	sram_mem[82473] = 16'b0000000000000000;
	sram_mem[82474] = 16'b0000000000000000;
	sram_mem[82475] = 16'b0000000000000000;
	sram_mem[82476] = 16'b0000000000000000;
	sram_mem[82477] = 16'b0000000000000000;
	sram_mem[82478] = 16'b0000000000000000;
	sram_mem[82479] = 16'b0000000000000000;
	sram_mem[82480] = 16'b0000000000000000;
	sram_mem[82481] = 16'b0000000000000000;
	sram_mem[82482] = 16'b0000000000000000;
	sram_mem[82483] = 16'b0000000000000000;
	sram_mem[82484] = 16'b0000000000000000;
	sram_mem[82485] = 16'b0000000000000000;
	sram_mem[82486] = 16'b0000000000000000;
	sram_mem[82487] = 16'b0000000000000000;
	sram_mem[82488] = 16'b0000000000000000;
	sram_mem[82489] = 16'b0000000000000000;
	sram_mem[82490] = 16'b0000000000000000;
	sram_mem[82491] = 16'b0000000000000000;
	sram_mem[82492] = 16'b0000000000000000;
	sram_mem[82493] = 16'b0000000000000000;
	sram_mem[82494] = 16'b0000000000000000;
	sram_mem[82495] = 16'b0000000000000000;
	sram_mem[82496] = 16'b0000000000000000;
	sram_mem[82497] = 16'b0000000000000000;
	sram_mem[82498] = 16'b0000000000000000;
	sram_mem[82499] = 16'b0000000000000000;
	sram_mem[82500] = 16'b0000000000000000;
	sram_mem[82501] = 16'b0000000000000000;
	sram_mem[82502] = 16'b0000000000000000;
	sram_mem[82503] = 16'b0000000000000000;
	sram_mem[82504] = 16'b0000000000000000;
	sram_mem[82505] = 16'b0000000000000000;
	sram_mem[82506] = 16'b0000000000000000;
	sram_mem[82507] = 16'b0000000000000000;
	sram_mem[82508] = 16'b0000000000000000;
	sram_mem[82509] = 16'b0000000000000000;
	sram_mem[82510] = 16'b0000000000000000;
	sram_mem[82511] = 16'b0000000000000000;
	sram_mem[82512] = 16'b0000000000000000;
	sram_mem[82513] = 16'b0000000000000000;
	sram_mem[82514] = 16'b0000000000000000;
	sram_mem[82515] = 16'b0000000000000000;
	sram_mem[82516] = 16'b0000000000000000;
	sram_mem[82517] = 16'b0000000000000000;
	sram_mem[82518] = 16'b0000000000000000;
	sram_mem[82519] = 16'b0000000000000000;
	sram_mem[82520] = 16'b0000000000000000;
	sram_mem[82521] = 16'b0000000000000000;
	sram_mem[82522] = 16'b0000000000000000;
	sram_mem[82523] = 16'b0000000000000000;
	sram_mem[82524] = 16'b0000000000000000;
	sram_mem[82525] = 16'b0000000000000000;
	sram_mem[82526] = 16'b0000000000000000;
	sram_mem[82527] = 16'b0000000000000000;
	sram_mem[82528] = 16'b0000000000000000;
	sram_mem[82529] = 16'b0000000000000000;
	sram_mem[82530] = 16'b0000000000000000;
	sram_mem[82531] = 16'b0000000000000000;
	sram_mem[82532] = 16'b0000000000000000;
	sram_mem[82533] = 16'b0000000000000000;
	sram_mem[82534] = 16'b0000000000000000;
	sram_mem[82535] = 16'b0000000000000000;
	sram_mem[82536] = 16'b0000000000000000;
	sram_mem[82537] = 16'b0000000000000000;
	sram_mem[82538] = 16'b0000000000000000;
	sram_mem[82539] = 16'b0000000000000000;
	sram_mem[82540] = 16'b0000000000000000;
	sram_mem[82541] = 16'b0000000000000000;
	sram_mem[82542] = 16'b0000000000000000;
	sram_mem[82543] = 16'b0000000000000000;
	sram_mem[82544] = 16'b0000000000000000;
	sram_mem[82545] = 16'b0000000000000000;
	sram_mem[82546] = 16'b0000000000000000;
	sram_mem[82547] = 16'b0000000000000000;
	sram_mem[82548] = 16'b0000000000000000;
	sram_mem[82549] = 16'b0000000000000000;
	sram_mem[82550] = 16'b0000000000000000;
	sram_mem[82551] = 16'b0000000000000000;
	sram_mem[82552] = 16'b0000000000000000;
	sram_mem[82553] = 16'b0000000000000000;
	sram_mem[82554] = 16'b0000000000000000;
	sram_mem[82555] = 16'b0000000000000000;
	sram_mem[82556] = 16'b0000000000000000;
	sram_mem[82557] = 16'b0000000000000000;
	sram_mem[82558] = 16'b0000000000000000;
	sram_mem[82559] = 16'b0000000000000000;
	sram_mem[82560] = 16'b0000000000000000;
	sram_mem[82561] = 16'b0000000000000000;
	sram_mem[82562] = 16'b0000000000000000;
	sram_mem[82563] = 16'b0000000000000000;
	sram_mem[82564] = 16'b0000000000000000;
	sram_mem[82565] = 16'b0000000000000000;
	sram_mem[82566] = 16'b0000000000000000;
	sram_mem[82567] = 16'b0000000000000000;
	sram_mem[82568] = 16'b0000000000000000;
	sram_mem[82569] = 16'b0000000000000000;
	sram_mem[82570] = 16'b0000000000000000;
	sram_mem[82571] = 16'b0000000000000000;
	sram_mem[82572] = 16'b0000000000000000;
	sram_mem[82573] = 16'b0000000000000000;
	sram_mem[82574] = 16'b0000000000000000;
	sram_mem[82575] = 16'b0000000000000000;
	sram_mem[82576] = 16'b0000000000000000;
	sram_mem[82577] = 16'b0000000000000000;
	sram_mem[82578] = 16'b0000000000000000;
	sram_mem[82579] = 16'b0000000000000000;
	sram_mem[82580] = 16'b0000000000000000;
	sram_mem[82581] = 16'b0000000000000000;
	sram_mem[82582] = 16'b0000000000000000;
	sram_mem[82583] = 16'b0000000000000000;
	sram_mem[82584] = 16'b0000000000000000;
	sram_mem[82585] = 16'b0000000000000000;
	sram_mem[82586] = 16'b0000000000000000;
	sram_mem[82587] = 16'b0000000000000000;
	sram_mem[82588] = 16'b0000000000000000;
	sram_mem[82589] = 16'b0000000000000000;
	sram_mem[82590] = 16'b0000000000000000;
	sram_mem[82591] = 16'b0000000000000000;
	sram_mem[82592] = 16'b0000000000000000;
	sram_mem[82593] = 16'b0000000000000000;
	sram_mem[82594] = 16'b0000000000000000;
	sram_mem[82595] = 16'b0000000000000000;
	sram_mem[82596] = 16'b0000000000000000;
	sram_mem[82597] = 16'b0000000000000000;
	sram_mem[82598] = 16'b0000000000000000;
	sram_mem[82599] = 16'b0000000000000000;
	sram_mem[82600] = 16'b0000000000000000;
	sram_mem[82601] = 16'b0000000000000000;
	sram_mem[82602] = 16'b0000000000000000;
	sram_mem[82603] = 16'b0000000000000000;
	sram_mem[82604] = 16'b0000000000000000;
	sram_mem[82605] = 16'b0000000000000000;
	sram_mem[82606] = 16'b0000000000000000;
	sram_mem[82607] = 16'b0000000000000000;
	sram_mem[82608] = 16'b0000000000000000;
	sram_mem[82609] = 16'b0000000000000000;
	sram_mem[82610] = 16'b0000000000000000;
	sram_mem[82611] = 16'b0000000000000000;
	sram_mem[82612] = 16'b0000000000000000;
	sram_mem[82613] = 16'b0000000000000000;
	sram_mem[82614] = 16'b0000000000000000;
	sram_mem[82615] = 16'b0000000000000000;
	sram_mem[82616] = 16'b0000000000000000;
	sram_mem[82617] = 16'b0000000000000000;
	sram_mem[82618] = 16'b0000000000000000;
	sram_mem[82619] = 16'b0000000000000000;
	sram_mem[82620] = 16'b0000000000000000;
	sram_mem[82621] = 16'b0000000000000000;
	sram_mem[82622] = 16'b0000000000000000;
	sram_mem[82623] = 16'b0000000000000000;
	sram_mem[82624] = 16'b0000000000000000;
	sram_mem[82625] = 16'b0000000000000000;
	sram_mem[82626] = 16'b0000000000000000;
	sram_mem[82627] = 16'b0000000000000000;
	sram_mem[82628] = 16'b0000000000000000;
	sram_mem[82629] = 16'b0000000000000000;
	sram_mem[82630] = 16'b0000000000000000;
	sram_mem[82631] = 16'b0000000000000000;
	sram_mem[82632] = 16'b0000000000000000;
	sram_mem[82633] = 16'b0000000000000000;
	sram_mem[82634] = 16'b0000000000000000;
	sram_mem[82635] = 16'b0000000000000000;
	sram_mem[82636] = 16'b0000000000000000;
	sram_mem[82637] = 16'b0000000000000000;
	sram_mem[82638] = 16'b0000000000000000;
	sram_mem[82639] = 16'b0000000000000000;
	sram_mem[82640] = 16'b0000000000000000;
	sram_mem[82641] = 16'b0000000000000000;
	sram_mem[82642] = 16'b0000000000000000;
	sram_mem[82643] = 16'b0000000000000000;
	sram_mem[82644] = 16'b0000000000000000;
	sram_mem[82645] = 16'b0000000000000000;
	sram_mem[82646] = 16'b0000000000000000;
	sram_mem[82647] = 16'b0000000000000000;
	sram_mem[82648] = 16'b0000000000000000;
	sram_mem[82649] = 16'b0000000000000000;
	sram_mem[82650] = 16'b0000000000000000;
	sram_mem[82651] = 16'b0000000000000000;
	sram_mem[82652] = 16'b0000000000000000;
	sram_mem[82653] = 16'b0000000000000000;
	sram_mem[82654] = 16'b0000000000000000;
	sram_mem[82655] = 16'b0000000000000000;
	sram_mem[82656] = 16'b0000000000000000;
	sram_mem[82657] = 16'b0000000000000000;
	sram_mem[82658] = 16'b0000000000000000;
	sram_mem[82659] = 16'b0000000000000000;
	sram_mem[82660] = 16'b0000000000000000;
	sram_mem[82661] = 16'b0000000000000000;
	sram_mem[82662] = 16'b0000000000000000;
	sram_mem[82663] = 16'b0000000000000000;
	sram_mem[82664] = 16'b0000000000000000;
	sram_mem[82665] = 16'b0000000000000000;
	sram_mem[82666] = 16'b0000000000000000;
	sram_mem[82667] = 16'b0000000000000000;
	sram_mem[82668] = 16'b0000000000000000;
	sram_mem[82669] = 16'b0000000000000000;
	sram_mem[82670] = 16'b0000000000000000;
	sram_mem[82671] = 16'b0000000000000000;
	sram_mem[82672] = 16'b0000000000000000;
	sram_mem[82673] = 16'b0000000000000000;
	sram_mem[82674] = 16'b0000000000000000;
	sram_mem[82675] = 16'b0000000000000000;
	sram_mem[82676] = 16'b0000000000000000;
	sram_mem[82677] = 16'b0000000000000000;
	sram_mem[82678] = 16'b0000000000000000;
	sram_mem[82679] = 16'b0000000000000000;
	sram_mem[82680] = 16'b0000000000000000;
	sram_mem[82681] = 16'b0000000000000000;
	sram_mem[82682] = 16'b0000000000000000;
	sram_mem[82683] = 16'b0000000000000000;
	sram_mem[82684] = 16'b0000000000000000;
	sram_mem[82685] = 16'b0000000000000000;
	sram_mem[82686] = 16'b0000000000000000;
	sram_mem[82687] = 16'b0000000000000000;
	sram_mem[82688] = 16'b0000000000000000;
	sram_mem[82689] = 16'b0000000000000000;
	sram_mem[82690] = 16'b0000000000000000;
	sram_mem[82691] = 16'b0000000000000000;
	sram_mem[82692] = 16'b0000000000000000;
	sram_mem[82693] = 16'b0000000000000000;
	sram_mem[82694] = 16'b0000000000000000;
	sram_mem[82695] = 16'b0000000000000000;
	sram_mem[82696] = 16'b0000000000000000;
	sram_mem[82697] = 16'b0000000000000000;
	sram_mem[82698] = 16'b0000000000000000;
	sram_mem[82699] = 16'b0000000000000000;
	sram_mem[82700] = 16'b0000000000000000;
	sram_mem[82701] = 16'b0000000000000000;
	sram_mem[82702] = 16'b0000000000000000;
	sram_mem[82703] = 16'b0000000000000000;
	sram_mem[82704] = 16'b0000000000000000;
	sram_mem[82705] = 16'b0000000000000000;
	sram_mem[82706] = 16'b0000000000000000;
	sram_mem[82707] = 16'b0000000000000000;
	sram_mem[82708] = 16'b0000000000000000;
	sram_mem[82709] = 16'b0000000000000000;
	sram_mem[82710] = 16'b0000000000000000;
	sram_mem[82711] = 16'b0000000000000000;
	sram_mem[82712] = 16'b0000000000000000;
	sram_mem[82713] = 16'b0000000000000000;
	sram_mem[82714] = 16'b0000000000000000;
	sram_mem[82715] = 16'b0000000000000000;
	sram_mem[82716] = 16'b0000000000000000;
	sram_mem[82717] = 16'b0000000000000000;
	sram_mem[82718] = 16'b0000000000000000;
	sram_mem[82719] = 16'b0000000000000000;
	sram_mem[82720] = 16'b0000000000000000;
	sram_mem[82721] = 16'b0000000000000000;
	sram_mem[82722] = 16'b0000000000000000;
	sram_mem[82723] = 16'b0000000000000000;
	sram_mem[82724] = 16'b0000000000000000;
	sram_mem[82725] = 16'b0000000000000000;
	sram_mem[82726] = 16'b0000000000000000;
	sram_mem[82727] = 16'b0000000000000000;
	sram_mem[82728] = 16'b0000000000000000;
	sram_mem[82729] = 16'b0000000000000000;
	sram_mem[82730] = 16'b0000000000000000;
	sram_mem[82731] = 16'b0000000000000000;
	sram_mem[82732] = 16'b0000000000000000;
	sram_mem[82733] = 16'b0000000000000000;
	sram_mem[82734] = 16'b0000000000000000;
	sram_mem[82735] = 16'b0000000000000000;
	sram_mem[82736] = 16'b0000000000000000;
	sram_mem[82737] = 16'b0000000000000000;
	sram_mem[82738] = 16'b0000000000000000;
	sram_mem[82739] = 16'b0000000000000000;
	sram_mem[82740] = 16'b0000000000000000;
	sram_mem[82741] = 16'b0000000000000000;
	sram_mem[82742] = 16'b0000000000000000;
	sram_mem[82743] = 16'b0000000000000000;
	sram_mem[82744] = 16'b0000000000000000;
	sram_mem[82745] = 16'b0000000000000000;
	sram_mem[82746] = 16'b0000000000000000;
	sram_mem[82747] = 16'b0000000000000000;
	sram_mem[82748] = 16'b0000000000000000;
	sram_mem[82749] = 16'b0000000000000000;
	sram_mem[82750] = 16'b0000000000000000;
	sram_mem[82751] = 16'b0000000000000000;
	sram_mem[82752] = 16'b0000000000000000;
	sram_mem[82753] = 16'b0000000000000000;
	sram_mem[82754] = 16'b0000000000000000;
	sram_mem[82755] = 16'b0000000000000000;
	sram_mem[82756] = 16'b0000000000000000;
	sram_mem[82757] = 16'b0000000000000000;
	sram_mem[82758] = 16'b0000000000000000;
	sram_mem[82759] = 16'b0000000000000000;
	sram_mem[82760] = 16'b0000000000000000;
	sram_mem[82761] = 16'b0000000000000000;
	sram_mem[82762] = 16'b0000000000000000;
	sram_mem[82763] = 16'b0000000000000000;
	sram_mem[82764] = 16'b0000000000000000;
	sram_mem[82765] = 16'b0000000000000000;
	sram_mem[82766] = 16'b0000000000000000;
	sram_mem[82767] = 16'b0000000000000000;
	sram_mem[82768] = 16'b0000000000000000;
	sram_mem[82769] = 16'b0000000000000000;
	sram_mem[82770] = 16'b0000000000000000;
	sram_mem[82771] = 16'b0000000000000000;
	sram_mem[82772] = 16'b0000000000000000;
	sram_mem[82773] = 16'b0000000000000000;
	sram_mem[82774] = 16'b0000000000000000;
	sram_mem[82775] = 16'b0000000000000000;
	sram_mem[82776] = 16'b0000000000000000;
	sram_mem[82777] = 16'b0000000000000000;
	sram_mem[82778] = 16'b0000000000000000;
	sram_mem[82779] = 16'b0000000000000000;
	sram_mem[82780] = 16'b0000000000000000;
	sram_mem[82781] = 16'b0000000000000000;
	sram_mem[82782] = 16'b0000000000000000;
	sram_mem[82783] = 16'b0000000000000000;
	sram_mem[82784] = 16'b0000000000000000;
	sram_mem[82785] = 16'b0000000000000000;
	sram_mem[82786] = 16'b0000000000000000;
	sram_mem[82787] = 16'b0000000000000000;
	sram_mem[82788] = 16'b0000000000000000;
	sram_mem[82789] = 16'b0000000000000000;
	sram_mem[82790] = 16'b0000000000000000;
	sram_mem[82791] = 16'b0000000000000000;
	sram_mem[82792] = 16'b0000000000000000;
	sram_mem[82793] = 16'b0000000000000000;
	sram_mem[82794] = 16'b0000000000000000;
	sram_mem[82795] = 16'b0000000000000000;
	sram_mem[82796] = 16'b0000000000000000;
	sram_mem[82797] = 16'b0000000000000000;
	sram_mem[82798] = 16'b0000000000000000;
	sram_mem[82799] = 16'b0000000000000000;
	sram_mem[82800] = 16'b0000000000000000;
	sram_mem[82801] = 16'b0000000000000000;
	sram_mem[82802] = 16'b0000000000000000;
	sram_mem[82803] = 16'b0000000000000000;
	sram_mem[82804] = 16'b0000000000000000;
	sram_mem[82805] = 16'b0000000000000000;
	sram_mem[82806] = 16'b0000000000000000;
	sram_mem[82807] = 16'b0000000000000000;
	sram_mem[82808] = 16'b0000000000000000;
	sram_mem[82809] = 16'b0000000000000000;
	sram_mem[82810] = 16'b0000000000000000;
	sram_mem[82811] = 16'b0000000000000000;
	sram_mem[82812] = 16'b0000000000000000;
	sram_mem[82813] = 16'b0000000000000000;
	sram_mem[82814] = 16'b0000000000000000;
	sram_mem[82815] = 16'b0000000000000000;
	sram_mem[82816] = 16'b0000000000000000;
	sram_mem[82817] = 16'b0000000000000000;
	sram_mem[82818] = 16'b0000000000000000;
	sram_mem[82819] = 16'b0000000000000000;
	sram_mem[82820] = 16'b0000000000000000;
	sram_mem[82821] = 16'b0000000000000000;
	sram_mem[82822] = 16'b0000000000000000;
	sram_mem[82823] = 16'b0000000000000000;
	sram_mem[82824] = 16'b0000000000000000;
	sram_mem[82825] = 16'b0000000000000000;
	sram_mem[82826] = 16'b0000000000000000;
	sram_mem[82827] = 16'b0000000000000000;
	sram_mem[82828] = 16'b0000000000000000;
	sram_mem[82829] = 16'b0000000000000000;
	sram_mem[82830] = 16'b0000000000000000;
	sram_mem[82831] = 16'b0000000000000000;
	sram_mem[82832] = 16'b0000000000000000;
	sram_mem[82833] = 16'b0000000000000000;
	sram_mem[82834] = 16'b0000000000000000;
	sram_mem[82835] = 16'b0000000000000000;
	sram_mem[82836] = 16'b0000000000000000;
	sram_mem[82837] = 16'b0000000000000000;
	sram_mem[82838] = 16'b0000000000000000;
	sram_mem[82839] = 16'b0000000000000000;
	sram_mem[82840] = 16'b0000000000000000;
	sram_mem[82841] = 16'b0000000000000000;
	sram_mem[82842] = 16'b0000000000000000;
	sram_mem[82843] = 16'b0000000000000000;
	sram_mem[82844] = 16'b0000000000000000;
	sram_mem[82845] = 16'b0000000000000000;
	sram_mem[82846] = 16'b0000000000000000;
	sram_mem[82847] = 16'b0000000000000000;
	sram_mem[82848] = 16'b0000000000000000;
	sram_mem[82849] = 16'b0000000000000000;
	sram_mem[82850] = 16'b0000000000000000;
	sram_mem[82851] = 16'b0000000000000000;
	sram_mem[82852] = 16'b0000000000000000;
	sram_mem[82853] = 16'b0000000000000000;
	sram_mem[82854] = 16'b0000000000000000;
	sram_mem[82855] = 16'b0000000000000000;
	sram_mem[82856] = 16'b0000000000000000;
	sram_mem[82857] = 16'b0000000000000000;
	sram_mem[82858] = 16'b0000000000000000;
	sram_mem[82859] = 16'b0000000000000000;
	sram_mem[82860] = 16'b0000000000000000;
	sram_mem[82861] = 16'b0000000000000000;
	sram_mem[82862] = 16'b0000000000000000;
	sram_mem[82863] = 16'b0000000000000000;
	sram_mem[82864] = 16'b0000000000000000;
	sram_mem[82865] = 16'b0000000000000000;
	sram_mem[82866] = 16'b0000000000000000;
	sram_mem[82867] = 16'b0000000000000000;
	sram_mem[82868] = 16'b0000000000000000;
	sram_mem[82869] = 16'b0000000000000000;
	sram_mem[82870] = 16'b0000000000000000;
	sram_mem[82871] = 16'b0000000000000000;
	sram_mem[82872] = 16'b0000000000000000;
	sram_mem[82873] = 16'b0000000000000000;
	sram_mem[82874] = 16'b0000000000000000;
	sram_mem[82875] = 16'b0000000000000000;
	sram_mem[82876] = 16'b0000000000000000;
	sram_mem[82877] = 16'b0000000000000000;
	sram_mem[82878] = 16'b0000000000000000;
	sram_mem[82879] = 16'b0000000000000000;
	sram_mem[82880] = 16'b0000000000000000;
	sram_mem[82881] = 16'b0000000000000000;
	sram_mem[82882] = 16'b0000000000000000;
	sram_mem[82883] = 16'b0000000000000000;
	sram_mem[82884] = 16'b0000000000000000;
	sram_mem[82885] = 16'b0000000000000000;
	sram_mem[82886] = 16'b0000000000000000;
	sram_mem[82887] = 16'b0000000000000000;
	sram_mem[82888] = 16'b0000000000000000;
	sram_mem[82889] = 16'b0000000000000000;
	sram_mem[82890] = 16'b0000000000000000;
	sram_mem[82891] = 16'b0000000000000000;
	sram_mem[82892] = 16'b0000000000000000;
	sram_mem[82893] = 16'b0000000000000000;
	sram_mem[82894] = 16'b0000000000000000;
	sram_mem[82895] = 16'b0000000000000000;
	sram_mem[82896] = 16'b0000000000000000;
	sram_mem[82897] = 16'b0000000000000000;
	sram_mem[82898] = 16'b0000000000000000;
	sram_mem[82899] = 16'b0000000000000000;
	sram_mem[82900] = 16'b0000000000000000;
	sram_mem[82901] = 16'b0000000000000000;
	sram_mem[82902] = 16'b0000000000000000;
	sram_mem[82903] = 16'b0000000000000000;
	sram_mem[82904] = 16'b0000000000000000;
	sram_mem[82905] = 16'b0000000000000000;
	sram_mem[82906] = 16'b0000000000000000;
	sram_mem[82907] = 16'b0000000000000000;
	sram_mem[82908] = 16'b0000000000000000;
	sram_mem[82909] = 16'b0000000000000000;
	sram_mem[82910] = 16'b0000000000000000;
	sram_mem[82911] = 16'b0000000000000000;
	sram_mem[82912] = 16'b0000000000000000;
	sram_mem[82913] = 16'b0000000000000000;
	sram_mem[82914] = 16'b0000000000000000;
	sram_mem[82915] = 16'b0000000000000000;
	sram_mem[82916] = 16'b0000000000000000;
	sram_mem[82917] = 16'b0000000000000000;
	sram_mem[82918] = 16'b0000000000000000;
	sram_mem[82919] = 16'b0000000000000000;
	sram_mem[82920] = 16'b0000000000000000;
	sram_mem[82921] = 16'b0000000000000000;
	sram_mem[82922] = 16'b0000000000000000;
	sram_mem[82923] = 16'b0000000000000000;
	sram_mem[82924] = 16'b0000000000000000;
	sram_mem[82925] = 16'b0000000000000000;
	sram_mem[82926] = 16'b0000000000000000;
	sram_mem[82927] = 16'b0000000000000000;
	sram_mem[82928] = 16'b0000000000000000;
	sram_mem[82929] = 16'b0000000000000000;
	sram_mem[82930] = 16'b0000000000000000;
	sram_mem[82931] = 16'b0000000000000000;
	sram_mem[82932] = 16'b0000000000000000;
	sram_mem[82933] = 16'b0000000000000000;
	sram_mem[82934] = 16'b0000000000000000;
	sram_mem[82935] = 16'b0000000000000000;
	sram_mem[82936] = 16'b0000000000000000;
	sram_mem[82937] = 16'b0000000000000000;
	sram_mem[82938] = 16'b0000000000000000;
	sram_mem[82939] = 16'b0000000000000000;
	sram_mem[82940] = 16'b0000000000000000;
	sram_mem[82941] = 16'b0000000000000000;
	sram_mem[82942] = 16'b0000000000000000;
	sram_mem[82943] = 16'b0000000000000000;
	sram_mem[82944] = 16'b0000000000000000;
	sram_mem[82945] = 16'b0000000000000000;
	sram_mem[82946] = 16'b0000000000000000;
	sram_mem[82947] = 16'b0000000000000000;
	sram_mem[82948] = 16'b0000000000000000;
	sram_mem[82949] = 16'b0000000000000000;
	sram_mem[82950] = 16'b0000000000000000;
	sram_mem[82951] = 16'b0000000000000000;
	sram_mem[82952] = 16'b0000000000000000;
	sram_mem[82953] = 16'b0000000000000000;
	sram_mem[82954] = 16'b0000000000000000;
	sram_mem[82955] = 16'b0000000000000000;
	sram_mem[82956] = 16'b0000000000000000;
	sram_mem[82957] = 16'b0000000000000000;
	sram_mem[82958] = 16'b0000000000000000;
	sram_mem[82959] = 16'b0000000000000000;
	sram_mem[82960] = 16'b0000000000000000;
	sram_mem[82961] = 16'b0000000000000000;
	sram_mem[82962] = 16'b0000000000000000;
	sram_mem[82963] = 16'b0000000000000000;
	sram_mem[82964] = 16'b0000000000000000;
	sram_mem[82965] = 16'b0000000000000000;
	sram_mem[82966] = 16'b0000000000000000;
	sram_mem[82967] = 16'b0000000000000000;
	sram_mem[82968] = 16'b0000000000000000;
	sram_mem[82969] = 16'b0000000000000000;
	sram_mem[82970] = 16'b0000000000000000;
	sram_mem[82971] = 16'b0000000000000000;
	sram_mem[82972] = 16'b0000000000000000;
	sram_mem[82973] = 16'b0000000000000000;
	sram_mem[82974] = 16'b0000000000000000;
	sram_mem[82975] = 16'b0000000000000000;
	sram_mem[82976] = 16'b0000000000000000;
	sram_mem[82977] = 16'b0000000000000000;
	sram_mem[82978] = 16'b0000000000000000;
	sram_mem[82979] = 16'b0000000000000000;
	sram_mem[82980] = 16'b0000000000000000;
	sram_mem[82981] = 16'b0000000000000000;
	sram_mem[82982] = 16'b0000000000000000;
	sram_mem[82983] = 16'b0000000000000000;
	sram_mem[82984] = 16'b0000000000000000;
	sram_mem[82985] = 16'b0000000000000000;
	sram_mem[82986] = 16'b0000000000000000;
	sram_mem[82987] = 16'b0000000000000000;
	sram_mem[82988] = 16'b0000000000000000;
	sram_mem[82989] = 16'b0000000000000000;
	sram_mem[82990] = 16'b0000000000000000;
	sram_mem[82991] = 16'b0000000000000000;
	sram_mem[82992] = 16'b0000000000000000;
	sram_mem[82993] = 16'b0000000000000000;
	sram_mem[82994] = 16'b0000000000000000;
	sram_mem[82995] = 16'b0000000000000000;
	sram_mem[82996] = 16'b0000000000000000;
	sram_mem[82997] = 16'b0000000000000000;
	sram_mem[82998] = 16'b0000000000000000;
	sram_mem[82999] = 16'b0000000000000000;
	sram_mem[83000] = 16'b0000000000000000;
	sram_mem[83001] = 16'b0000000000000000;
	sram_mem[83002] = 16'b0000000000000000;
	sram_mem[83003] = 16'b0000000000000000;
	sram_mem[83004] = 16'b0000000000000000;
	sram_mem[83005] = 16'b0000000000000000;
	sram_mem[83006] = 16'b0000000000000000;
	sram_mem[83007] = 16'b0000000000000000;
	sram_mem[83008] = 16'b0000000000000000;
	sram_mem[83009] = 16'b0000000000000000;
	sram_mem[83010] = 16'b0000000000000000;
	sram_mem[83011] = 16'b0000000000000000;
	sram_mem[83012] = 16'b0000000000000000;
	sram_mem[83013] = 16'b0000000000000000;
	sram_mem[83014] = 16'b0000000000000000;
	sram_mem[83015] = 16'b0000000000000000;
	sram_mem[83016] = 16'b0000000000000000;
	sram_mem[83017] = 16'b0000000000000000;
	sram_mem[83018] = 16'b0000000000000000;
	sram_mem[83019] = 16'b0000000000000000;
	sram_mem[83020] = 16'b0000000000000000;
	sram_mem[83021] = 16'b0000000000000000;
	sram_mem[83022] = 16'b0000000000000000;
	sram_mem[83023] = 16'b0000000000000000;
	sram_mem[83024] = 16'b0000000000000000;
	sram_mem[83025] = 16'b0000000000000000;
	sram_mem[83026] = 16'b0000000000000000;
	sram_mem[83027] = 16'b0000000000000000;
	sram_mem[83028] = 16'b0000000000000000;
	sram_mem[83029] = 16'b0000000000000000;
	sram_mem[83030] = 16'b0000000000000000;
	sram_mem[83031] = 16'b0000000000000000;
	sram_mem[83032] = 16'b0000000000000000;
	sram_mem[83033] = 16'b0000000000000000;
	sram_mem[83034] = 16'b0000000000000000;
	sram_mem[83035] = 16'b0000000000000000;
	sram_mem[83036] = 16'b0000000000000000;
	sram_mem[83037] = 16'b0000000000000000;
	sram_mem[83038] = 16'b0000000000000000;
	sram_mem[83039] = 16'b0000000000000000;
	sram_mem[83040] = 16'b0000000000000000;
	sram_mem[83041] = 16'b0000000000000000;
	sram_mem[83042] = 16'b0000000000000000;
	sram_mem[83043] = 16'b0000000000000000;
	sram_mem[83044] = 16'b0000000000000000;
	sram_mem[83045] = 16'b0000000000000000;
	sram_mem[83046] = 16'b0000000000000000;
	sram_mem[83047] = 16'b0000000000000000;
	sram_mem[83048] = 16'b0000000000000000;
	sram_mem[83049] = 16'b0000000000000000;
	sram_mem[83050] = 16'b0000000000000000;
	sram_mem[83051] = 16'b0000000000000000;
	sram_mem[83052] = 16'b0000000000000000;
	sram_mem[83053] = 16'b0000000000000000;
	sram_mem[83054] = 16'b0000000000000000;
	sram_mem[83055] = 16'b0000000000000000;
	sram_mem[83056] = 16'b0000000000000000;
	sram_mem[83057] = 16'b0000000000000000;
	sram_mem[83058] = 16'b0000000000000000;
	sram_mem[83059] = 16'b0000000000000000;
	sram_mem[83060] = 16'b0000000000000000;
	sram_mem[83061] = 16'b0000000000000000;
	sram_mem[83062] = 16'b0000000000000000;
	sram_mem[83063] = 16'b0000000000000000;
	sram_mem[83064] = 16'b0000000000000000;
	sram_mem[83065] = 16'b0000000000000000;
	sram_mem[83066] = 16'b0000000000000000;
	sram_mem[83067] = 16'b0000000000000000;
	sram_mem[83068] = 16'b0000000000000000;
	sram_mem[83069] = 16'b0000000000000000;
	sram_mem[83070] = 16'b0000000000000000;
	sram_mem[83071] = 16'b0000000000000000;
	sram_mem[83072] = 16'b0000000000000000;
	sram_mem[83073] = 16'b0000000000000000;
	sram_mem[83074] = 16'b0000000000000000;
	sram_mem[83075] = 16'b0000000000000000;
	sram_mem[83076] = 16'b0000000000000000;
	sram_mem[83077] = 16'b0000000000000000;
	sram_mem[83078] = 16'b0000000000000000;
	sram_mem[83079] = 16'b0000000000000000;
	sram_mem[83080] = 16'b0000000000000000;
	sram_mem[83081] = 16'b0000000000000000;
	sram_mem[83082] = 16'b0000000000000000;
	sram_mem[83083] = 16'b0000000000000000;
	sram_mem[83084] = 16'b0000000000000000;
	sram_mem[83085] = 16'b0000000000000000;
	sram_mem[83086] = 16'b0000000000000000;
	sram_mem[83087] = 16'b0000000000000000;
	sram_mem[83088] = 16'b0000000000000000;
	sram_mem[83089] = 16'b0000000000000000;
	sram_mem[83090] = 16'b0000000000000000;
	sram_mem[83091] = 16'b0000000000000000;
	sram_mem[83092] = 16'b0000000000000000;
	sram_mem[83093] = 16'b0000000000000000;
	sram_mem[83094] = 16'b0000000000000000;
	sram_mem[83095] = 16'b0000000000000000;
	sram_mem[83096] = 16'b0000000000000000;
	sram_mem[83097] = 16'b0000000000000000;
	sram_mem[83098] = 16'b0000000000000000;
	sram_mem[83099] = 16'b0000000000000000;
	sram_mem[83100] = 16'b0000000000000000;
	sram_mem[83101] = 16'b0000000000000000;
	sram_mem[83102] = 16'b0000000000000000;
	sram_mem[83103] = 16'b0000000000000000;
	sram_mem[83104] = 16'b0000000000000000;
	sram_mem[83105] = 16'b0000000000000000;
	sram_mem[83106] = 16'b0000000000000000;
	sram_mem[83107] = 16'b0000000000000000;
	sram_mem[83108] = 16'b0000000000000000;
	sram_mem[83109] = 16'b0000000000000000;
	sram_mem[83110] = 16'b0000000000000000;
	sram_mem[83111] = 16'b0000000000000000;
	sram_mem[83112] = 16'b0000000000000000;
	sram_mem[83113] = 16'b0000000000000000;
	sram_mem[83114] = 16'b0000000000000000;
	sram_mem[83115] = 16'b0000000000000000;
	sram_mem[83116] = 16'b0000000000000000;
	sram_mem[83117] = 16'b0000000000000000;
	sram_mem[83118] = 16'b0000000000000000;
	sram_mem[83119] = 16'b0000000000000000;
	sram_mem[83120] = 16'b0000000000000000;
	sram_mem[83121] = 16'b0000000000000000;
	sram_mem[83122] = 16'b0000000000000000;
	sram_mem[83123] = 16'b0000000000000000;
	sram_mem[83124] = 16'b0000000000000000;
	sram_mem[83125] = 16'b0000000000000000;
	sram_mem[83126] = 16'b0000000000000000;
	sram_mem[83127] = 16'b0000000000000000;
	sram_mem[83128] = 16'b0000000000000000;
	sram_mem[83129] = 16'b0000000000000000;
	sram_mem[83130] = 16'b0000000000000000;
	sram_mem[83131] = 16'b0000000000000000;
	sram_mem[83132] = 16'b0000000000000000;
	sram_mem[83133] = 16'b0000000000000000;
	sram_mem[83134] = 16'b0000000000000000;
	sram_mem[83135] = 16'b0000000000000000;
	sram_mem[83136] = 16'b0000000000000000;
	sram_mem[83137] = 16'b0000000000000000;
	sram_mem[83138] = 16'b0000000000000000;
	sram_mem[83139] = 16'b0000000000000000;
	sram_mem[83140] = 16'b0000000000000000;
	sram_mem[83141] = 16'b0000000000000000;
	sram_mem[83142] = 16'b0000000000000000;
	sram_mem[83143] = 16'b0000000000000000;
	sram_mem[83144] = 16'b0000000000000000;
	sram_mem[83145] = 16'b0000000000000000;
	sram_mem[83146] = 16'b0000000000000000;
	sram_mem[83147] = 16'b0000000000000000;
	sram_mem[83148] = 16'b0000000000000000;
	sram_mem[83149] = 16'b0000000000000000;
	sram_mem[83150] = 16'b0000000000000000;
	sram_mem[83151] = 16'b0000000000000000;
	sram_mem[83152] = 16'b0000000000000000;
	sram_mem[83153] = 16'b0000000000000000;
	sram_mem[83154] = 16'b0000000000000000;
	sram_mem[83155] = 16'b0000000000000000;
	sram_mem[83156] = 16'b0000000000000000;
	sram_mem[83157] = 16'b0000000000000000;
	sram_mem[83158] = 16'b0000000000000000;
	sram_mem[83159] = 16'b0000000000000000;
	sram_mem[83160] = 16'b0000000000000000;
	sram_mem[83161] = 16'b0000000000000000;
	sram_mem[83162] = 16'b0000000000000000;
	sram_mem[83163] = 16'b0000000000000000;
	sram_mem[83164] = 16'b0000000000000000;
	sram_mem[83165] = 16'b0000000000000000;
	sram_mem[83166] = 16'b0000000000000000;
	sram_mem[83167] = 16'b0000000000000000;
	sram_mem[83168] = 16'b0000000000000000;
	sram_mem[83169] = 16'b0000000000000000;
	sram_mem[83170] = 16'b0000000000000000;
	sram_mem[83171] = 16'b0000000000000000;
	sram_mem[83172] = 16'b0000000000000000;
	sram_mem[83173] = 16'b0000000000000000;
	sram_mem[83174] = 16'b0000000000000000;
	sram_mem[83175] = 16'b0000000000000000;
	sram_mem[83176] = 16'b0000000000000000;
	sram_mem[83177] = 16'b0000000000000000;
	sram_mem[83178] = 16'b0000000000000000;
	sram_mem[83179] = 16'b0000000000000000;
	sram_mem[83180] = 16'b0000000000000000;
	sram_mem[83181] = 16'b0000000000000000;
	sram_mem[83182] = 16'b0000000000000000;
	sram_mem[83183] = 16'b0000000000000000;
	sram_mem[83184] = 16'b0000000000000000;
	sram_mem[83185] = 16'b0000000000000000;
	sram_mem[83186] = 16'b0000000000000000;
	sram_mem[83187] = 16'b0000000000000000;
	sram_mem[83188] = 16'b0000000000000000;
	sram_mem[83189] = 16'b0000000000000000;
	sram_mem[83190] = 16'b0000000000000000;
	sram_mem[83191] = 16'b0000000000000000;
	sram_mem[83192] = 16'b0000000000000000;
	sram_mem[83193] = 16'b0000000000000000;
	sram_mem[83194] = 16'b0000000000000000;
	sram_mem[83195] = 16'b0000000000000000;
	sram_mem[83196] = 16'b0000000000000000;
	sram_mem[83197] = 16'b0000000000000000;
	sram_mem[83198] = 16'b0000000000000000;
	sram_mem[83199] = 16'b0000000000000000;
	sram_mem[83200] = 16'b0000000000000000;
	sram_mem[83201] = 16'b0000000000000000;
	sram_mem[83202] = 16'b0000000000000000;
	sram_mem[83203] = 16'b0000000000000000;
	sram_mem[83204] = 16'b0000000000000000;
	sram_mem[83205] = 16'b0000000000000000;
	sram_mem[83206] = 16'b0000000000000000;
	sram_mem[83207] = 16'b0000000000000000;
	sram_mem[83208] = 16'b0000000000000000;
	sram_mem[83209] = 16'b0000000000000000;
	sram_mem[83210] = 16'b0000000000000000;
	sram_mem[83211] = 16'b0000000000000000;
	sram_mem[83212] = 16'b0000000000000000;
	sram_mem[83213] = 16'b0000000000000000;
	sram_mem[83214] = 16'b0000000000000000;
	sram_mem[83215] = 16'b0000000000000000;
	sram_mem[83216] = 16'b0000000000000000;
	sram_mem[83217] = 16'b0000000000000000;
	sram_mem[83218] = 16'b0000000000000000;
	sram_mem[83219] = 16'b0000000000000000;
	sram_mem[83220] = 16'b0000000000000000;
	sram_mem[83221] = 16'b0000000000000000;
	sram_mem[83222] = 16'b0000000000000000;
	sram_mem[83223] = 16'b0000000000000000;
	sram_mem[83224] = 16'b0000000000000000;
	sram_mem[83225] = 16'b0000000000000000;
	sram_mem[83226] = 16'b0000000000000000;
	sram_mem[83227] = 16'b0000000000000000;
	sram_mem[83228] = 16'b0000000000000000;
	sram_mem[83229] = 16'b0000000000000000;
	sram_mem[83230] = 16'b0000000000000000;
	sram_mem[83231] = 16'b0000000000000000;
	sram_mem[83232] = 16'b0000000000000000;
	sram_mem[83233] = 16'b0000000000000000;
	sram_mem[83234] = 16'b0000000000000000;
	sram_mem[83235] = 16'b0000000000000000;
	sram_mem[83236] = 16'b0000000000000000;
	sram_mem[83237] = 16'b0000000000000000;
	sram_mem[83238] = 16'b0000000000000000;
	sram_mem[83239] = 16'b0000000000000000;
	sram_mem[83240] = 16'b0000000000000000;
	sram_mem[83241] = 16'b0000000000000000;
	sram_mem[83242] = 16'b0000000000000000;
	sram_mem[83243] = 16'b0000000000000000;
	sram_mem[83244] = 16'b0000000000000000;
	sram_mem[83245] = 16'b0000000000000000;
	sram_mem[83246] = 16'b0000000000000000;
	sram_mem[83247] = 16'b0000000000000000;
	sram_mem[83248] = 16'b0000000000000000;
	sram_mem[83249] = 16'b0000000000000000;
	sram_mem[83250] = 16'b0000000000000000;
	sram_mem[83251] = 16'b0000000000000000;
	sram_mem[83252] = 16'b0000000000000000;
	sram_mem[83253] = 16'b0000000000000000;
	sram_mem[83254] = 16'b0000000000000000;
	sram_mem[83255] = 16'b0000000000000000;
	sram_mem[83256] = 16'b0000000000000000;
	sram_mem[83257] = 16'b0000000000000000;
	sram_mem[83258] = 16'b0000000000000000;
	sram_mem[83259] = 16'b0000000000000000;
	sram_mem[83260] = 16'b0000000000000000;
	sram_mem[83261] = 16'b0000000000000000;
	sram_mem[83262] = 16'b0000000000000000;
	sram_mem[83263] = 16'b0000000000000000;
	sram_mem[83264] = 16'b0000000000000000;
	sram_mem[83265] = 16'b0000000000000000;
	sram_mem[83266] = 16'b0000000000000000;
	sram_mem[83267] = 16'b0000000000000000;
	sram_mem[83268] = 16'b0000000000000000;
	sram_mem[83269] = 16'b0000000000000000;
	sram_mem[83270] = 16'b0000000000000000;
	sram_mem[83271] = 16'b0000000000000000;
	sram_mem[83272] = 16'b0000000000000000;
	sram_mem[83273] = 16'b0000000000000000;
	sram_mem[83274] = 16'b0000000000000000;
	sram_mem[83275] = 16'b0000000000000000;
	sram_mem[83276] = 16'b0000000000000000;
	sram_mem[83277] = 16'b0000000000000000;
	sram_mem[83278] = 16'b0000000000000000;
	sram_mem[83279] = 16'b0000000000000000;
	sram_mem[83280] = 16'b0000000000000000;
	sram_mem[83281] = 16'b0000000000000000;
	sram_mem[83282] = 16'b0000000000000000;
	sram_mem[83283] = 16'b0000000000000000;
	sram_mem[83284] = 16'b0000000000000000;
	sram_mem[83285] = 16'b0000000000000000;
	sram_mem[83286] = 16'b0000000000000000;
	sram_mem[83287] = 16'b0000000000000000;
	sram_mem[83288] = 16'b0000000000000000;
	sram_mem[83289] = 16'b0000000000000000;
	sram_mem[83290] = 16'b0000000000000000;
	sram_mem[83291] = 16'b0000000000000000;
	sram_mem[83292] = 16'b0000000000000000;
	sram_mem[83293] = 16'b0000000000000000;
	sram_mem[83294] = 16'b0000000000000000;
	sram_mem[83295] = 16'b0000000000000000;
	sram_mem[83296] = 16'b0000000000000000;
	sram_mem[83297] = 16'b0000000000000000;
	sram_mem[83298] = 16'b0000000000000000;
	sram_mem[83299] = 16'b0000000000000000;
	sram_mem[83300] = 16'b0000000000000000;
	sram_mem[83301] = 16'b0000000000000000;
	sram_mem[83302] = 16'b0000000000000000;
	sram_mem[83303] = 16'b0000000000000000;
	sram_mem[83304] = 16'b0000000000000000;
	sram_mem[83305] = 16'b0000000000000000;
	sram_mem[83306] = 16'b0000000000000000;
	sram_mem[83307] = 16'b0000000000000000;
	sram_mem[83308] = 16'b0000000000000000;
	sram_mem[83309] = 16'b0000000000000000;
	sram_mem[83310] = 16'b0000000000000000;
	sram_mem[83311] = 16'b0000000000000000;
	sram_mem[83312] = 16'b0000000000000000;
	sram_mem[83313] = 16'b0000000000000000;
	sram_mem[83314] = 16'b0000000000000000;
	sram_mem[83315] = 16'b0000000000000000;
	sram_mem[83316] = 16'b0000000000000000;
	sram_mem[83317] = 16'b0000000000000000;
	sram_mem[83318] = 16'b0000000000000000;
	sram_mem[83319] = 16'b0000000000000000;
	sram_mem[83320] = 16'b0000000000000000;
	sram_mem[83321] = 16'b0000000000000000;
	sram_mem[83322] = 16'b0000000000000000;
	sram_mem[83323] = 16'b0000000000000000;
	sram_mem[83324] = 16'b0000000000000000;
	sram_mem[83325] = 16'b0000000000000000;
	sram_mem[83326] = 16'b0000000000000000;
	sram_mem[83327] = 16'b0000000000000000;
	sram_mem[83328] = 16'b0000000000000000;
	sram_mem[83329] = 16'b0000000000000000;
	sram_mem[83330] = 16'b0000000000000000;
	sram_mem[83331] = 16'b0000000000000000;
	sram_mem[83332] = 16'b0000000000000000;
	sram_mem[83333] = 16'b0000000000000000;
	sram_mem[83334] = 16'b0000000000000000;
	sram_mem[83335] = 16'b0000000000000000;
	sram_mem[83336] = 16'b0000000000000000;
	sram_mem[83337] = 16'b0000000000000000;
	sram_mem[83338] = 16'b0000000000000000;
	sram_mem[83339] = 16'b0000000000000000;
	sram_mem[83340] = 16'b0000000000000000;
	sram_mem[83341] = 16'b0000000000000000;
	sram_mem[83342] = 16'b0000000000000000;
	sram_mem[83343] = 16'b0000000000000000;
	sram_mem[83344] = 16'b0000000000000000;
	sram_mem[83345] = 16'b0000000000000000;
	sram_mem[83346] = 16'b0000000000000000;
	sram_mem[83347] = 16'b0000000000000000;
	sram_mem[83348] = 16'b0000000000000000;
	sram_mem[83349] = 16'b0000000000000000;
	sram_mem[83350] = 16'b0000000000000000;
	sram_mem[83351] = 16'b0000000000000000;
	sram_mem[83352] = 16'b0000000000000000;
	sram_mem[83353] = 16'b0000000000000000;
	sram_mem[83354] = 16'b0000000000000000;
	sram_mem[83355] = 16'b0000000000000000;
	sram_mem[83356] = 16'b0000000000000000;
	sram_mem[83357] = 16'b0000000000000000;
	sram_mem[83358] = 16'b0000000000000000;
	sram_mem[83359] = 16'b0000000000000000;
	sram_mem[83360] = 16'b0000000000000000;
	sram_mem[83361] = 16'b0000000000000000;
	sram_mem[83362] = 16'b0000000000000000;
	sram_mem[83363] = 16'b0000000000000000;
	sram_mem[83364] = 16'b0000000000000000;
	sram_mem[83365] = 16'b0000000000000000;
	sram_mem[83366] = 16'b0000000000000000;
	sram_mem[83367] = 16'b0000000000000000;
	sram_mem[83368] = 16'b0000000000000000;
	sram_mem[83369] = 16'b0000000000000000;
	sram_mem[83370] = 16'b0000000000000000;
	sram_mem[83371] = 16'b0000000000000000;
	sram_mem[83372] = 16'b0000000000000000;
	sram_mem[83373] = 16'b0000000000000000;
	sram_mem[83374] = 16'b0000000000000000;
	sram_mem[83375] = 16'b0000000000000000;
	sram_mem[83376] = 16'b0000000000000000;
	sram_mem[83377] = 16'b0000000000000000;
	sram_mem[83378] = 16'b0000000000000000;
	sram_mem[83379] = 16'b0000000000000000;
	sram_mem[83380] = 16'b0000000000000000;
	sram_mem[83381] = 16'b0000000000000000;
	sram_mem[83382] = 16'b0000000000000000;
	sram_mem[83383] = 16'b0000000000000000;
	sram_mem[83384] = 16'b0000000000000000;
	sram_mem[83385] = 16'b0000000000000000;
	sram_mem[83386] = 16'b0000000000000000;
	sram_mem[83387] = 16'b0000000000000000;
	sram_mem[83388] = 16'b0000000000000000;
	sram_mem[83389] = 16'b0000000000000000;
	sram_mem[83390] = 16'b0000000000000000;
	sram_mem[83391] = 16'b0000000000000000;
	sram_mem[83392] = 16'b0000000000000000;
	sram_mem[83393] = 16'b0000000000000000;
	sram_mem[83394] = 16'b0000000000000000;
	sram_mem[83395] = 16'b0000000000000000;
	sram_mem[83396] = 16'b0000000000000000;
	sram_mem[83397] = 16'b0000000000000000;
	sram_mem[83398] = 16'b0000000000000000;
	sram_mem[83399] = 16'b0000000000000000;
	sram_mem[83400] = 16'b0000000000000000;
	sram_mem[83401] = 16'b0000000000000000;
	sram_mem[83402] = 16'b0000000000000000;
	sram_mem[83403] = 16'b0000000000000000;
	sram_mem[83404] = 16'b0000000000000000;
	sram_mem[83405] = 16'b0000000000000000;
	sram_mem[83406] = 16'b0000000000000000;
	sram_mem[83407] = 16'b0000000000000000;
	sram_mem[83408] = 16'b0000000000000000;
	sram_mem[83409] = 16'b0000000000000000;
	sram_mem[83410] = 16'b0000000000000000;
	sram_mem[83411] = 16'b0000000000000000;
	sram_mem[83412] = 16'b0000000000000000;
	sram_mem[83413] = 16'b0000000000000000;
	sram_mem[83414] = 16'b0000000000000000;
	sram_mem[83415] = 16'b0000000000000000;
	sram_mem[83416] = 16'b0000000000000000;
	sram_mem[83417] = 16'b0000000000000000;
	sram_mem[83418] = 16'b0000000000000000;
	sram_mem[83419] = 16'b0000000000000000;
	sram_mem[83420] = 16'b0000000000000000;
	sram_mem[83421] = 16'b0000000000000000;
	sram_mem[83422] = 16'b0000000000000000;
	sram_mem[83423] = 16'b0000000000000000;
	sram_mem[83424] = 16'b0000000000000000;
	sram_mem[83425] = 16'b0000000000000000;
	sram_mem[83426] = 16'b0000000000000000;
	sram_mem[83427] = 16'b0000000000000000;
	sram_mem[83428] = 16'b0000000000000000;
	sram_mem[83429] = 16'b0000000000000000;
	sram_mem[83430] = 16'b0000000000000000;
	sram_mem[83431] = 16'b0000000000000000;
	sram_mem[83432] = 16'b0000000000000000;
	sram_mem[83433] = 16'b0000000000000000;
	sram_mem[83434] = 16'b0000000000000000;
	sram_mem[83435] = 16'b0000000000000000;
	sram_mem[83436] = 16'b0000000000000000;
	sram_mem[83437] = 16'b0000000000000000;
	sram_mem[83438] = 16'b0000000000000000;
	sram_mem[83439] = 16'b0000000000000000;
	sram_mem[83440] = 16'b0000000000000000;
	sram_mem[83441] = 16'b0000000000000000;
	sram_mem[83442] = 16'b0000000000000000;
	sram_mem[83443] = 16'b0000000000000000;
	sram_mem[83444] = 16'b0000000000000000;
	sram_mem[83445] = 16'b0000000000000000;
	sram_mem[83446] = 16'b0000000000000000;
	sram_mem[83447] = 16'b0000000000000000;
	sram_mem[83448] = 16'b0000000000000000;
	sram_mem[83449] = 16'b0000000000000000;
	sram_mem[83450] = 16'b0000000000000000;
	sram_mem[83451] = 16'b0000000000000000;
	sram_mem[83452] = 16'b0000000000000000;
	sram_mem[83453] = 16'b0000000000000000;
	sram_mem[83454] = 16'b0000000000000000;
	sram_mem[83455] = 16'b0000000000000000;
	sram_mem[83456] = 16'b0000000000000000;
	sram_mem[83457] = 16'b0000000000000000;
	sram_mem[83458] = 16'b0000000000000000;
	sram_mem[83459] = 16'b0000000000000000;
	sram_mem[83460] = 16'b0000000000000000;
	sram_mem[83461] = 16'b0000000000000000;
	sram_mem[83462] = 16'b0000000000000000;
	sram_mem[83463] = 16'b0000000000000000;
	sram_mem[83464] = 16'b0000000000000000;
	sram_mem[83465] = 16'b0000000000000000;
	sram_mem[83466] = 16'b0000000000000000;
	sram_mem[83467] = 16'b0000000000000000;
	sram_mem[83468] = 16'b0000000000000000;
	sram_mem[83469] = 16'b0000000000000000;
	sram_mem[83470] = 16'b0000000000000000;
	sram_mem[83471] = 16'b0000000000000000;
	sram_mem[83472] = 16'b0000000000000000;
	sram_mem[83473] = 16'b0000000000000000;
	sram_mem[83474] = 16'b0000000000000000;
	sram_mem[83475] = 16'b0000000000000000;
	sram_mem[83476] = 16'b0000000000000000;
	sram_mem[83477] = 16'b0000000000000000;
	sram_mem[83478] = 16'b0000000000000000;
	sram_mem[83479] = 16'b0000000000000000;
	sram_mem[83480] = 16'b0000000000000000;
	sram_mem[83481] = 16'b0000000000000000;
	sram_mem[83482] = 16'b0000000000000000;
	sram_mem[83483] = 16'b0000000000000000;
	sram_mem[83484] = 16'b0000000000000000;
	sram_mem[83485] = 16'b0000000000000000;
	sram_mem[83486] = 16'b0000000000000000;
	sram_mem[83487] = 16'b0000000000000000;
	sram_mem[83488] = 16'b0000000000000000;
	sram_mem[83489] = 16'b0000000000000000;
	sram_mem[83490] = 16'b0000000000000000;
	sram_mem[83491] = 16'b0000000000000000;
	sram_mem[83492] = 16'b0000000000000000;
	sram_mem[83493] = 16'b0000000000000000;
	sram_mem[83494] = 16'b0000000000000000;
	sram_mem[83495] = 16'b0000000000000000;
	sram_mem[83496] = 16'b0000000000000000;
	sram_mem[83497] = 16'b0000000000000000;
	sram_mem[83498] = 16'b0000000000000000;
	sram_mem[83499] = 16'b0000000000000000;
	sram_mem[83500] = 16'b0000000000000000;
	sram_mem[83501] = 16'b0000000000000000;
	sram_mem[83502] = 16'b0000000000000000;
	sram_mem[83503] = 16'b0000000000000000;
	sram_mem[83504] = 16'b0000000000000000;
	sram_mem[83505] = 16'b0000000000000000;
	sram_mem[83506] = 16'b0000000000000000;
	sram_mem[83507] = 16'b0000000000000000;
	sram_mem[83508] = 16'b0000000000000000;
	sram_mem[83509] = 16'b0000000000000000;
	sram_mem[83510] = 16'b0000000000000000;
	sram_mem[83511] = 16'b0000000000000000;
	sram_mem[83512] = 16'b0000000000000000;
	sram_mem[83513] = 16'b0000000000000000;
	sram_mem[83514] = 16'b0000000000000000;
	sram_mem[83515] = 16'b0000000000000000;
	sram_mem[83516] = 16'b0000000000000000;
	sram_mem[83517] = 16'b0000000000000000;
	sram_mem[83518] = 16'b0000000000000000;
	sram_mem[83519] = 16'b0000000000000000;
	sram_mem[83520] = 16'b0000000000000000;
	sram_mem[83521] = 16'b0000000000000000;
	sram_mem[83522] = 16'b0000000000000000;
	sram_mem[83523] = 16'b0000000000000000;
	sram_mem[83524] = 16'b0000000000000000;
	sram_mem[83525] = 16'b0000000000000000;
	sram_mem[83526] = 16'b0000000000000000;
	sram_mem[83527] = 16'b0000000000000000;
	sram_mem[83528] = 16'b0000000000000000;
	sram_mem[83529] = 16'b0000000000000000;
	sram_mem[83530] = 16'b0000000000000000;
	sram_mem[83531] = 16'b0000000000000000;
	sram_mem[83532] = 16'b0000000000000000;
	sram_mem[83533] = 16'b0000000000000000;
	sram_mem[83534] = 16'b0000000000000000;
	sram_mem[83535] = 16'b0000000000000000;
	sram_mem[83536] = 16'b0000000000000000;
	sram_mem[83537] = 16'b0000000000000000;
	sram_mem[83538] = 16'b0000000000000000;
	sram_mem[83539] = 16'b0000000000000000;
	sram_mem[83540] = 16'b0000000000000000;
	sram_mem[83541] = 16'b0000000000000000;
	sram_mem[83542] = 16'b0000000000000000;
	sram_mem[83543] = 16'b0000000000000000;
	sram_mem[83544] = 16'b0000000000000000;
	sram_mem[83545] = 16'b0000000000000000;
	sram_mem[83546] = 16'b0000000000000000;
	sram_mem[83547] = 16'b0000000000000000;
	sram_mem[83548] = 16'b0000000000000000;
	sram_mem[83549] = 16'b0000000000000000;
	sram_mem[83550] = 16'b0000000000000000;
	sram_mem[83551] = 16'b0000000000000000;
	sram_mem[83552] = 16'b0000000000000000;
	sram_mem[83553] = 16'b0000000000000000;
	sram_mem[83554] = 16'b0000000000000000;
	sram_mem[83555] = 16'b0000000000000000;
	sram_mem[83556] = 16'b0000000000000000;
	sram_mem[83557] = 16'b0000000000000000;
	sram_mem[83558] = 16'b0000000000000000;
	sram_mem[83559] = 16'b0000000000000000;
	sram_mem[83560] = 16'b0000000000000000;
	sram_mem[83561] = 16'b0000000000000000;
	sram_mem[83562] = 16'b0000000000000000;
	sram_mem[83563] = 16'b0000000000000000;
	sram_mem[83564] = 16'b0000000000000000;
	sram_mem[83565] = 16'b0000000000000000;
	sram_mem[83566] = 16'b0000000000000000;
	sram_mem[83567] = 16'b0000000000000000;
	sram_mem[83568] = 16'b0000000000000000;
	sram_mem[83569] = 16'b0000000000000000;
	sram_mem[83570] = 16'b0000000000000000;
	sram_mem[83571] = 16'b0000000000000000;
	sram_mem[83572] = 16'b0000000000000000;
	sram_mem[83573] = 16'b0000000000000000;
	sram_mem[83574] = 16'b0000000000000000;
	sram_mem[83575] = 16'b0000000000000000;
	sram_mem[83576] = 16'b0000000000000000;
	sram_mem[83577] = 16'b0000000000000000;
	sram_mem[83578] = 16'b0000000000000000;
	sram_mem[83579] = 16'b0000000000000000;
	sram_mem[83580] = 16'b0000000000000000;
	sram_mem[83581] = 16'b0000000000000000;
	sram_mem[83582] = 16'b0000000000000000;
	sram_mem[83583] = 16'b0000000000000000;
	sram_mem[83584] = 16'b0000000000000000;
	sram_mem[83585] = 16'b0000000000000000;
	sram_mem[83586] = 16'b0000000000000000;
	sram_mem[83587] = 16'b0000000000000000;
	sram_mem[83588] = 16'b0000000000000000;
	sram_mem[83589] = 16'b0000000000000000;
	sram_mem[83590] = 16'b0000000000000000;
	sram_mem[83591] = 16'b0000000000000000;
	sram_mem[83592] = 16'b0000000000000000;
	sram_mem[83593] = 16'b0000000000000000;
	sram_mem[83594] = 16'b0000000000000000;
	sram_mem[83595] = 16'b0000000000000000;
	sram_mem[83596] = 16'b0000000000000000;
	sram_mem[83597] = 16'b0000000000000000;
	sram_mem[83598] = 16'b0000000000000000;
	sram_mem[83599] = 16'b0000000000000000;
	sram_mem[83600] = 16'b0000000000000000;
	sram_mem[83601] = 16'b0000000000000000;
	sram_mem[83602] = 16'b0000000000000000;
	sram_mem[83603] = 16'b0000000000000000;
	sram_mem[83604] = 16'b0000000000000000;
	sram_mem[83605] = 16'b0000000000000000;
	sram_mem[83606] = 16'b0000000000000000;
	sram_mem[83607] = 16'b0000000000000000;
	sram_mem[83608] = 16'b0000000000000000;
	sram_mem[83609] = 16'b0000000000000000;
	sram_mem[83610] = 16'b0000000000000000;
	sram_mem[83611] = 16'b0000000000000000;
	sram_mem[83612] = 16'b0000000000000000;
	sram_mem[83613] = 16'b0000000000000000;
	sram_mem[83614] = 16'b0000000000000000;
	sram_mem[83615] = 16'b0000000000000000;
	sram_mem[83616] = 16'b0000000000000000;
	sram_mem[83617] = 16'b0000000000000000;
	sram_mem[83618] = 16'b0000000000000000;
	sram_mem[83619] = 16'b0000000000000000;
	sram_mem[83620] = 16'b0000000000000000;
	sram_mem[83621] = 16'b0000000000000000;
	sram_mem[83622] = 16'b0000000000000000;
	sram_mem[83623] = 16'b0000000000000000;
	sram_mem[83624] = 16'b0000000000000000;
	sram_mem[83625] = 16'b0000000000000000;
	sram_mem[83626] = 16'b0000000000000000;
	sram_mem[83627] = 16'b0000000000000000;
	sram_mem[83628] = 16'b0000000000000000;
	sram_mem[83629] = 16'b0000000000000000;
	sram_mem[83630] = 16'b0000000000000000;
	sram_mem[83631] = 16'b0000000000000000;
	sram_mem[83632] = 16'b0000000000000000;
	sram_mem[83633] = 16'b0000000000000000;
	sram_mem[83634] = 16'b0000000000000000;
	sram_mem[83635] = 16'b0000000000000000;
	sram_mem[83636] = 16'b0000000000000000;
	sram_mem[83637] = 16'b0000000000000000;
	sram_mem[83638] = 16'b0000000000000000;
	sram_mem[83639] = 16'b0000000000000000;
	sram_mem[83640] = 16'b0000000000000000;
	sram_mem[83641] = 16'b0000000000000000;
	sram_mem[83642] = 16'b0000000000000000;
	sram_mem[83643] = 16'b0000000000000000;
	sram_mem[83644] = 16'b0000000000000000;
	sram_mem[83645] = 16'b0000000000000000;
	sram_mem[83646] = 16'b0000000000000000;
	sram_mem[83647] = 16'b0000000000000000;
	sram_mem[83648] = 16'b0000000000000000;
	sram_mem[83649] = 16'b0000000000000000;
	sram_mem[83650] = 16'b0000000000000000;
	sram_mem[83651] = 16'b0000000000000000;
	sram_mem[83652] = 16'b0000000000000000;
	sram_mem[83653] = 16'b0000000000000000;
	sram_mem[83654] = 16'b0000000000000000;
	sram_mem[83655] = 16'b0000000000000000;
	sram_mem[83656] = 16'b0000000000000000;
	sram_mem[83657] = 16'b0000000000000000;
	sram_mem[83658] = 16'b0000000000000000;
	sram_mem[83659] = 16'b0000000000000000;
	sram_mem[83660] = 16'b0000000000000000;
	sram_mem[83661] = 16'b0000000000000000;
	sram_mem[83662] = 16'b0000000000000000;
	sram_mem[83663] = 16'b0000000000000000;
	sram_mem[83664] = 16'b0000000000000000;
	sram_mem[83665] = 16'b0000000000000000;
	sram_mem[83666] = 16'b0000000000000000;
	sram_mem[83667] = 16'b0000000000000000;
	sram_mem[83668] = 16'b0000000000000000;
	sram_mem[83669] = 16'b0000000000000000;
	sram_mem[83670] = 16'b0000000000000000;
	sram_mem[83671] = 16'b0000000000000000;
	sram_mem[83672] = 16'b0000000000000000;
	sram_mem[83673] = 16'b0000000000000000;
	sram_mem[83674] = 16'b0000000000000000;
	sram_mem[83675] = 16'b0000000000000000;
	sram_mem[83676] = 16'b0000000000000000;
	sram_mem[83677] = 16'b0000000000000000;
	sram_mem[83678] = 16'b0000000000000000;
	sram_mem[83679] = 16'b0000000000000000;
	sram_mem[83680] = 16'b0000000000000000;
	sram_mem[83681] = 16'b0000000000000000;
	sram_mem[83682] = 16'b0000000000000000;
	sram_mem[83683] = 16'b0000000000000000;
	sram_mem[83684] = 16'b0000000000000000;
	sram_mem[83685] = 16'b0000000000000000;
	sram_mem[83686] = 16'b0000000000000000;
	sram_mem[83687] = 16'b0000000000000000;
	sram_mem[83688] = 16'b0000000000000000;
	sram_mem[83689] = 16'b0000000000000000;
	sram_mem[83690] = 16'b0000000000000000;
	sram_mem[83691] = 16'b0000000000000000;
	sram_mem[83692] = 16'b0000000000000000;
	sram_mem[83693] = 16'b0000000000000000;
	sram_mem[83694] = 16'b0000000000000000;
	sram_mem[83695] = 16'b0000000000000000;
	sram_mem[83696] = 16'b0000000000000000;
	sram_mem[83697] = 16'b0000000000000000;
	sram_mem[83698] = 16'b0000000000000000;
	sram_mem[83699] = 16'b0000000000000000;
	sram_mem[83700] = 16'b0000000000000000;
	sram_mem[83701] = 16'b0000000000000000;
	sram_mem[83702] = 16'b0000000000000000;
	sram_mem[83703] = 16'b0000000000000000;
	sram_mem[83704] = 16'b0000000000000000;
	sram_mem[83705] = 16'b0000000000000000;
	sram_mem[83706] = 16'b0000000000000000;
	sram_mem[83707] = 16'b0000000000000000;
	sram_mem[83708] = 16'b0000000000000000;
	sram_mem[83709] = 16'b0000000000000000;
	sram_mem[83710] = 16'b0000000000000000;
	sram_mem[83711] = 16'b0000000000000000;
	sram_mem[83712] = 16'b0000000000000000;
	sram_mem[83713] = 16'b0000000000000000;
	sram_mem[83714] = 16'b0000000000000000;
	sram_mem[83715] = 16'b0000000000000000;
	sram_mem[83716] = 16'b0000000000000000;
	sram_mem[83717] = 16'b0000000000000000;
	sram_mem[83718] = 16'b0000000000000000;
	sram_mem[83719] = 16'b0000000000000000;
	sram_mem[83720] = 16'b0000000000000000;
	sram_mem[83721] = 16'b0000000000000000;
	sram_mem[83722] = 16'b0000000000000000;
	sram_mem[83723] = 16'b0000000000000000;
	sram_mem[83724] = 16'b0000000000000000;
	sram_mem[83725] = 16'b0000000000000000;
	sram_mem[83726] = 16'b0000000000000000;
	sram_mem[83727] = 16'b0000000000000000;
	sram_mem[83728] = 16'b0000000000000000;
	sram_mem[83729] = 16'b0000000000000000;
	sram_mem[83730] = 16'b0000000000000000;
	sram_mem[83731] = 16'b0000000000000000;
	sram_mem[83732] = 16'b0000000000000000;
	sram_mem[83733] = 16'b0000000000000000;
	sram_mem[83734] = 16'b0000000000000000;
	sram_mem[83735] = 16'b0000000000000000;
	sram_mem[83736] = 16'b0000000000000000;
	sram_mem[83737] = 16'b0000000000000000;
	sram_mem[83738] = 16'b0000000000000000;
	sram_mem[83739] = 16'b0000000000000000;
	sram_mem[83740] = 16'b0000000000000000;
	sram_mem[83741] = 16'b0000000000000000;
	sram_mem[83742] = 16'b0000000000000000;
	sram_mem[83743] = 16'b0000000000000000;
	sram_mem[83744] = 16'b0000000000000000;
	sram_mem[83745] = 16'b0000000000000000;
	sram_mem[83746] = 16'b0000000000000000;
	sram_mem[83747] = 16'b0000000000000000;
	sram_mem[83748] = 16'b0000000000000000;
	sram_mem[83749] = 16'b0000000000000000;
	sram_mem[83750] = 16'b0000000000000000;
	sram_mem[83751] = 16'b0000000000000000;
	sram_mem[83752] = 16'b0000000000000000;
	sram_mem[83753] = 16'b0000000000000000;
	sram_mem[83754] = 16'b0000000000000000;
	sram_mem[83755] = 16'b0000000000000000;
	sram_mem[83756] = 16'b0000000000000000;
	sram_mem[83757] = 16'b0000000000000000;
	sram_mem[83758] = 16'b0000000000000000;
	sram_mem[83759] = 16'b0000000000000000;
	sram_mem[83760] = 16'b0000000000000000;
	sram_mem[83761] = 16'b0000000000000000;
	sram_mem[83762] = 16'b0000000000000000;
	sram_mem[83763] = 16'b0000000000000000;
	sram_mem[83764] = 16'b0000000000000000;
	sram_mem[83765] = 16'b0000000000000000;
	sram_mem[83766] = 16'b0000000000000000;
	sram_mem[83767] = 16'b0000000000000000;
	sram_mem[83768] = 16'b0000000000000000;
	sram_mem[83769] = 16'b0000000000000000;
	sram_mem[83770] = 16'b0000000000000000;
	sram_mem[83771] = 16'b0000000000000000;
	sram_mem[83772] = 16'b0000000000000000;
	sram_mem[83773] = 16'b0000000000000000;
	sram_mem[83774] = 16'b0000000000000000;
	sram_mem[83775] = 16'b0000000000000000;
	sram_mem[83776] = 16'b0000000000000000;
	sram_mem[83777] = 16'b0000000000000000;
	sram_mem[83778] = 16'b0000000000000000;
	sram_mem[83779] = 16'b0000000000000000;
	sram_mem[83780] = 16'b0000000000000000;
	sram_mem[83781] = 16'b0000000000000000;
	sram_mem[83782] = 16'b0000000000000000;
	sram_mem[83783] = 16'b0000000000000000;
	sram_mem[83784] = 16'b0000000000000000;
	sram_mem[83785] = 16'b0000000000000000;
	sram_mem[83786] = 16'b0000000000000000;
	sram_mem[83787] = 16'b0000000000000000;
	sram_mem[83788] = 16'b0000000000000000;
	sram_mem[83789] = 16'b0000000000000000;
	sram_mem[83790] = 16'b0000000000000000;
	sram_mem[83791] = 16'b0000000000000000;
	sram_mem[83792] = 16'b0000000000000000;
	sram_mem[83793] = 16'b0000000000000000;
	sram_mem[83794] = 16'b0000000000000000;
	sram_mem[83795] = 16'b0000000000000000;
	sram_mem[83796] = 16'b0000000000000000;
	sram_mem[83797] = 16'b0000000000000000;
	sram_mem[83798] = 16'b0000000000000000;
	sram_mem[83799] = 16'b0000000000000000;
	sram_mem[83800] = 16'b0000000000000000;
	sram_mem[83801] = 16'b0000000000000000;
	sram_mem[83802] = 16'b0000000000000000;
	sram_mem[83803] = 16'b0000000000000000;
	sram_mem[83804] = 16'b0000000000000000;
	sram_mem[83805] = 16'b0000000000000000;
	sram_mem[83806] = 16'b0000000000000000;
	sram_mem[83807] = 16'b0000000000000000;
	sram_mem[83808] = 16'b0000000000000000;
	sram_mem[83809] = 16'b0000000000000000;
	sram_mem[83810] = 16'b0000000000000000;
	sram_mem[83811] = 16'b0000000000000000;
	sram_mem[83812] = 16'b0000000000000000;
	sram_mem[83813] = 16'b0000000000000000;
	sram_mem[83814] = 16'b0000000000000000;
	sram_mem[83815] = 16'b0000000000000000;
	sram_mem[83816] = 16'b0000000000000000;
	sram_mem[83817] = 16'b0000000000000000;
	sram_mem[83818] = 16'b0000000000000000;
	sram_mem[83819] = 16'b0000000000000000;
	sram_mem[83820] = 16'b0000000000000000;
	sram_mem[83821] = 16'b0000000000000000;
	sram_mem[83822] = 16'b0000000000000000;
	sram_mem[83823] = 16'b0000000000000000;
	sram_mem[83824] = 16'b0000000000000000;
	sram_mem[83825] = 16'b0000000000000000;
	sram_mem[83826] = 16'b0000000000000000;
	sram_mem[83827] = 16'b0000000000000000;
	sram_mem[83828] = 16'b0000000000000000;
	sram_mem[83829] = 16'b0000000000000000;
	sram_mem[83830] = 16'b0000000000000000;
	sram_mem[83831] = 16'b0000000000000000;
	sram_mem[83832] = 16'b0000000000000000;
	sram_mem[83833] = 16'b0000000000000000;
	sram_mem[83834] = 16'b0000000000000000;
	sram_mem[83835] = 16'b0000000000000000;
	sram_mem[83836] = 16'b0000000000000000;
	sram_mem[83837] = 16'b0000000000000000;
	sram_mem[83838] = 16'b0000000000000000;
	sram_mem[83839] = 16'b0000000000000000;
	sram_mem[83840] = 16'b0000000000000000;
	sram_mem[83841] = 16'b0000000000000000;
	sram_mem[83842] = 16'b0000000000000000;
	sram_mem[83843] = 16'b0000000000000000;
	sram_mem[83844] = 16'b0000000000000000;
	sram_mem[83845] = 16'b0000000000000000;
	sram_mem[83846] = 16'b0000000000000000;
	sram_mem[83847] = 16'b0000000000000000;
	sram_mem[83848] = 16'b0000000000000000;
	sram_mem[83849] = 16'b0000000000000000;
	sram_mem[83850] = 16'b0000000000000000;
	sram_mem[83851] = 16'b0000000000000000;
	sram_mem[83852] = 16'b0000000000000000;
	sram_mem[83853] = 16'b0000000000000000;
	sram_mem[83854] = 16'b0000000000000000;
	sram_mem[83855] = 16'b0000000000000000;
	sram_mem[83856] = 16'b0000000000000000;
	sram_mem[83857] = 16'b0000000000000000;
	sram_mem[83858] = 16'b0000000000000000;
	sram_mem[83859] = 16'b0000000000000000;
	sram_mem[83860] = 16'b0000000000000000;
	sram_mem[83861] = 16'b0000000000000000;
	sram_mem[83862] = 16'b0000000000000000;
	sram_mem[83863] = 16'b0000000000000000;
	sram_mem[83864] = 16'b0000000000000000;
	sram_mem[83865] = 16'b0000000000000000;
	sram_mem[83866] = 16'b0000000000000000;
	sram_mem[83867] = 16'b0000000000000000;
	sram_mem[83868] = 16'b0000000000000000;
	sram_mem[83869] = 16'b0000000000000000;
	sram_mem[83870] = 16'b0000000000000000;
	sram_mem[83871] = 16'b0000000000000000;
	sram_mem[83872] = 16'b0000000000000000;
	sram_mem[83873] = 16'b0000000000000000;
	sram_mem[83874] = 16'b0000000000000000;
	sram_mem[83875] = 16'b0000000000000000;
	sram_mem[83876] = 16'b0000000000000000;
	sram_mem[83877] = 16'b0000000000000000;
	sram_mem[83878] = 16'b0000000000000000;
	sram_mem[83879] = 16'b0000000000000000;
	sram_mem[83880] = 16'b0000000000000000;
	sram_mem[83881] = 16'b0000000000000000;
	sram_mem[83882] = 16'b0000000000000000;
	sram_mem[83883] = 16'b0000000000000000;
	sram_mem[83884] = 16'b0000000000000000;
	sram_mem[83885] = 16'b0000000000000000;
	sram_mem[83886] = 16'b0000000000000000;
	sram_mem[83887] = 16'b0000000000000000;
	sram_mem[83888] = 16'b0000000000000000;
	sram_mem[83889] = 16'b0000000000000000;
	sram_mem[83890] = 16'b0000000000000000;
	sram_mem[83891] = 16'b0000000000000000;
	sram_mem[83892] = 16'b0000000000000000;
	sram_mem[83893] = 16'b0000000000000000;
	sram_mem[83894] = 16'b0000000000000000;
	sram_mem[83895] = 16'b0000000000000000;
	sram_mem[83896] = 16'b0000000000000000;
	sram_mem[83897] = 16'b0000000000000000;
	sram_mem[83898] = 16'b0000000000000000;
	sram_mem[83899] = 16'b0000000000000000;
	sram_mem[83900] = 16'b0000000000000000;
	sram_mem[83901] = 16'b0000000000000000;
	sram_mem[83902] = 16'b0000000000000000;
	sram_mem[83903] = 16'b0000000000000000;
	sram_mem[83904] = 16'b0000000000000000;
	sram_mem[83905] = 16'b0000000000000000;
	sram_mem[83906] = 16'b0000000000000000;
	sram_mem[83907] = 16'b0000000000000000;
	sram_mem[83908] = 16'b0000000000000000;
	sram_mem[83909] = 16'b0000000000000000;
	sram_mem[83910] = 16'b0000000000000000;
	sram_mem[83911] = 16'b0000000000000000;
	sram_mem[83912] = 16'b0000000000000000;
	sram_mem[83913] = 16'b0000000000000000;
	sram_mem[83914] = 16'b0000000000000000;
	sram_mem[83915] = 16'b0000000000000000;
	sram_mem[83916] = 16'b0000000000000000;
	sram_mem[83917] = 16'b0000000000000000;
	sram_mem[83918] = 16'b0000000000000000;
	sram_mem[83919] = 16'b0000000000000000;
	sram_mem[83920] = 16'b0000000000000000;
	sram_mem[83921] = 16'b0000000000000000;
	sram_mem[83922] = 16'b0000000000000000;
	sram_mem[83923] = 16'b0000000000000000;
	sram_mem[83924] = 16'b0000000000000000;
	sram_mem[83925] = 16'b0000000000000000;
	sram_mem[83926] = 16'b0000000000000000;
	sram_mem[83927] = 16'b0000000000000000;
	sram_mem[83928] = 16'b0000000000000000;
	sram_mem[83929] = 16'b0000000000000000;
	sram_mem[83930] = 16'b0000000000000000;
	sram_mem[83931] = 16'b0000000000000000;
	sram_mem[83932] = 16'b0000000000000000;
	sram_mem[83933] = 16'b0000000000000000;
	sram_mem[83934] = 16'b0000000000000000;
	sram_mem[83935] = 16'b0000000000000000;
	sram_mem[83936] = 16'b0000000000000000;
	sram_mem[83937] = 16'b0000000000000000;
	sram_mem[83938] = 16'b0000000000000000;
	sram_mem[83939] = 16'b0000000000000000;
	sram_mem[83940] = 16'b0000000000000000;
	sram_mem[83941] = 16'b0000000000000000;
	sram_mem[83942] = 16'b0000000000000000;
	sram_mem[83943] = 16'b0000000000000000;
	sram_mem[83944] = 16'b0000000000000000;
	sram_mem[83945] = 16'b0000000000000000;
	sram_mem[83946] = 16'b0000000000000000;
	sram_mem[83947] = 16'b0000000000000000;
	sram_mem[83948] = 16'b0000000000000000;
	sram_mem[83949] = 16'b0000000000000000;
	sram_mem[83950] = 16'b0000000000000000;
	sram_mem[83951] = 16'b0000000000000000;
	sram_mem[83952] = 16'b0000000000000000;
	sram_mem[83953] = 16'b0000000000000000;
	sram_mem[83954] = 16'b0000000000000000;
	sram_mem[83955] = 16'b0000000000000000;
	sram_mem[83956] = 16'b0000000000000000;
	sram_mem[83957] = 16'b0000000000000000;
	sram_mem[83958] = 16'b0000000000000000;
	sram_mem[83959] = 16'b0000000000000000;
	sram_mem[83960] = 16'b0000000000000000;
	sram_mem[83961] = 16'b0000000000000000;
	sram_mem[83962] = 16'b0000000000000000;
	sram_mem[83963] = 16'b0000000000000000;
	sram_mem[83964] = 16'b0000000000000000;
	sram_mem[83965] = 16'b0000000000000000;
	sram_mem[83966] = 16'b0000000000000000;
	sram_mem[83967] = 16'b0000000000000000;
	sram_mem[83968] = 16'b0000000000000000;
	sram_mem[83969] = 16'b0000000000000000;
	sram_mem[83970] = 16'b0000000000000000;
	sram_mem[83971] = 16'b0000000000000000;
	sram_mem[83972] = 16'b0000000000000000;
	sram_mem[83973] = 16'b0000000000000000;
	sram_mem[83974] = 16'b0000000000000000;
	sram_mem[83975] = 16'b0000000000000000;
	sram_mem[83976] = 16'b0000000000000000;
	sram_mem[83977] = 16'b0000000000000000;
	sram_mem[83978] = 16'b0000000000000000;
	sram_mem[83979] = 16'b0000000000000000;
	sram_mem[83980] = 16'b0000000000000000;
	sram_mem[83981] = 16'b0000000000000000;
	sram_mem[83982] = 16'b0000000000000000;
	sram_mem[83983] = 16'b0000000000000000;
	sram_mem[83984] = 16'b0000000000000000;
	sram_mem[83985] = 16'b0000000000000000;
	sram_mem[83986] = 16'b0000000000000000;
	sram_mem[83987] = 16'b0000000000000000;
	sram_mem[83988] = 16'b0000000000000000;
	sram_mem[83989] = 16'b0000000000000000;
	sram_mem[83990] = 16'b0000000000000000;
	sram_mem[83991] = 16'b0000000000000000;
	sram_mem[83992] = 16'b0000000000000000;
	sram_mem[83993] = 16'b0000000000000000;
	sram_mem[83994] = 16'b0000000000000000;
	sram_mem[83995] = 16'b0000000000000000;
	sram_mem[83996] = 16'b0000000000000000;
	sram_mem[83997] = 16'b0000000000000000;
	sram_mem[83998] = 16'b0000000000000000;
	sram_mem[83999] = 16'b0000000000000000;
	sram_mem[84000] = 16'b0000000000000000;
	sram_mem[84001] = 16'b0000000000000000;
	sram_mem[84002] = 16'b0000000000000000;
	sram_mem[84003] = 16'b0000000000000000;
	sram_mem[84004] = 16'b0000000000000000;
	sram_mem[84005] = 16'b0000000000000000;
	sram_mem[84006] = 16'b0000000000000000;
	sram_mem[84007] = 16'b0000000000000000;
	sram_mem[84008] = 16'b0000000000000000;
	sram_mem[84009] = 16'b0000000000000000;
	sram_mem[84010] = 16'b0000000000000000;
	sram_mem[84011] = 16'b0000000000000000;
	sram_mem[84012] = 16'b0000000000000000;
	sram_mem[84013] = 16'b0000000000000000;
	sram_mem[84014] = 16'b0000000000000000;
	sram_mem[84015] = 16'b0000000000000000;
	sram_mem[84016] = 16'b0000000000000000;
	sram_mem[84017] = 16'b0000000000000000;
	sram_mem[84018] = 16'b0000000000000000;
	sram_mem[84019] = 16'b0000000000000000;
	sram_mem[84020] = 16'b0000000000000000;
	sram_mem[84021] = 16'b0000000000000000;
	sram_mem[84022] = 16'b0000000000000000;
	sram_mem[84023] = 16'b0000000000000000;
	sram_mem[84024] = 16'b0000000000000000;
	sram_mem[84025] = 16'b0000000000000000;
	sram_mem[84026] = 16'b0000000000000000;
	sram_mem[84027] = 16'b0000000000000000;
	sram_mem[84028] = 16'b0000000000000000;
	sram_mem[84029] = 16'b0000000000000000;
	sram_mem[84030] = 16'b0000000000000000;
	sram_mem[84031] = 16'b0000000000000000;
	sram_mem[84032] = 16'b0000000000000000;
	sram_mem[84033] = 16'b0000000000000000;
	sram_mem[84034] = 16'b0000000000000000;
	sram_mem[84035] = 16'b0000000000000000;
	sram_mem[84036] = 16'b0000000000000000;
	sram_mem[84037] = 16'b0000000000000000;
	sram_mem[84038] = 16'b0000000000000000;
	sram_mem[84039] = 16'b0000000000000000;
	sram_mem[84040] = 16'b0000000000000000;
	sram_mem[84041] = 16'b0000000000000000;
	sram_mem[84042] = 16'b0000000000000000;
	sram_mem[84043] = 16'b0000000000000000;
	sram_mem[84044] = 16'b0000000000000000;
	sram_mem[84045] = 16'b0000000000000000;
	sram_mem[84046] = 16'b0000000000000000;
	sram_mem[84047] = 16'b0000000000000000;
	sram_mem[84048] = 16'b0000000000000000;
	sram_mem[84049] = 16'b0000000000000000;
	sram_mem[84050] = 16'b0000000000000000;
	sram_mem[84051] = 16'b0000000000000000;
	sram_mem[84052] = 16'b0000000000000000;
	sram_mem[84053] = 16'b0000000000000000;
	sram_mem[84054] = 16'b0000000000000000;
	sram_mem[84055] = 16'b0000000000000000;
	sram_mem[84056] = 16'b0000000000000000;
	sram_mem[84057] = 16'b0000000000000000;
	sram_mem[84058] = 16'b0000000000000000;
	sram_mem[84059] = 16'b0000000000000000;
	sram_mem[84060] = 16'b0000000000000000;
	sram_mem[84061] = 16'b0000000000000000;
	sram_mem[84062] = 16'b0000000000000000;
	sram_mem[84063] = 16'b0000000000000000;
	sram_mem[84064] = 16'b0000000000000000;
	sram_mem[84065] = 16'b0000000000000000;
	sram_mem[84066] = 16'b0000000000000000;
	sram_mem[84067] = 16'b0000000000000000;
	sram_mem[84068] = 16'b0000000000000000;
	sram_mem[84069] = 16'b0000000000000000;
	sram_mem[84070] = 16'b0000000000000000;
	sram_mem[84071] = 16'b0000000000000000;
	sram_mem[84072] = 16'b0000000000000000;
	sram_mem[84073] = 16'b0000000000000000;
	sram_mem[84074] = 16'b0000000000000000;
	sram_mem[84075] = 16'b0000000000000000;
	sram_mem[84076] = 16'b0000000000000000;
	sram_mem[84077] = 16'b0000000000000000;
	sram_mem[84078] = 16'b0000000000000000;
	sram_mem[84079] = 16'b0000000000000000;
	sram_mem[84080] = 16'b0000000000000000;
	sram_mem[84081] = 16'b0000000000000000;
	sram_mem[84082] = 16'b0000000000000000;
	sram_mem[84083] = 16'b0000000000000000;
	sram_mem[84084] = 16'b0000000000000000;
	sram_mem[84085] = 16'b0000000000000000;
	sram_mem[84086] = 16'b0000000000000000;
	sram_mem[84087] = 16'b0000000000000000;
	sram_mem[84088] = 16'b0000000000000000;
	sram_mem[84089] = 16'b0000000000000000;
	sram_mem[84090] = 16'b0000000000000000;
	sram_mem[84091] = 16'b0000000000000000;
	sram_mem[84092] = 16'b0000000000000000;
	sram_mem[84093] = 16'b0000000000000000;
	sram_mem[84094] = 16'b0000000000000000;
	sram_mem[84095] = 16'b0000000000000000;
	sram_mem[84096] = 16'b0000000000000000;
	sram_mem[84097] = 16'b0000000000000000;
	sram_mem[84098] = 16'b0000000000000000;
	sram_mem[84099] = 16'b0000000000000000;
	sram_mem[84100] = 16'b0000000000000000;
	sram_mem[84101] = 16'b0000000000000000;
	sram_mem[84102] = 16'b0000000000000000;
	sram_mem[84103] = 16'b0000000000000000;
	sram_mem[84104] = 16'b0000000000000000;
	sram_mem[84105] = 16'b0000000000000000;
	sram_mem[84106] = 16'b0000000000000000;
	sram_mem[84107] = 16'b0000000000000000;
	sram_mem[84108] = 16'b0000000000000000;
	sram_mem[84109] = 16'b0000000000000000;
	sram_mem[84110] = 16'b0000000000000000;
	sram_mem[84111] = 16'b0000000000000000;
	sram_mem[84112] = 16'b0000000000000000;
	sram_mem[84113] = 16'b0000000000000000;
	sram_mem[84114] = 16'b0000000000000000;
	sram_mem[84115] = 16'b0000000000000000;
	sram_mem[84116] = 16'b0000000000000000;
	sram_mem[84117] = 16'b0000000000000000;
	sram_mem[84118] = 16'b0000000000000000;
	sram_mem[84119] = 16'b0000000000000000;
	sram_mem[84120] = 16'b0000000000000000;
	sram_mem[84121] = 16'b0000000000000000;
	sram_mem[84122] = 16'b0000000000000000;
	sram_mem[84123] = 16'b0000000000000000;
	sram_mem[84124] = 16'b0000000000000000;
	sram_mem[84125] = 16'b0000000000000000;
	sram_mem[84126] = 16'b0000000000000000;
	sram_mem[84127] = 16'b0000000000000000;
	sram_mem[84128] = 16'b0000000000000000;
	sram_mem[84129] = 16'b0000000000000000;
	sram_mem[84130] = 16'b0000000000000000;
	sram_mem[84131] = 16'b0000000000000000;
	sram_mem[84132] = 16'b0000000000000000;
	sram_mem[84133] = 16'b0000000000000000;
	sram_mem[84134] = 16'b0000000000000000;
	sram_mem[84135] = 16'b0000000000000000;
	sram_mem[84136] = 16'b0000000000000000;
	sram_mem[84137] = 16'b0000000000000000;
	sram_mem[84138] = 16'b0000000000000000;
	sram_mem[84139] = 16'b0000000000000000;
	sram_mem[84140] = 16'b0000000000000000;
	sram_mem[84141] = 16'b0000000000000000;
	sram_mem[84142] = 16'b0000000000000000;
	sram_mem[84143] = 16'b0000000000000000;
	sram_mem[84144] = 16'b0000000000000000;
	sram_mem[84145] = 16'b0000000000000000;
	sram_mem[84146] = 16'b0000000000000000;
	sram_mem[84147] = 16'b0000000000000000;
	sram_mem[84148] = 16'b0000000000000000;
	sram_mem[84149] = 16'b0000000000000000;
	sram_mem[84150] = 16'b0000000000000000;
	sram_mem[84151] = 16'b0000000000000000;
	sram_mem[84152] = 16'b0000000000000000;
	sram_mem[84153] = 16'b0000000000000000;
	sram_mem[84154] = 16'b0000000000000000;
	sram_mem[84155] = 16'b0000000000000000;
	sram_mem[84156] = 16'b0000000000000000;
	sram_mem[84157] = 16'b0000000000000000;
	sram_mem[84158] = 16'b0000000000000000;
	sram_mem[84159] = 16'b0000000000000000;
	sram_mem[84160] = 16'b0000000000000000;
	sram_mem[84161] = 16'b0000000000000000;
	sram_mem[84162] = 16'b0000000000000000;
	sram_mem[84163] = 16'b0000000000000000;
	sram_mem[84164] = 16'b0000000000000000;
	sram_mem[84165] = 16'b0000000000000000;
	sram_mem[84166] = 16'b0000000000000000;
	sram_mem[84167] = 16'b0000000000000000;
	sram_mem[84168] = 16'b0000000000000000;
	sram_mem[84169] = 16'b0000000000000000;
	sram_mem[84170] = 16'b0000000000000000;
	sram_mem[84171] = 16'b0000000000000000;
	sram_mem[84172] = 16'b0000000000000000;
	sram_mem[84173] = 16'b0000000000000000;
	sram_mem[84174] = 16'b0000000000000000;
	sram_mem[84175] = 16'b0000000000000000;
	sram_mem[84176] = 16'b0000000000000000;
	sram_mem[84177] = 16'b0000000000000000;
	sram_mem[84178] = 16'b0000000000000000;
	sram_mem[84179] = 16'b0000000000000000;
	sram_mem[84180] = 16'b0000000000000000;
	sram_mem[84181] = 16'b0000000000000000;
	sram_mem[84182] = 16'b0000000000000000;
	sram_mem[84183] = 16'b0000000000000000;
	sram_mem[84184] = 16'b0000000000000000;
	sram_mem[84185] = 16'b0000000000000000;
	sram_mem[84186] = 16'b0000000000000000;
	sram_mem[84187] = 16'b0000000000000000;
	sram_mem[84188] = 16'b0000000000000000;
	sram_mem[84189] = 16'b0000000000000000;
	sram_mem[84190] = 16'b0000000000000000;
	sram_mem[84191] = 16'b0000000000000000;
	sram_mem[84192] = 16'b0000000000000000;
	sram_mem[84193] = 16'b0000000000000000;
	sram_mem[84194] = 16'b0000000000000000;
	sram_mem[84195] = 16'b0000000000000000;
	sram_mem[84196] = 16'b0000000000000000;
	sram_mem[84197] = 16'b0000000000000000;
	sram_mem[84198] = 16'b0000000000000000;
	sram_mem[84199] = 16'b0000000000000000;
	sram_mem[84200] = 16'b0000000000000000;
	sram_mem[84201] = 16'b0000000000000000;
	sram_mem[84202] = 16'b0000000000000000;
	sram_mem[84203] = 16'b0000000000000000;
	sram_mem[84204] = 16'b0000000000000000;
	sram_mem[84205] = 16'b0000000000000000;
	sram_mem[84206] = 16'b0000000000000000;
	sram_mem[84207] = 16'b0000000000000000;
	sram_mem[84208] = 16'b0000000000000000;
	sram_mem[84209] = 16'b0000000000000000;
	sram_mem[84210] = 16'b0000000000000000;
	sram_mem[84211] = 16'b0000000000000000;
	sram_mem[84212] = 16'b0000000000000000;
	sram_mem[84213] = 16'b0000000000000000;
	sram_mem[84214] = 16'b0000000000000000;
	sram_mem[84215] = 16'b0000000000000000;
	sram_mem[84216] = 16'b0000000000000000;
	sram_mem[84217] = 16'b0000000000000000;
	sram_mem[84218] = 16'b0000000000000000;
	sram_mem[84219] = 16'b0000000000000000;
	sram_mem[84220] = 16'b0000000000000000;
	sram_mem[84221] = 16'b0000000000000000;
	sram_mem[84222] = 16'b0000000000000000;
	sram_mem[84223] = 16'b0000000000000000;
	sram_mem[84224] = 16'b0000000000000000;
	sram_mem[84225] = 16'b0000000000000000;
	sram_mem[84226] = 16'b0000000000000000;
	sram_mem[84227] = 16'b0000000000000000;
	sram_mem[84228] = 16'b0000000000000000;
	sram_mem[84229] = 16'b0000000000000000;
	sram_mem[84230] = 16'b0000000000000000;
	sram_mem[84231] = 16'b0000000000000000;
	sram_mem[84232] = 16'b0000000000000000;
	sram_mem[84233] = 16'b0000000000000000;
	sram_mem[84234] = 16'b0000000000000000;
	sram_mem[84235] = 16'b0000000000000000;
	sram_mem[84236] = 16'b0000000000000000;
	sram_mem[84237] = 16'b0000000000000000;
	sram_mem[84238] = 16'b0000000000000000;
	sram_mem[84239] = 16'b0000000000000000;
	sram_mem[84240] = 16'b0000000000000000;
	sram_mem[84241] = 16'b0000000000000000;
	sram_mem[84242] = 16'b0000000000000000;
	sram_mem[84243] = 16'b0000000000000000;
	sram_mem[84244] = 16'b0000000000000000;
	sram_mem[84245] = 16'b0000000000000000;
	sram_mem[84246] = 16'b0000000000000000;
	sram_mem[84247] = 16'b0000000000000000;
	sram_mem[84248] = 16'b0000000000000000;
	sram_mem[84249] = 16'b0000000000000000;
	sram_mem[84250] = 16'b0000000000000000;
	sram_mem[84251] = 16'b0000000000000000;
	sram_mem[84252] = 16'b0000000000000000;
	sram_mem[84253] = 16'b0000000000000000;
	sram_mem[84254] = 16'b0000000000000000;
	sram_mem[84255] = 16'b0000000000000000;
	sram_mem[84256] = 16'b0000000000000000;
	sram_mem[84257] = 16'b0000000000000000;
	sram_mem[84258] = 16'b0000000000000000;
	sram_mem[84259] = 16'b0000000000000000;
	sram_mem[84260] = 16'b0000000000000000;
	sram_mem[84261] = 16'b0000000000000000;
	sram_mem[84262] = 16'b0000000000000000;
	sram_mem[84263] = 16'b0000000000000000;
	sram_mem[84264] = 16'b0000000000000000;
	sram_mem[84265] = 16'b0000000000000000;
	sram_mem[84266] = 16'b0000000000000000;
	sram_mem[84267] = 16'b0000000000000000;
	sram_mem[84268] = 16'b0000000000000000;
	sram_mem[84269] = 16'b0000000000000000;
	sram_mem[84270] = 16'b0000000000000000;
	sram_mem[84271] = 16'b0000000000000000;
	sram_mem[84272] = 16'b0000000000000000;
	sram_mem[84273] = 16'b0000000000000000;
	sram_mem[84274] = 16'b0000000000000000;
	sram_mem[84275] = 16'b0000000000000000;
	sram_mem[84276] = 16'b0000000000000000;
	sram_mem[84277] = 16'b0000000000000000;
	sram_mem[84278] = 16'b0000000000000000;
	sram_mem[84279] = 16'b0000000000000000;
	sram_mem[84280] = 16'b0000000000000000;
	sram_mem[84281] = 16'b0000000000000000;
	sram_mem[84282] = 16'b0000000000000000;
	sram_mem[84283] = 16'b0000000000000000;
	sram_mem[84284] = 16'b0000000000000000;
	sram_mem[84285] = 16'b0000000000000000;
	sram_mem[84286] = 16'b0000000000000000;
	sram_mem[84287] = 16'b0000000000000000;
	sram_mem[84288] = 16'b0000000000000000;
	sram_mem[84289] = 16'b0000000000000000;
	sram_mem[84290] = 16'b0000000000000000;
	sram_mem[84291] = 16'b0000000000000000;
	sram_mem[84292] = 16'b0000000000000000;
	sram_mem[84293] = 16'b0000000000000000;
	sram_mem[84294] = 16'b0000000000000000;
	sram_mem[84295] = 16'b0000000000000000;
	sram_mem[84296] = 16'b0000000000000000;
	sram_mem[84297] = 16'b0000000000000000;
	sram_mem[84298] = 16'b0000000000000000;
	sram_mem[84299] = 16'b0000000000000000;
	sram_mem[84300] = 16'b0000000000000000;
	sram_mem[84301] = 16'b0000000000000000;
	sram_mem[84302] = 16'b0000000000000000;
	sram_mem[84303] = 16'b0000000000000000;
	sram_mem[84304] = 16'b0000000000000000;
	sram_mem[84305] = 16'b0000000000000000;
	sram_mem[84306] = 16'b0000000000000000;
	sram_mem[84307] = 16'b0000000000000000;
	sram_mem[84308] = 16'b0000000000000000;
	sram_mem[84309] = 16'b0000000000000000;
	sram_mem[84310] = 16'b0000000000000000;
	sram_mem[84311] = 16'b0000000000000000;
	sram_mem[84312] = 16'b0000000000000000;
	sram_mem[84313] = 16'b0000000000000000;
	sram_mem[84314] = 16'b0000000000000000;
	sram_mem[84315] = 16'b0000000000000000;
	sram_mem[84316] = 16'b0000000000000000;
	sram_mem[84317] = 16'b0000000000000000;
	sram_mem[84318] = 16'b0000000000000000;
	sram_mem[84319] = 16'b0000000000000000;
	sram_mem[84320] = 16'b0000000000000000;
	sram_mem[84321] = 16'b0000000000000000;
	sram_mem[84322] = 16'b0000000000000000;
	sram_mem[84323] = 16'b0000000000000000;
	sram_mem[84324] = 16'b0000000000000000;
	sram_mem[84325] = 16'b0000000000000000;
	sram_mem[84326] = 16'b0000000000000000;
	sram_mem[84327] = 16'b0000000000000000;
	sram_mem[84328] = 16'b0000000000000000;
	sram_mem[84329] = 16'b0000000000000000;
	sram_mem[84330] = 16'b0000000000000000;
	sram_mem[84331] = 16'b0000000000000000;
	sram_mem[84332] = 16'b0000000000000000;
	sram_mem[84333] = 16'b0000000000000000;
	sram_mem[84334] = 16'b0000000000000000;
	sram_mem[84335] = 16'b0000000000000000;
	sram_mem[84336] = 16'b0000000000000000;
	sram_mem[84337] = 16'b0000000000000000;
	sram_mem[84338] = 16'b0000000000000000;
	sram_mem[84339] = 16'b0000000000000000;
	sram_mem[84340] = 16'b0000000000000000;
	sram_mem[84341] = 16'b0000000000000000;
	sram_mem[84342] = 16'b0000000000000000;
	sram_mem[84343] = 16'b0000000000000000;
	sram_mem[84344] = 16'b0000000000000000;
	sram_mem[84345] = 16'b0000000000000000;
	sram_mem[84346] = 16'b0000000000000000;
	sram_mem[84347] = 16'b0000000000000000;
	sram_mem[84348] = 16'b0000000000000000;
	sram_mem[84349] = 16'b0000000000000000;
	sram_mem[84350] = 16'b0000000000000000;
	sram_mem[84351] = 16'b0000000000000000;
	sram_mem[84352] = 16'b0000000000000000;
	sram_mem[84353] = 16'b0000000000000000;
	sram_mem[84354] = 16'b0000000000000000;
	sram_mem[84355] = 16'b0000000000000000;
	sram_mem[84356] = 16'b0000000000000000;
	sram_mem[84357] = 16'b0000000000000000;
	sram_mem[84358] = 16'b0000000000000000;
	sram_mem[84359] = 16'b0000000000000000;
	sram_mem[84360] = 16'b0000000000000000;
	sram_mem[84361] = 16'b0000000000000000;
	sram_mem[84362] = 16'b0000000000000000;
	sram_mem[84363] = 16'b0000000000000000;
	sram_mem[84364] = 16'b0000000000000000;
	sram_mem[84365] = 16'b0000000000000000;
	sram_mem[84366] = 16'b0000000000000000;
	sram_mem[84367] = 16'b0000000000000000;
	sram_mem[84368] = 16'b0000000000000000;
	sram_mem[84369] = 16'b0000000000000000;
	sram_mem[84370] = 16'b0000000000000000;
	sram_mem[84371] = 16'b0000000000000000;
	sram_mem[84372] = 16'b0000000000000000;
	sram_mem[84373] = 16'b0000000000000000;
	sram_mem[84374] = 16'b0000000000000000;
	sram_mem[84375] = 16'b0000000000000000;
	sram_mem[84376] = 16'b0000000000000000;
	sram_mem[84377] = 16'b0000000000000000;
	sram_mem[84378] = 16'b0000000000000000;
	sram_mem[84379] = 16'b0000000000000000;
	sram_mem[84380] = 16'b0000000000000000;
	sram_mem[84381] = 16'b0000000000000000;
	sram_mem[84382] = 16'b0000000000000000;
	sram_mem[84383] = 16'b0000000000000000;
	sram_mem[84384] = 16'b0000000000000000;
	sram_mem[84385] = 16'b0000000000000000;
	sram_mem[84386] = 16'b0000000000000000;
	sram_mem[84387] = 16'b0000000000000000;
	sram_mem[84388] = 16'b0000000000000000;
	sram_mem[84389] = 16'b0000000000000000;
	sram_mem[84390] = 16'b0000000000000000;
	sram_mem[84391] = 16'b0000000000000000;
	sram_mem[84392] = 16'b0000000000000000;
	sram_mem[84393] = 16'b0000000000000000;
	sram_mem[84394] = 16'b0000000000000000;
	sram_mem[84395] = 16'b0000000000000000;
	sram_mem[84396] = 16'b0000000000000000;
	sram_mem[84397] = 16'b0000000000000000;
	sram_mem[84398] = 16'b0000000000000000;
	sram_mem[84399] = 16'b0000000000000000;
	sram_mem[84400] = 16'b0000000000000000;
	sram_mem[84401] = 16'b0000000000000000;
	sram_mem[84402] = 16'b0000000000000000;
	sram_mem[84403] = 16'b0000000000000000;
	sram_mem[84404] = 16'b0000000000000000;
	sram_mem[84405] = 16'b0000000000000000;
	sram_mem[84406] = 16'b0000000000000000;
	sram_mem[84407] = 16'b0000000000000000;
	sram_mem[84408] = 16'b0000000000000000;
	sram_mem[84409] = 16'b0000000000000000;
	sram_mem[84410] = 16'b0000000000000000;
	sram_mem[84411] = 16'b0000000000000000;
	sram_mem[84412] = 16'b0000000000000000;
	sram_mem[84413] = 16'b0000000000000000;
	sram_mem[84414] = 16'b0000000000000000;
	sram_mem[84415] = 16'b0000000000000000;
	sram_mem[84416] = 16'b0000000000000000;
	sram_mem[84417] = 16'b0000000000000000;
	sram_mem[84418] = 16'b0000000000000000;
	sram_mem[84419] = 16'b0000000000000000;
	sram_mem[84420] = 16'b0000000000000000;
	sram_mem[84421] = 16'b0000000000000000;
	sram_mem[84422] = 16'b0000000000000000;
	sram_mem[84423] = 16'b0000000000000000;
	sram_mem[84424] = 16'b0000000000000000;
	sram_mem[84425] = 16'b0000000000000000;
	sram_mem[84426] = 16'b0000000000000000;
	sram_mem[84427] = 16'b0000000000000000;
	sram_mem[84428] = 16'b0000000000000000;
	sram_mem[84429] = 16'b0000000000000000;
	sram_mem[84430] = 16'b0000000000000000;
	sram_mem[84431] = 16'b0000000000000000;
	sram_mem[84432] = 16'b0000000000000000;
	sram_mem[84433] = 16'b0000000000000000;
	sram_mem[84434] = 16'b0000000000000000;
	sram_mem[84435] = 16'b0000000000000000;
	sram_mem[84436] = 16'b0000000000000000;
	sram_mem[84437] = 16'b0000000000000000;
	sram_mem[84438] = 16'b0000000000000000;
	sram_mem[84439] = 16'b0000000000000000;
	sram_mem[84440] = 16'b0000000000000000;
	sram_mem[84441] = 16'b0000000000000000;
	sram_mem[84442] = 16'b0000000000000000;
	sram_mem[84443] = 16'b0000000000000000;
	sram_mem[84444] = 16'b0000000000000000;
	sram_mem[84445] = 16'b0000000000000000;
	sram_mem[84446] = 16'b0000000000000000;
	sram_mem[84447] = 16'b0000000000000000;
	sram_mem[84448] = 16'b0000000000000000;
	sram_mem[84449] = 16'b0000000000000000;
	sram_mem[84450] = 16'b0000000000000000;
	sram_mem[84451] = 16'b0000000000000000;
	sram_mem[84452] = 16'b0000000000000000;
	sram_mem[84453] = 16'b0000000000000000;
	sram_mem[84454] = 16'b0000000000000000;
	sram_mem[84455] = 16'b0000000000000000;
	sram_mem[84456] = 16'b0000000000000000;
	sram_mem[84457] = 16'b0000000000000000;
	sram_mem[84458] = 16'b0000000000000000;
	sram_mem[84459] = 16'b0000000000000000;
	sram_mem[84460] = 16'b0000000000000000;
	sram_mem[84461] = 16'b0000000000000000;
	sram_mem[84462] = 16'b0000000000000000;
	sram_mem[84463] = 16'b0000000000000000;
	sram_mem[84464] = 16'b0000000000000000;
	sram_mem[84465] = 16'b0000000000000000;
	sram_mem[84466] = 16'b0000000000000000;
	sram_mem[84467] = 16'b0000000000000000;
	sram_mem[84468] = 16'b0000000000000000;
	sram_mem[84469] = 16'b0000000000000000;
	sram_mem[84470] = 16'b0000000000000000;
	sram_mem[84471] = 16'b0000000000000000;
	sram_mem[84472] = 16'b0000000000000000;
	sram_mem[84473] = 16'b0000000000000000;
	sram_mem[84474] = 16'b0000000000000000;
	sram_mem[84475] = 16'b0000000000000000;
	sram_mem[84476] = 16'b0000000000000000;
	sram_mem[84477] = 16'b0000000000000000;
	sram_mem[84478] = 16'b0000000000000000;
	sram_mem[84479] = 16'b0000000000000000;
	sram_mem[84480] = 16'b0000000000000000;
	sram_mem[84481] = 16'b0000000000000000;
	sram_mem[84482] = 16'b0000000000000000;
	sram_mem[84483] = 16'b0000000000000000;
	sram_mem[84484] = 16'b0000000000000000;
	sram_mem[84485] = 16'b0000000000000000;
	sram_mem[84486] = 16'b0000000000000000;
	sram_mem[84487] = 16'b0000000000000000;
	sram_mem[84488] = 16'b0000000000000000;
	sram_mem[84489] = 16'b0000000000000000;
	sram_mem[84490] = 16'b0000000000000000;
	sram_mem[84491] = 16'b0000000000000000;
	sram_mem[84492] = 16'b0000000000000000;
	sram_mem[84493] = 16'b0000000000000000;
	sram_mem[84494] = 16'b0000000000000000;
	sram_mem[84495] = 16'b0000000000000000;
	sram_mem[84496] = 16'b0000000000000000;
	sram_mem[84497] = 16'b0000000000000000;
	sram_mem[84498] = 16'b0000000000000000;
	sram_mem[84499] = 16'b0000000000000000;
	sram_mem[84500] = 16'b0000000000000000;
	sram_mem[84501] = 16'b0000000000000000;
	sram_mem[84502] = 16'b0000000000000000;
	sram_mem[84503] = 16'b0000000000000000;
	sram_mem[84504] = 16'b0000000000000000;
	sram_mem[84505] = 16'b0000000000000000;
	sram_mem[84506] = 16'b0000000000000000;
	sram_mem[84507] = 16'b0000000000000000;
	sram_mem[84508] = 16'b0000000000000000;
	sram_mem[84509] = 16'b0000000000000000;
	sram_mem[84510] = 16'b0000000000000000;
	sram_mem[84511] = 16'b0000000000000000;
	sram_mem[84512] = 16'b0000000000000000;
	sram_mem[84513] = 16'b0000000000000000;
	sram_mem[84514] = 16'b0000000000000000;
	sram_mem[84515] = 16'b0000000000000000;
	sram_mem[84516] = 16'b0000000000000000;
	sram_mem[84517] = 16'b0000000000000000;
	sram_mem[84518] = 16'b0000000000000000;
	sram_mem[84519] = 16'b0000000000000000;
	sram_mem[84520] = 16'b0000000000000000;
	sram_mem[84521] = 16'b0000000000000000;
	sram_mem[84522] = 16'b0000000000000000;
	sram_mem[84523] = 16'b0000000000000000;
	sram_mem[84524] = 16'b0000000000000000;
	sram_mem[84525] = 16'b0000000000000000;
	sram_mem[84526] = 16'b0000000000000000;
	sram_mem[84527] = 16'b0000000000000000;
	sram_mem[84528] = 16'b0000000000000000;
	sram_mem[84529] = 16'b0000000000000000;
	sram_mem[84530] = 16'b0000000000000000;
	sram_mem[84531] = 16'b0000000000000000;
	sram_mem[84532] = 16'b0000000000000000;
	sram_mem[84533] = 16'b0000000000000000;
	sram_mem[84534] = 16'b0000000000000000;
	sram_mem[84535] = 16'b0000000000000000;
	sram_mem[84536] = 16'b0000000000000000;
	sram_mem[84537] = 16'b0000000000000000;
	sram_mem[84538] = 16'b0000000000000000;
	sram_mem[84539] = 16'b0000000000000000;
	sram_mem[84540] = 16'b0000000000000000;
	sram_mem[84541] = 16'b0000000000000000;
	sram_mem[84542] = 16'b0000000000000000;
	sram_mem[84543] = 16'b0000000000000000;
	sram_mem[84544] = 16'b0000000000000000;
	sram_mem[84545] = 16'b0000000000000000;
	sram_mem[84546] = 16'b0000000000000000;
	sram_mem[84547] = 16'b0000000000000000;
	sram_mem[84548] = 16'b0000000000000000;
	sram_mem[84549] = 16'b0000000000000000;
	sram_mem[84550] = 16'b0000000000000000;
	sram_mem[84551] = 16'b0000000000000000;
	sram_mem[84552] = 16'b0000000000000000;
	sram_mem[84553] = 16'b0000000000000000;
	sram_mem[84554] = 16'b0000000000000000;
	sram_mem[84555] = 16'b0000000000000000;
	sram_mem[84556] = 16'b0000000000000000;
	sram_mem[84557] = 16'b0000000000000000;
	sram_mem[84558] = 16'b0000000000000000;
	sram_mem[84559] = 16'b0000000000000000;
	sram_mem[84560] = 16'b0000000000000000;
	sram_mem[84561] = 16'b0000000000000000;
	sram_mem[84562] = 16'b0000000000000000;
	sram_mem[84563] = 16'b0000000000000000;
	sram_mem[84564] = 16'b0000000000000000;
	sram_mem[84565] = 16'b0000000000000000;
	sram_mem[84566] = 16'b0000000000000000;
	sram_mem[84567] = 16'b0000000000000000;
	sram_mem[84568] = 16'b0000000000000000;
	sram_mem[84569] = 16'b0000000000000000;
	sram_mem[84570] = 16'b0000000000000000;
	sram_mem[84571] = 16'b0000000000000000;
	sram_mem[84572] = 16'b0000000000000000;
	sram_mem[84573] = 16'b0000000000000000;
	sram_mem[84574] = 16'b0000000000000000;
	sram_mem[84575] = 16'b0000000000000000;
	sram_mem[84576] = 16'b0000000000000000;
	sram_mem[84577] = 16'b0000000000000000;
	sram_mem[84578] = 16'b0000000000000000;
	sram_mem[84579] = 16'b0000000000000000;
	sram_mem[84580] = 16'b0000000000000000;
	sram_mem[84581] = 16'b0000000000000000;
	sram_mem[84582] = 16'b0000000000000000;
	sram_mem[84583] = 16'b0000000000000000;
	sram_mem[84584] = 16'b0000000000000000;
	sram_mem[84585] = 16'b0000000000000000;
	sram_mem[84586] = 16'b0000000000000000;
	sram_mem[84587] = 16'b0000000000000000;
	sram_mem[84588] = 16'b0000000000000000;
	sram_mem[84589] = 16'b0000000000000000;
	sram_mem[84590] = 16'b0000000000000000;
	sram_mem[84591] = 16'b0000000000000000;
	sram_mem[84592] = 16'b0000000000000000;
	sram_mem[84593] = 16'b0000000000000000;
	sram_mem[84594] = 16'b0000000000000000;
	sram_mem[84595] = 16'b0000000000000000;
	sram_mem[84596] = 16'b0000000000000000;
	sram_mem[84597] = 16'b0000000000000000;
	sram_mem[84598] = 16'b0000000000000000;
	sram_mem[84599] = 16'b0000000000000000;
	sram_mem[84600] = 16'b0000000000000000;
	sram_mem[84601] = 16'b0000000000000000;
	sram_mem[84602] = 16'b0000000000000000;
	sram_mem[84603] = 16'b0000000000000000;
	sram_mem[84604] = 16'b0000000000000000;
	sram_mem[84605] = 16'b0000000000000000;
	sram_mem[84606] = 16'b0000000000000000;
	sram_mem[84607] = 16'b0000000000000000;
	sram_mem[84608] = 16'b0000000000000000;
	sram_mem[84609] = 16'b0000000000000000;
	sram_mem[84610] = 16'b0000000000000000;
	sram_mem[84611] = 16'b0000000000000000;
	sram_mem[84612] = 16'b0000000000000000;
	sram_mem[84613] = 16'b0000000000000000;
	sram_mem[84614] = 16'b0000000000000000;
	sram_mem[84615] = 16'b0000000000000000;
	sram_mem[84616] = 16'b0000000000000000;
	sram_mem[84617] = 16'b0000000000000000;
	sram_mem[84618] = 16'b0000000000000000;
	sram_mem[84619] = 16'b0000000000000000;
	sram_mem[84620] = 16'b0000000000000000;
	sram_mem[84621] = 16'b0000000000000000;
	sram_mem[84622] = 16'b0000000000000000;
	sram_mem[84623] = 16'b0000000000000000;
	sram_mem[84624] = 16'b0000000000000000;
	sram_mem[84625] = 16'b0000000000000000;
	sram_mem[84626] = 16'b0000000000000000;
	sram_mem[84627] = 16'b0000000000000000;
	sram_mem[84628] = 16'b0000000000000000;
	sram_mem[84629] = 16'b0000000000000000;
	sram_mem[84630] = 16'b0000000000000000;
	sram_mem[84631] = 16'b0000000000000000;
	sram_mem[84632] = 16'b0000000000000000;
	sram_mem[84633] = 16'b0000000000000000;
	sram_mem[84634] = 16'b0000000000000000;
	sram_mem[84635] = 16'b0000000000000000;
	sram_mem[84636] = 16'b0000000000000000;
	sram_mem[84637] = 16'b0000000000000000;
	sram_mem[84638] = 16'b0000000000000000;
	sram_mem[84639] = 16'b0000000000000000;
	sram_mem[84640] = 16'b0000000000000000;
	sram_mem[84641] = 16'b0000000000000000;
	sram_mem[84642] = 16'b0000000000000000;
	sram_mem[84643] = 16'b0000000000000000;
	sram_mem[84644] = 16'b0000000000000000;
	sram_mem[84645] = 16'b0000000000000000;
	sram_mem[84646] = 16'b0000000000000000;
	sram_mem[84647] = 16'b0000000000000000;
	sram_mem[84648] = 16'b0000000000000000;
	sram_mem[84649] = 16'b0000000000000000;
	sram_mem[84650] = 16'b0000000000000000;
	sram_mem[84651] = 16'b0000000000000000;
	sram_mem[84652] = 16'b0000000000000000;
	sram_mem[84653] = 16'b0000000000000000;
	sram_mem[84654] = 16'b0000000000000000;
	sram_mem[84655] = 16'b0000000000000000;
	sram_mem[84656] = 16'b0000000000000000;
	sram_mem[84657] = 16'b0000000000000000;
	sram_mem[84658] = 16'b0000000000000000;
	sram_mem[84659] = 16'b0000000000000000;
	sram_mem[84660] = 16'b0000000000000000;
	sram_mem[84661] = 16'b0000000000000000;
	sram_mem[84662] = 16'b0000000000000000;
	sram_mem[84663] = 16'b0000000000000000;
	sram_mem[84664] = 16'b0000000000000000;
	sram_mem[84665] = 16'b0000000000000000;
	sram_mem[84666] = 16'b0000000000000000;
	sram_mem[84667] = 16'b0000000000000000;
	sram_mem[84668] = 16'b0000000000000000;
	sram_mem[84669] = 16'b0000000000000000;
	sram_mem[84670] = 16'b0000000000000000;
	sram_mem[84671] = 16'b0000000000000000;
	sram_mem[84672] = 16'b0000000000000000;
	sram_mem[84673] = 16'b0000000000000000;
	sram_mem[84674] = 16'b0000000000000000;
	sram_mem[84675] = 16'b0000000000000000;
	sram_mem[84676] = 16'b0000000000000000;
	sram_mem[84677] = 16'b0000000000000000;
	sram_mem[84678] = 16'b0000000000000000;
	sram_mem[84679] = 16'b0000000000000000;
	sram_mem[84680] = 16'b0000000000000000;
	sram_mem[84681] = 16'b0000000000000000;
	sram_mem[84682] = 16'b0000000000000000;
	sram_mem[84683] = 16'b0000000000000000;
	sram_mem[84684] = 16'b0000000000000000;
	sram_mem[84685] = 16'b0000000000000000;
	sram_mem[84686] = 16'b0000000000000000;
	sram_mem[84687] = 16'b0000000000000000;
	sram_mem[84688] = 16'b0000000000000000;
	sram_mem[84689] = 16'b0000000000000000;
	sram_mem[84690] = 16'b0000000000000000;
	sram_mem[84691] = 16'b0000000000000000;
	sram_mem[84692] = 16'b0000000000000000;
	sram_mem[84693] = 16'b0000000000000000;
	sram_mem[84694] = 16'b0000000000000000;
	sram_mem[84695] = 16'b0000000000000000;
	sram_mem[84696] = 16'b0000000000000000;
	sram_mem[84697] = 16'b0000000000000000;
	sram_mem[84698] = 16'b0000000000000000;
	sram_mem[84699] = 16'b0000000000000000;
	sram_mem[84700] = 16'b0000000000000000;
	sram_mem[84701] = 16'b0000000000000000;
	sram_mem[84702] = 16'b0000000000000000;
	sram_mem[84703] = 16'b0000000000000000;
	sram_mem[84704] = 16'b0000000000000000;
	sram_mem[84705] = 16'b0000000000000000;
	sram_mem[84706] = 16'b0000000000000000;
	sram_mem[84707] = 16'b0000000000000000;
	sram_mem[84708] = 16'b0000000000000000;
	sram_mem[84709] = 16'b0000000000000000;
	sram_mem[84710] = 16'b0000000000000000;
	sram_mem[84711] = 16'b0000000000000000;
	sram_mem[84712] = 16'b0000000000000000;
	sram_mem[84713] = 16'b0000000000000000;
	sram_mem[84714] = 16'b0000000000000000;
	sram_mem[84715] = 16'b0000000000000000;
	sram_mem[84716] = 16'b0000000000000000;
	sram_mem[84717] = 16'b0000000000000000;
	sram_mem[84718] = 16'b0000000000000000;
	sram_mem[84719] = 16'b0000000000000000;
	sram_mem[84720] = 16'b0000000000000000;
	sram_mem[84721] = 16'b0000000000000000;
	sram_mem[84722] = 16'b0000000000000000;
	sram_mem[84723] = 16'b0000000000000000;
	sram_mem[84724] = 16'b0000000000000000;
	sram_mem[84725] = 16'b0000000000000000;
	sram_mem[84726] = 16'b0000000000000000;
	sram_mem[84727] = 16'b0000000000000000;
	sram_mem[84728] = 16'b0000000000000000;
	sram_mem[84729] = 16'b0000000000000000;
	sram_mem[84730] = 16'b0000000000000000;
	sram_mem[84731] = 16'b0000000000000000;
	sram_mem[84732] = 16'b0000000000000000;
	sram_mem[84733] = 16'b0000000000000000;
	sram_mem[84734] = 16'b0000000000000000;
	sram_mem[84735] = 16'b0000000000000000;
	sram_mem[84736] = 16'b0000000000000000;
	sram_mem[84737] = 16'b0000000000000000;
	sram_mem[84738] = 16'b0000000000000000;
	sram_mem[84739] = 16'b0000000000000000;
	sram_mem[84740] = 16'b0000000000000000;
	sram_mem[84741] = 16'b0000000000000000;
	sram_mem[84742] = 16'b0000000000000000;
	sram_mem[84743] = 16'b0000000000000000;
	sram_mem[84744] = 16'b0000000000000000;
	sram_mem[84745] = 16'b0000000000000000;
	sram_mem[84746] = 16'b0000000000000000;
	sram_mem[84747] = 16'b0000000000000000;
	sram_mem[84748] = 16'b0000000000000000;
	sram_mem[84749] = 16'b0000000000000000;
	sram_mem[84750] = 16'b0000000000000000;
	sram_mem[84751] = 16'b0000000000000000;
	sram_mem[84752] = 16'b0000000000000000;
	sram_mem[84753] = 16'b0000000000000000;
	sram_mem[84754] = 16'b0000000000000000;
	sram_mem[84755] = 16'b0000000000000000;
	sram_mem[84756] = 16'b0000000000000000;
	sram_mem[84757] = 16'b0000000000000000;
	sram_mem[84758] = 16'b0000000000000000;
	sram_mem[84759] = 16'b0000000000000000;
	sram_mem[84760] = 16'b0000000000000000;
	sram_mem[84761] = 16'b0000000000000000;
	sram_mem[84762] = 16'b0000000000000000;
	sram_mem[84763] = 16'b0000000000000000;
	sram_mem[84764] = 16'b0000000000000000;
	sram_mem[84765] = 16'b0000000000000000;
	sram_mem[84766] = 16'b0000000000000000;
	sram_mem[84767] = 16'b0000000000000000;
	sram_mem[84768] = 16'b0000000000000000;
	sram_mem[84769] = 16'b0000000000000000;
	sram_mem[84770] = 16'b0000000000000000;
	sram_mem[84771] = 16'b0000000000000000;
	sram_mem[84772] = 16'b0000000000000000;
	sram_mem[84773] = 16'b0000000000000000;
	sram_mem[84774] = 16'b0000000000000000;
	sram_mem[84775] = 16'b0000000000000000;
	sram_mem[84776] = 16'b0000000000000000;
	sram_mem[84777] = 16'b0000000000000000;
	sram_mem[84778] = 16'b0000000000000000;
	sram_mem[84779] = 16'b0000000000000000;
	sram_mem[84780] = 16'b0000000000000000;
	sram_mem[84781] = 16'b0000000000000000;
	sram_mem[84782] = 16'b0000000000000000;
	sram_mem[84783] = 16'b0000000000000000;
	sram_mem[84784] = 16'b0000000000000000;
	sram_mem[84785] = 16'b0000000000000000;
	sram_mem[84786] = 16'b0000000000000000;
	sram_mem[84787] = 16'b0000000000000000;
	sram_mem[84788] = 16'b0000000000000000;
	sram_mem[84789] = 16'b0000000000000000;
	sram_mem[84790] = 16'b0000000000000000;
	sram_mem[84791] = 16'b0000000000000000;
	sram_mem[84792] = 16'b0000000000000000;
	sram_mem[84793] = 16'b0000000000000000;
	sram_mem[84794] = 16'b0000000000000000;
	sram_mem[84795] = 16'b0000000000000000;
	sram_mem[84796] = 16'b0000000000000000;
	sram_mem[84797] = 16'b0000000000000000;
	sram_mem[84798] = 16'b0000000000000000;
	sram_mem[84799] = 16'b0000000000000000;
	sram_mem[84800] = 16'b0000000000000000;
	sram_mem[84801] = 16'b0000000000000000;
	sram_mem[84802] = 16'b0000000000000000;
	sram_mem[84803] = 16'b0000000000000000;
	sram_mem[84804] = 16'b0000000000000000;
	sram_mem[84805] = 16'b0000000000000000;
	sram_mem[84806] = 16'b0000000000000000;
	sram_mem[84807] = 16'b0000000000000000;
	sram_mem[84808] = 16'b0000000000000000;
	sram_mem[84809] = 16'b0000000000000000;
	sram_mem[84810] = 16'b0000000000000000;
	sram_mem[84811] = 16'b0000000000000000;
	sram_mem[84812] = 16'b0000000000000000;
	sram_mem[84813] = 16'b0000000000000000;
	sram_mem[84814] = 16'b0000000000000000;
	sram_mem[84815] = 16'b0000000000000000;
	sram_mem[84816] = 16'b0000000000000000;
	sram_mem[84817] = 16'b0000000000000000;
	sram_mem[84818] = 16'b0000000000000000;
	sram_mem[84819] = 16'b0000000000000000;
	sram_mem[84820] = 16'b0000000000000000;
	sram_mem[84821] = 16'b0000000000000000;
	sram_mem[84822] = 16'b0000000000000000;
	sram_mem[84823] = 16'b0000000000000000;
	sram_mem[84824] = 16'b0000000000000000;
	sram_mem[84825] = 16'b0000000000000000;
	sram_mem[84826] = 16'b0000000000000000;
	sram_mem[84827] = 16'b0000000000000000;
	sram_mem[84828] = 16'b0000000000000000;
	sram_mem[84829] = 16'b0000000000000000;
	sram_mem[84830] = 16'b0000000000000000;
	sram_mem[84831] = 16'b0000000000000000;
	sram_mem[84832] = 16'b0000000000000000;
	sram_mem[84833] = 16'b0000000000000000;
	sram_mem[84834] = 16'b0000000000000000;
	sram_mem[84835] = 16'b0000000000000000;
	sram_mem[84836] = 16'b0000000000000000;
	sram_mem[84837] = 16'b0000000000000000;
	sram_mem[84838] = 16'b0000000000000000;
	sram_mem[84839] = 16'b0000000000000000;
	sram_mem[84840] = 16'b0000000000000000;
	sram_mem[84841] = 16'b0000000000000000;
	sram_mem[84842] = 16'b0000000000000000;
	sram_mem[84843] = 16'b0000000000000000;
	sram_mem[84844] = 16'b0000000000000000;
	sram_mem[84845] = 16'b0000000000000000;
	sram_mem[84846] = 16'b0000000000000000;
	sram_mem[84847] = 16'b0000000000000000;
	sram_mem[84848] = 16'b0000000000000000;
	sram_mem[84849] = 16'b0000000000000000;
	sram_mem[84850] = 16'b0000000000000000;
	sram_mem[84851] = 16'b0000000000000000;
	sram_mem[84852] = 16'b0000000000000000;
	sram_mem[84853] = 16'b0000000000000000;
	sram_mem[84854] = 16'b0000000000000000;
	sram_mem[84855] = 16'b0000000000000000;
	sram_mem[84856] = 16'b0000000000000000;
	sram_mem[84857] = 16'b0000000000000000;
	sram_mem[84858] = 16'b0000000000000000;
	sram_mem[84859] = 16'b0000000000000000;
	sram_mem[84860] = 16'b0000000000000000;
	sram_mem[84861] = 16'b0000000000000000;
	sram_mem[84862] = 16'b0000000000000000;
	sram_mem[84863] = 16'b0000000000000000;
	sram_mem[84864] = 16'b0000000000000000;
	sram_mem[84865] = 16'b0000000000000000;
	sram_mem[84866] = 16'b0000000000000000;
	sram_mem[84867] = 16'b0000000000000000;
	sram_mem[84868] = 16'b0000000000000000;
	sram_mem[84869] = 16'b0000000000000000;
	sram_mem[84870] = 16'b0000000000000000;
	sram_mem[84871] = 16'b0000000000000000;
	sram_mem[84872] = 16'b0000000000000000;
	sram_mem[84873] = 16'b0000000000000000;
	sram_mem[84874] = 16'b0000000000000000;
	sram_mem[84875] = 16'b0000000000000000;
	sram_mem[84876] = 16'b0000000000000000;
	sram_mem[84877] = 16'b0000000000000000;
	sram_mem[84878] = 16'b0000000000000000;
	sram_mem[84879] = 16'b0000000000000000;
	sram_mem[84880] = 16'b0000000000000000;
	sram_mem[84881] = 16'b0000000000000000;
	sram_mem[84882] = 16'b0000000000000000;
	sram_mem[84883] = 16'b0000000000000000;
	sram_mem[84884] = 16'b0000000000000000;
	sram_mem[84885] = 16'b0000000000000000;
	sram_mem[84886] = 16'b0000000000000000;
	sram_mem[84887] = 16'b0000000000000000;
	sram_mem[84888] = 16'b0000000000000000;
	sram_mem[84889] = 16'b0000000000000000;
	sram_mem[84890] = 16'b0000000000000000;
	sram_mem[84891] = 16'b0000000000000000;
	sram_mem[84892] = 16'b0000000000000000;
	sram_mem[84893] = 16'b0000000000000000;
	sram_mem[84894] = 16'b0000000000000000;
	sram_mem[84895] = 16'b0000000000000000;
	sram_mem[84896] = 16'b0000000000000000;
	sram_mem[84897] = 16'b0000000000000000;
	sram_mem[84898] = 16'b0000000000000000;
	sram_mem[84899] = 16'b0000000000000000;
	sram_mem[84900] = 16'b0000000000000000;
	sram_mem[84901] = 16'b0000000000000000;
	sram_mem[84902] = 16'b0000000000000000;
	sram_mem[84903] = 16'b0000000000000000;
	sram_mem[84904] = 16'b0000000000000000;
	sram_mem[84905] = 16'b0000000000000000;
	sram_mem[84906] = 16'b0000000000000000;
	sram_mem[84907] = 16'b0000000000000000;
	sram_mem[84908] = 16'b0000000000000000;
	sram_mem[84909] = 16'b0000000000000000;
	sram_mem[84910] = 16'b0000000000000000;
	sram_mem[84911] = 16'b0000000000000000;
	sram_mem[84912] = 16'b0000000000000000;
	sram_mem[84913] = 16'b0000000000000000;
	sram_mem[84914] = 16'b0000000000000000;
	sram_mem[84915] = 16'b0000000000000000;
	sram_mem[84916] = 16'b0000000000000000;
	sram_mem[84917] = 16'b0000000000000000;
	sram_mem[84918] = 16'b0000000000000000;
	sram_mem[84919] = 16'b0000000000000000;
	sram_mem[84920] = 16'b0000000000000000;
	sram_mem[84921] = 16'b0000000000000000;
	sram_mem[84922] = 16'b0000000000000000;
	sram_mem[84923] = 16'b0000000000000000;
	sram_mem[84924] = 16'b0000000000000000;
	sram_mem[84925] = 16'b0000000000000000;
	sram_mem[84926] = 16'b0000000000000000;
	sram_mem[84927] = 16'b0000000000000000;
	sram_mem[84928] = 16'b0000000000000000;
	sram_mem[84929] = 16'b0000000000000000;
	sram_mem[84930] = 16'b0000000000000000;
	sram_mem[84931] = 16'b0000000000000000;
	sram_mem[84932] = 16'b0000000000000000;
	sram_mem[84933] = 16'b0000000000000000;
	sram_mem[84934] = 16'b0000000000000000;
	sram_mem[84935] = 16'b0000000000000000;
	sram_mem[84936] = 16'b0000000000000000;
	sram_mem[84937] = 16'b0000000000000000;
	sram_mem[84938] = 16'b0000000000000000;
	sram_mem[84939] = 16'b0000000000000000;
	sram_mem[84940] = 16'b0000000000000000;
	sram_mem[84941] = 16'b0000000000000000;
	sram_mem[84942] = 16'b0000000000000000;
	sram_mem[84943] = 16'b0000000000000000;
	sram_mem[84944] = 16'b0000000000000000;
	sram_mem[84945] = 16'b0000000000000000;
	sram_mem[84946] = 16'b0000000000000000;
	sram_mem[84947] = 16'b0000000000000000;
	sram_mem[84948] = 16'b0000000000000000;
	sram_mem[84949] = 16'b0000000000000000;
	sram_mem[84950] = 16'b0000000000000000;
	sram_mem[84951] = 16'b0000000000000000;
	sram_mem[84952] = 16'b0000000000000000;
	sram_mem[84953] = 16'b0000000000000000;
	sram_mem[84954] = 16'b0000000000000000;
	sram_mem[84955] = 16'b0000000000000000;
	sram_mem[84956] = 16'b0000000000000000;
	sram_mem[84957] = 16'b0000000000000000;
	sram_mem[84958] = 16'b0000000000000000;
	sram_mem[84959] = 16'b0000000000000000;
	sram_mem[84960] = 16'b0000000000000000;
	sram_mem[84961] = 16'b0000000000000000;
	sram_mem[84962] = 16'b0000000000000000;
	sram_mem[84963] = 16'b0000000000000000;
	sram_mem[84964] = 16'b0000000000000000;
	sram_mem[84965] = 16'b0000000000000000;
	sram_mem[84966] = 16'b0000000000000000;
	sram_mem[84967] = 16'b0000000000000000;
	sram_mem[84968] = 16'b0000000000000000;
	sram_mem[84969] = 16'b0000000000000000;
	sram_mem[84970] = 16'b0000000000000000;
	sram_mem[84971] = 16'b0000000000000000;
	sram_mem[84972] = 16'b0000000000000000;
	sram_mem[84973] = 16'b0000000000000000;
	sram_mem[84974] = 16'b0000000000000000;
	sram_mem[84975] = 16'b0000000000000000;
	sram_mem[84976] = 16'b0000000000000000;
	sram_mem[84977] = 16'b0000000000000000;
	sram_mem[84978] = 16'b0000000000000000;
	sram_mem[84979] = 16'b0000000000000000;
	sram_mem[84980] = 16'b0000000000000000;
	sram_mem[84981] = 16'b0000000000000000;
	sram_mem[84982] = 16'b0000000000000000;
	sram_mem[84983] = 16'b0000000000000000;
	sram_mem[84984] = 16'b0000000000000000;
	sram_mem[84985] = 16'b0000000000000000;
	sram_mem[84986] = 16'b0000000000000000;
	sram_mem[84987] = 16'b0000000000000000;
	sram_mem[84988] = 16'b0000000000000000;
	sram_mem[84989] = 16'b0000000000000000;
	sram_mem[84990] = 16'b0000000000000000;
	sram_mem[84991] = 16'b0000000000000000;
	sram_mem[84992] = 16'b0000000000000000;
	sram_mem[84993] = 16'b0000000000000000;
	sram_mem[84994] = 16'b0000000000000000;
	sram_mem[84995] = 16'b0000000000000000;
	sram_mem[84996] = 16'b0000000000000000;
	sram_mem[84997] = 16'b0000000000000000;
	sram_mem[84998] = 16'b0000000000000000;
	sram_mem[84999] = 16'b0000000000000000;
	sram_mem[85000] = 16'b0000000000000000;
	sram_mem[85001] = 16'b0000000000000000;
	sram_mem[85002] = 16'b0000000000000000;
	sram_mem[85003] = 16'b0000000000000000;
	sram_mem[85004] = 16'b0000000000000000;
	sram_mem[85005] = 16'b0000000000000000;
	sram_mem[85006] = 16'b0000000000000000;
	sram_mem[85007] = 16'b0000000000000000;
	sram_mem[85008] = 16'b0000000000000000;
	sram_mem[85009] = 16'b0000000000000000;
	sram_mem[85010] = 16'b0000000000000000;
	sram_mem[85011] = 16'b0000000000000000;
	sram_mem[85012] = 16'b0000000000000000;
	sram_mem[85013] = 16'b0000000000000000;
	sram_mem[85014] = 16'b0000000000000000;
	sram_mem[85015] = 16'b0000000000000000;
	sram_mem[85016] = 16'b0000000000000000;
	sram_mem[85017] = 16'b0000000000000000;
	sram_mem[85018] = 16'b0000000000000000;
	sram_mem[85019] = 16'b0000000000000000;
	sram_mem[85020] = 16'b0000000000000000;
	sram_mem[85021] = 16'b0000000000000000;
	sram_mem[85022] = 16'b0000000000000000;
	sram_mem[85023] = 16'b0000000000000000;
	sram_mem[85024] = 16'b0000000000000000;
	sram_mem[85025] = 16'b0000000000000000;
	sram_mem[85026] = 16'b0000000000000000;
	sram_mem[85027] = 16'b0000000000000000;
	sram_mem[85028] = 16'b0000000000000000;
	sram_mem[85029] = 16'b0000000000000000;
	sram_mem[85030] = 16'b0000000000000000;
	sram_mem[85031] = 16'b0000000000000000;
	sram_mem[85032] = 16'b0000000000000000;
	sram_mem[85033] = 16'b0000000000000000;
	sram_mem[85034] = 16'b0000000000000000;
	sram_mem[85035] = 16'b0000000000000000;
	sram_mem[85036] = 16'b0000000000000000;
	sram_mem[85037] = 16'b0000000000000000;
	sram_mem[85038] = 16'b0000000000000000;
	sram_mem[85039] = 16'b0000000000000000;
	sram_mem[85040] = 16'b0000000000000000;
	sram_mem[85041] = 16'b0000000000000000;
	sram_mem[85042] = 16'b0000000000000000;
	sram_mem[85043] = 16'b0000000000000000;
	sram_mem[85044] = 16'b0000000000000000;
	sram_mem[85045] = 16'b0000000000000000;
	sram_mem[85046] = 16'b0000000000000000;
	sram_mem[85047] = 16'b0000000000000000;
	sram_mem[85048] = 16'b0000000000000000;
	sram_mem[85049] = 16'b0000000000000000;
	sram_mem[85050] = 16'b0000000000000000;
	sram_mem[85051] = 16'b0000000000000000;
	sram_mem[85052] = 16'b0000000000000000;
	sram_mem[85053] = 16'b0000000000000000;
	sram_mem[85054] = 16'b0000000000000000;
	sram_mem[85055] = 16'b0000000000000000;
	sram_mem[85056] = 16'b0000000000000000;
	sram_mem[85057] = 16'b0000000000000000;
	sram_mem[85058] = 16'b0000000000000000;
	sram_mem[85059] = 16'b0000000000000000;
	sram_mem[85060] = 16'b0000000000000000;
	sram_mem[85061] = 16'b0000000000000000;
	sram_mem[85062] = 16'b0000000000000000;
	sram_mem[85063] = 16'b0000000000000000;
	sram_mem[85064] = 16'b0000000000000000;
	sram_mem[85065] = 16'b0000000000000000;
	sram_mem[85066] = 16'b0000000000000000;
	sram_mem[85067] = 16'b0000000000000000;
	sram_mem[85068] = 16'b0000000000000000;
	sram_mem[85069] = 16'b0000000000000000;
	sram_mem[85070] = 16'b0000000000000000;
	sram_mem[85071] = 16'b0000000000000000;
	sram_mem[85072] = 16'b0000000000000000;
	sram_mem[85073] = 16'b0000000000000000;
	sram_mem[85074] = 16'b0000000000000000;
	sram_mem[85075] = 16'b0000000000000000;
	sram_mem[85076] = 16'b0000000000000000;
	sram_mem[85077] = 16'b0000000000000000;
	sram_mem[85078] = 16'b0000000000000000;
	sram_mem[85079] = 16'b0000000000000000;
	sram_mem[85080] = 16'b0000000000000000;
	sram_mem[85081] = 16'b0000000000000000;
	sram_mem[85082] = 16'b0000000000000000;
	sram_mem[85083] = 16'b0000000000000000;
	sram_mem[85084] = 16'b0000000000000000;
	sram_mem[85085] = 16'b0000000000000000;
	sram_mem[85086] = 16'b0000000000000000;
	sram_mem[85087] = 16'b0000000000000000;
	sram_mem[85088] = 16'b0000000000000000;
	sram_mem[85089] = 16'b0000000000000000;
	sram_mem[85090] = 16'b0000000000000000;
	sram_mem[85091] = 16'b0000000000000000;
	sram_mem[85092] = 16'b0000000000000000;
	sram_mem[85093] = 16'b0000000000000000;
	sram_mem[85094] = 16'b0000000000000000;
	sram_mem[85095] = 16'b0000000000000000;
	sram_mem[85096] = 16'b0000000000000000;
	sram_mem[85097] = 16'b0000000000000000;
	sram_mem[85098] = 16'b0000000000000000;
	sram_mem[85099] = 16'b0000000000000000;
	sram_mem[85100] = 16'b0000000000000000;
	sram_mem[85101] = 16'b0000000000000000;
	sram_mem[85102] = 16'b0000000000000000;
	sram_mem[85103] = 16'b0000000000000000;
	sram_mem[85104] = 16'b0000000000000000;
	sram_mem[85105] = 16'b0000000000000000;
	sram_mem[85106] = 16'b0000000000000000;
	sram_mem[85107] = 16'b0000000000000000;
	sram_mem[85108] = 16'b0000000000000000;
	sram_mem[85109] = 16'b0000000000000000;
	sram_mem[85110] = 16'b0000000000000000;
	sram_mem[85111] = 16'b0000000000000000;
	sram_mem[85112] = 16'b0000000000000000;
	sram_mem[85113] = 16'b0000000000000000;
	sram_mem[85114] = 16'b0000000000000000;
	sram_mem[85115] = 16'b0000000000000000;
	sram_mem[85116] = 16'b0000000000000000;
	sram_mem[85117] = 16'b0000000000000000;
	sram_mem[85118] = 16'b0000000000000000;
	sram_mem[85119] = 16'b0000000000000000;
	sram_mem[85120] = 16'b0000000000000000;
	sram_mem[85121] = 16'b0000000000000000;
	sram_mem[85122] = 16'b0000000000000000;
	sram_mem[85123] = 16'b0000000000000000;
	sram_mem[85124] = 16'b0000000000000000;
	sram_mem[85125] = 16'b0000000000000000;
	sram_mem[85126] = 16'b0000000000000000;
	sram_mem[85127] = 16'b0000000000000000;
	sram_mem[85128] = 16'b0000000000000000;
	sram_mem[85129] = 16'b0000000000000000;
	sram_mem[85130] = 16'b0000000000000000;
	sram_mem[85131] = 16'b0000000000000000;
	sram_mem[85132] = 16'b0000000000000000;
	sram_mem[85133] = 16'b0000000000000000;
	sram_mem[85134] = 16'b0000000000000000;
	sram_mem[85135] = 16'b0000000000000000;
	sram_mem[85136] = 16'b0000000000000000;
	sram_mem[85137] = 16'b0000000000000000;
	sram_mem[85138] = 16'b0000000000000000;
	sram_mem[85139] = 16'b0000000000000000;
	sram_mem[85140] = 16'b0000000000000000;
	sram_mem[85141] = 16'b0000000000000000;
	sram_mem[85142] = 16'b0000000000000000;
	sram_mem[85143] = 16'b0000000000000000;
	sram_mem[85144] = 16'b0000000000000000;
	sram_mem[85145] = 16'b0000000000000000;
	sram_mem[85146] = 16'b0000000000000000;
	sram_mem[85147] = 16'b0000000000000000;
	sram_mem[85148] = 16'b0000000000000000;
	sram_mem[85149] = 16'b0000000000000000;
	sram_mem[85150] = 16'b0000000000000000;
	sram_mem[85151] = 16'b0000000000000000;
	sram_mem[85152] = 16'b0000000000000000;
	sram_mem[85153] = 16'b0000000000000000;
	sram_mem[85154] = 16'b0000000000000000;
	sram_mem[85155] = 16'b0000000000000000;
	sram_mem[85156] = 16'b0000000000000000;
	sram_mem[85157] = 16'b0000000000000000;
	sram_mem[85158] = 16'b0000000000000000;
	sram_mem[85159] = 16'b0000000000000000;
	sram_mem[85160] = 16'b0000000000000000;
	sram_mem[85161] = 16'b0000000000000000;
	sram_mem[85162] = 16'b0000000000000000;
	sram_mem[85163] = 16'b0000000000000000;
	sram_mem[85164] = 16'b0000000000000000;
	sram_mem[85165] = 16'b0000000000000000;
	sram_mem[85166] = 16'b0000000000000000;
	sram_mem[85167] = 16'b0000000000000000;
	sram_mem[85168] = 16'b0000000000000000;
	sram_mem[85169] = 16'b0000000000000000;
	sram_mem[85170] = 16'b0000000000000000;
	sram_mem[85171] = 16'b0000000000000000;
	sram_mem[85172] = 16'b0000000000000000;
	sram_mem[85173] = 16'b0000000000000000;
	sram_mem[85174] = 16'b0000000000000000;
	sram_mem[85175] = 16'b0000000000000000;
	sram_mem[85176] = 16'b0000000000000000;
	sram_mem[85177] = 16'b0000000000000000;
	sram_mem[85178] = 16'b0000000000000000;
	sram_mem[85179] = 16'b0000000000000000;
	sram_mem[85180] = 16'b0000000000000000;
	sram_mem[85181] = 16'b0000000000000000;
	sram_mem[85182] = 16'b0000000000000000;
	sram_mem[85183] = 16'b0000000000000000;
	sram_mem[85184] = 16'b0000000000000000;
	sram_mem[85185] = 16'b0000000000000000;
	sram_mem[85186] = 16'b0000000000000000;
	sram_mem[85187] = 16'b0000000000000000;
	sram_mem[85188] = 16'b0000000000000000;
	sram_mem[85189] = 16'b0000000000000000;
	sram_mem[85190] = 16'b0000000000000000;
	sram_mem[85191] = 16'b0000000000000000;
	sram_mem[85192] = 16'b0000000000000000;
	sram_mem[85193] = 16'b0000000000000000;
	sram_mem[85194] = 16'b0000000000000000;
	sram_mem[85195] = 16'b0000000000000000;
	sram_mem[85196] = 16'b0000000000000000;
	sram_mem[85197] = 16'b0000000000000000;
	sram_mem[85198] = 16'b0000000000000000;
	sram_mem[85199] = 16'b0000000000000000;
	sram_mem[85200] = 16'b0000000000000000;
	sram_mem[85201] = 16'b0000000000000000;
	sram_mem[85202] = 16'b0000000000000000;
	sram_mem[85203] = 16'b0000000000000000;
	sram_mem[85204] = 16'b0000000000000000;
	sram_mem[85205] = 16'b0000000000000000;
	sram_mem[85206] = 16'b0000000000000000;
	sram_mem[85207] = 16'b0000000000000000;
	sram_mem[85208] = 16'b0000000000000000;
	sram_mem[85209] = 16'b0000000000000000;
	sram_mem[85210] = 16'b0000000000000000;
	sram_mem[85211] = 16'b0000000000000000;
	sram_mem[85212] = 16'b0000000000000000;
	sram_mem[85213] = 16'b0000000000000000;
	sram_mem[85214] = 16'b0000000000000000;
	sram_mem[85215] = 16'b0000000000000000;
	sram_mem[85216] = 16'b0000000000000000;
	sram_mem[85217] = 16'b0000000000000000;
	sram_mem[85218] = 16'b0000000000000000;
	sram_mem[85219] = 16'b0000000000000000;
	sram_mem[85220] = 16'b0000000000000000;
	sram_mem[85221] = 16'b0000000000000000;
	sram_mem[85222] = 16'b0000000000000000;
	sram_mem[85223] = 16'b0000000000000000;
	sram_mem[85224] = 16'b0000000000000000;
	sram_mem[85225] = 16'b0000000000000000;
	sram_mem[85226] = 16'b0000000000000000;
	sram_mem[85227] = 16'b0000000000000000;
	sram_mem[85228] = 16'b0000000000000000;
	sram_mem[85229] = 16'b0000000000000000;
	sram_mem[85230] = 16'b0000000000000000;
	sram_mem[85231] = 16'b0000000000000000;
	sram_mem[85232] = 16'b0000000000000000;
	sram_mem[85233] = 16'b0000000000000000;
	sram_mem[85234] = 16'b0000000000000000;
	sram_mem[85235] = 16'b0000000000000000;
	sram_mem[85236] = 16'b0000000000000000;
	sram_mem[85237] = 16'b0000000000000000;
	sram_mem[85238] = 16'b0000000000000000;
	sram_mem[85239] = 16'b0000000000000000;
	sram_mem[85240] = 16'b0000000000000000;
	sram_mem[85241] = 16'b0000000000000000;
	sram_mem[85242] = 16'b0000000000000000;
	sram_mem[85243] = 16'b0000000000000000;
	sram_mem[85244] = 16'b0000000000000000;
	sram_mem[85245] = 16'b0000000000000000;
	sram_mem[85246] = 16'b0000000000000000;
	sram_mem[85247] = 16'b0000000000000000;
	sram_mem[85248] = 16'b0000000000000000;
	sram_mem[85249] = 16'b0000000000000000;
	sram_mem[85250] = 16'b0000000000000000;
	sram_mem[85251] = 16'b0000000000000000;
	sram_mem[85252] = 16'b0000000000000000;
	sram_mem[85253] = 16'b0000000000000000;
	sram_mem[85254] = 16'b0000000000000000;
	sram_mem[85255] = 16'b0000000000000000;
	sram_mem[85256] = 16'b0000000000000000;
	sram_mem[85257] = 16'b0000000000000000;
	sram_mem[85258] = 16'b0000000000000000;
	sram_mem[85259] = 16'b0000000000000000;
	sram_mem[85260] = 16'b0000000000000000;
	sram_mem[85261] = 16'b0000000000000000;
	sram_mem[85262] = 16'b0000000000000000;
	sram_mem[85263] = 16'b0000000000000000;
	sram_mem[85264] = 16'b0000000000000000;
	sram_mem[85265] = 16'b0000000000000000;
	sram_mem[85266] = 16'b0000000000000000;
	sram_mem[85267] = 16'b0000000000000000;
	sram_mem[85268] = 16'b0000000000000000;
	sram_mem[85269] = 16'b0000000000000000;
	sram_mem[85270] = 16'b0000000000000000;
	sram_mem[85271] = 16'b0000000000000000;
	sram_mem[85272] = 16'b0000000000000000;
	sram_mem[85273] = 16'b0000000000000000;
	sram_mem[85274] = 16'b0000000000000000;
	sram_mem[85275] = 16'b0000000000000000;
	sram_mem[85276] = 16'b0000000000000000;
	sram_mem[85277] = 16'b0000000000000000;
	sram_mem[85278] = 16'b0000000000000000;
	sram_mem[85279] = 16'b0000000000000000;
	sram_mem[85280] = 16'b0000000000000000;
	sram_mem[85281] = 16'b0000000000000000;
	sram_mem[85282] = 16'b0000000000000000;
	sram_mem[85283] = 16'b0000000000000000;
	sram_mem[85284] = 16'b0000000000000000;
	sram_mem[85285] = 16'b0000000000000000;
	sram_mem[85286] = 16'b0000000000000000;
	sram_mem[85287] = 16'b0000000000000000;
	sram_mem[85288] = 16'b0000000000000000;
	sram_mem[85289] = 16'b0000000000000000;
	sram_mem[85290] = 16'b0000000000000000;
	sram_mem[85291] = 16'b0000000000000000;
	sram_mem[85292] = 16'b0000000000000000;
	sram_mem[85293] = 16'b0000000000000000;
	sram_mem[85294] = 16'b0000000000000000;
	sram_mem[85295] = 16'b0000000000000000;
	sram_mem[85296] = 16'b0000000000000000;
	sram_mem[85297] = 16'b0000000000000000;
	sram_mem[85298] = 16'b0000000000000000;
	sram_mem[85299] = 16'b0000000000000000;
	sram_mem[85300] = 16'b0000000000000000;
	sram_mem[85301] = 16'b0000000000000000;
	sram_mem[85302] = 16'b0000000000000000;
	sram_mem[85303] = 16'b0000000000000000;
	sram_mem[85304] = 16'b0000000000000000;
	sram_mem[85305] = 16'b0000000000000000;
	sram_mem[85306] = 16'b0000000000000000;
	sram_mem[85307] = 16'b0000000000000000;
	sram_mem[85308] = 16'b0000000000000000;
	sram_mem[85309] = 16'b0000000000000000;
	sram_mem[85310] = 16'b0000000000000000;
	sram_mem[85311] = 16'b0000000000000000;
	sram_mem[85312] = 16'b0000000000000000;
	sram_mem[85313] = 16'b0000000000000000;
	sram_mem[85314] = 16'b0000000000000000;
	sram_mem[85315] = 16'b0000000000000000;
	sram_mem[85316] = 16'b0000000000000000;
	sram_mem[85317] = 16'b0000000000000000;
	sram_mem[85318] = 16'b0000000000000000;
	sram_mem[85319] = 16'b0000000000000000;
	sram_mem[85320] = 16'b0000000000000000;
	sram_mem[85321] = 16'b0000000000000000;
	sram_mem[85322] = 16'b0000000000000000;
	sram_mem[85323] = 16'b0000000000000000;
	sram_mem[85324] = 16'b0000000000000000;
	sram_mem[85325] = 16'b0000000000000000;
	sram_mem[85326] = 16'b0000000000000000;
	sram_mem[85327] = 16'b0000000000000000;
	sram_mem[85328] = 16'b0000000000000000;
	sram_mem[85329] = 16'b0000000000000000;
	sram_mem[85330] = 16'b0000000000000000;
	sram_mem[85331] = 16'b0000000000000000;
	sram_mem[85332] = 16'b0000000000000000;
	sram_mem[85333] = 16'b0000000000000000;
	sram_mem[85334] = 16'b0000000000000000;
	sram_mem[85335] = 16'b0000000000000000;
	sram_mem[85336] = 16'b0000000000000000;
	sram_mem[85337] = 16'b0000000000000000;
	sram_mem[85338] = 16'b0000000000000000;
	sram_mem[85339] = 16'b0000000000000000;
	sram_mem[85340] = 16'b0000000000000000;
	sram_mem[85341] = 16'b0000000000000000;
	sram_mem[85342] = 16'b0000000000000000;
	sram_mem[85343] = 16'b0000000000000000;
	sram_mem[85344] = 16'b0000000000000000;
	sram_mem[85345] = 16'b0000000000000000;
	sram_mem[85346] = 16'b0000000000000000;
	sram_mem[85347] = 16'b0000000000000000;
	sram_mem[85348] = 16'b0000000000000000;
	sram_mem[85349] = 16'b0000000000000000;
	sram_mem[85350] = 16'b0000000000000000;
	sram_mem[85351] = 16'b0000000000000000;
	sram_mem[85352] = 16'b0000000000000000;
	sram_mem[85353] = 16'b0000000000000000;
	sram_mem[85354] = 16'b0000000000000000;
	sram_mem[85355] = 16'b0000000000000000;
	sram_mem[85356] = 16'b0000000000000000;
	sram_mem[85357] = 16'b0000000000000000;
	sram_mem[85358] = 16'b0000000000000000;
	sram_mem[85359] = 16'b0000000000000000;
	sram_mem[85360] = 16'b0000000000000000;
	sram_mem[85361] = 16'b0000000000000000;
	sram_mem[85362] = 16'b0000000000000000;
	sram_mem[85363] = 16'b0000000000000000;
	sram_mem[85364] = 16'b0000000000000000;
	sram_mem[85365] = 16'b0000000000000000;
	sram_mem[85366] = 16'b0000000000000000;
	sram_mem[85367] = 16'b0000000000000000;
	sram_mem[85368] = 16'b0000000000000000;
	sram_mem[85369] = 16'b0000000000000000;
	sram_mem[85370] = 16'b0000000000000000;
	sram_mem[85371] = 16'b0000000000000000;
	sram_mem[85372] = 16'b0000000000000000;
	sram_mem[85373] = 16'b0000000000000000;
	sram_mem[85374] = 16'b0000000000000000;
	sram_mem[85375] = 16'b0000000000000000;
	sram_mem[85376] = 16'b0000000000000000;
	sram_mem[85377] = 16'b0000000000000000;
	sram_mem[85378] = 16'b0000000000000000;
	sram_mem[85379] = 16'b0000000000000000;
	sram_mem[85380] = 16'b0000000000000000;
	sram_mem[85381] = 16'b0000000000000000;
	sram_mem[85382] = 16'b0000000000000000;
	sram_mem[85383] = 16'b0000000000000000;
	sram_mem[85384] = 16'b0000000000000000;
	sram_mem[85385] = 16'b0000000000000000;
	sram_mem[85386] = 16'b0000000000000000;
	sram_mem[85387] = 16'b0000000000000000;
	sram_mem[85388] = 16'b0000000000000000;
	sram_mem[85389] = 16'b0000000000000000;
	sram_mem[85390] = 16'b0000000000000000;
	sram_mem[85391] = 16'b0000000000000000;
	sram_mem[85392] = 16'b0000000000000000;
	sram_mem[85393] = 16'b0000000000000000;
	sram_mem[85394] = 16'b0000000000000000;
	sram_mem[85395] = 16'b0000000000000000;
	sram_mem[85396] = 16'b0000000000000000;
	sram_mem[85397] = 16'b0000000000000000;
	sram_mem[85398] = 16'b0000000000000000;
	sram_mem[85399] = 16'b0000000000000000;
	sram_mem[85400] = 16'b0000000000000000;
	sram_mem[85401] = 16'b0000000000000000;
	sram_mem[85402] = 16'b0000000000000000;
	sram_mem[85403] = 16'b0000000000000000;
	sram_mem[85404] = 16'b0000000000000000;
	sram_mem[85405] = 16'b0000000000000000;
	sram_mem[85406] = 16'b0000000000000000;
	sram_mem[85407] = 16'b0000000000000000;
	sram_mem[85408] = 16'b0000000000000000;
	sram_mem[85409] = 16'b0000000000000000;
	sram_mem[85410] = 16'b0000000000000000;
	sram_mem[85411] = 16'b0000000000000000;
	sram_mem[85412] = 16'b0000000000000000;
	sram_mem[85413] = 16'b0000000000000000;
	sram_mem[85414] = 16'b0000000000000000;
	sram_mem[85415] = 16'b0000000000000000;
	sram_mem[85416] = 16'b0000000000000000;
	sram_mem[85417] = 16'b0000000000000000;
	sram_mem[85418] = 16'b0000000000000000;
	sram_mem[85419] = 16'b0000000000000000;
	sram_mem[85420] = 16'b0000000000000000;
	sram_mem[85421] = 16'b0000000000000000;
	sram_mem[85422] = 16'b0000000000000000;
	sram_mem[85423] = 16'b0000000000000000;
	sram_mem[85424] = 16'b0000000000000000;
	sram_mem[85425] = 16'b0000000000000000;
	sram_mem[85426] = 16'b0000000000000000;
	sram_mem[85427] = 16'b0000000000000000;
	sram_mem[85428] = 16'b0000000000000000;
	sram_mem[85429] = 16'b0000000000000000;
	sram_mem[85430] = 16'b0000000000000000;
	sram_mem[85431] = 16'b0000000000000000;
	sram_mem[85432] = 16'b0000000000000000;
	sram_mem[85433] = 16'b0000000000000000;
	sram_mem[85434] = 16'b0000000000000000;
	sram_mem[85435] = 16'b0000000000000000;
	sram_mem[85436] = 16'b0000000000000000;
	sram_mem[85437] = 16'b0000000000000000;
	sram_mem[85438] = 16'b0000000000000000;
	sram_mem[85439] = 16'b0000000000000000;
	sram_mem[85440] = 16'b0000000000000000;
	sram_mem[85441] = 16'b0000000000000000;
	sram_mem[85442] = 16'b0000000000000000;
	sram_mem[85443] = 16'b0000000000000000;
	sram_mem[85444] = 16'b0000000000000000;
	sram_mem[85445] = 16'b0000000000000000;
	sram_mem[85446] = 16'b0000000000000000;
	sram_mem[85447] = 16'b0000000000000000;
	sram_mem[85448] = 16'b0000000000000000;
	sram_mem[85449] = 16'b0000000000000000;
	sram_mem[85450] = 16'b0000000000000000;
	sram_mem[85451] = 16'b0000000000000000;
	sram_mem[85452] = 16'b0000000000000000;
	sram_mem[85453] = 16'b0000000000000000;
	sram_mem[85454] = 16'b0000000000000000;
	sram_mem[85455] = 16'b0000000000000000;
	sram_mem[85456] = 16'b0000000000000000;
	sram_mem[85457] = 16'b0000000000000000;
	sram_mem[85458] = 16'b0000000000000000;
	sram_mem[85459] = 16'b0000000000000000;
	sram_mem[85460] = 16'b0000000000000000;
	sram_mem[85461] = 16'b0000000000000000;
	sram_mem[85462] = 16'b0000000000000000;
	sram_mem[85463] = 16'b0000000000000000;
	sram_mem[85464] = 16'b0000000000000000;
	sram_mem[85465] = 16'b0000000000000000;
	sram_mem[85466] = 16'b0000000000000000;
	sram_mem[85467] = 16'b0000000000000000;
	sram_mem[85468] = 16'b0000000000000000;
	sram_mem[85469] = 16'b0000000000000000;
	sram_mem[85470] = 16'b0000000000000000;
	sram_mem[85471] = 16'b0000000000000000;
	sram_mem[85472] = 16'b0000000000000000;
	sram_mem[85473] = 16'b0000000000000000;
	sram_mem[85474] = 16'b0000000000000000;
	sram_mem[85475] = 16'b0000000000000000;
	sram_mem[85476] = 16'b0000000000000000;
	sram_mem[85477] = 16'b0000000000000000;
	sram_mem[85478] = 16'b0000000000000000;
	sram_mem[85479] = 16'b0000000000000000;
	sram_mem[85480] = 16'b0000000000000000;
	sram_mem[85481] = 16'b0000000000000000;
	sram_mem[85482] = 16'b0000000000000000;
	sram_mem[85483] = 16'b0000000000000000;
	sram_mem[85484] = 16'b0000000000000000;
	sram_mem[85485] = 16'b0000000000000000;
	sram_mem[85486] = 16'b0000000000000000;
	sram_mem[85487] = 16'b0000000000000000;
	sram_mem[85488] = 16'b0000000000000000;
	sram_mem[85489] = 16'b0000000000000000;
	sram_mem[85490] = 16'b0000000000000000;
	sram_mem[85491] = 16'b0000000000000000;
	sram_mem[85492] = 16'b0000000000000000;
	sram_mem[85493] = 16'b0000000000000000;
	sram_mem[85494] = 16'b0000000000000000;
	sram_mem[85495] = 16'b0000000000000000;
	sram_mem[85496] = 16'b0000000000000000;
	sram_mem[85497] = 16'b0000000000000000;
	sram_mem[85498] = 16'b0000000000000000;
	sram_mem[85499] = 16'b0000000000000000;
	sram_mem[85500] = 16'b0000000000000000;
	sram_mem[85501] = 16'b0000000000000000;
	sram_mem[85502] = 16'b0000000000000000;
	sram_mem[85503] = 16'b0000000000000000;
	sram_mem[85504] = 16'b0000000000000000;
	sram_mem[85505] = 16'b0000000000000000;
	sram_mem[85506] = 16'b0000000000000000;
	sram_mem[85507] = 16'b0000000000000000;
	sram_mem[85508] = 16'b0000000000000000;
	sram_mem[85509] = 16'b0000000000000000;
	sram_mem[85510] = 16'b0000000000000000;
	sram_mem[85511] = 16'b0000000000000000;
	sram_mem[85512] = 16'b0000000000000000;
	sram_mem[85513] = 16'b0000000000000000;
	sram_mem[85514] = 16'b0000000000000000;
	sram_mem[85515] = 16'b0000000000000000;
	sram_mem[85516] = 16'b0000000000000000;
	sram_mem[85517] = 16'b0000000000000000;
	sram_mem[85518] = 16'b0000000000000000;
	sram_mem[85519] = 16'b0000000000000000;
	sram_mem[85520] = 16'b0000000000000000;
	sram_mem[85521] = 16'b0000000000000000;
	sram_mem[85522] = 16'b0000000000000000;
	sram_mem[85523] = 16'b0000000000000000;
	sram_mem[85524] = 16'b0000000000000000;
	sram_mem[85525] = 16'b0000000000000000;
	sram_mem[85526] = 16'b0000000000000000;
	sram_mem[85527] = 16'b0000000000000000;
	sram_mem[85528] = 16'b0000000000000000;
	sram_mem[85529] = 16'b0000000000000000;
	sram_mem[85530] = 16'b0000000000000000;
	sram_mem[85531] = 16'b0000000000000000;
	sram_mem[85532] = 16'b0000000000000000;
	sram_mem[85533] = 16'b0000000000000000;
	sram_mem[85534] = 16'b0000000000000000;
	sram_mem[85535] = 16'b0000000000000000;
	sram_mem[85536] = 16'b0000000000000000;
	sram_mem[85537] = 16'b0000000000000000;
	sram_mem[85538] = 16'b0000000000000000;
	sram_mem[85539] = 16'b0000000000000000;
	sram_mem[85540] = 16'b0000000000000000;
	sram_mem[85541] = 16'b0000000000000000;
	sram_mem[85542] = 16'b0000000000000000;
	sram_mem[85543] = 16'b0000000000000000;
	sram_mem[85544] = 16'b0000000000000000;
	sram_mem[85545] = 16'b0000000000000000;
	sram_mem[85546] = 16'b0000000000000000;
	sram_mem[85547] = 16'b0000000000000000;
	sram_mem[85548] = 16'b0000000000000000;
	sram_mem[85549] = 16'b0000000000000000;
	sram_mem[85550] = 16'b0000000000000000;
	sram_mem[85551] = 16'b0000000000000000;
	sram_mem[85552] = 16'b0000000000000000;
	sram_mem[85553] = 16'b0000000000000000;
	sram_mem[85554] = 16'b0000000000000000;
	sram_mem[85555] = 16'b0000000000000000;
	sram_mem[85556] = 16'b0000000000000000;
	sram_mem[85557] = 16'b0000000000000000;
	sram_mem[85558] = 16'b0000000000000000;
	sram_mem[85559] = 16'b0000000000000000;
	sram_mem[85560] = 16'b0000000000000000;
	sram_mem[85561] = 16'b0000000000000000;
	sram_mem[85562] = 16'b0000000000000000;
	sram_mem[85563] = 16'b0000000000000000;
	sram_mem[85564] = 16'b0000000000000000;
	sram_mem[85565] = 16'b0000000000000000;
	sram_mem[85566] = 16'b0000000000000000;
	sram_mem[85567] = 16'b0000000000000000;
	sram_mem[85568] = 16'b0000000000000000;
	sram_mem[85569] = 16'b0000000000000000;
	sram_mem[85570] = 16'b0000000000000000;
	sram_mem[85571] = 16'b0000000000000000;
	sram_mem[85572] = 16'b0000000000000000;
	sram_mem[85573] = 16'b0000000000000000;
	sram_mem[85574] = 16'b0000000000000000;
	sram_mem[85575] = 16'b0000000000000000;
	sram_mem[85576] = 16'b0000000000000000;
	sram_mem[85577] = 16'b0000000000000000;
	sram_mem[85578] = 16'b0000000000000000;
	sram_mem[85579] = 16'b0000000000000000;
	sram_mem[85580] = 16'b0000000000000000;
	sram_mem[85581] = 16'b0000000000000000;
	sram_mem[85582] = 16'b0000000000000000;
	sram_mem[85583] = 16'b0000000000000000;
	sram_mem[85584] = 16'b0000000000000000;
	sram_mem[85585] = 16'b0000000000000000;
	sram_mem[85586] = 16'b0000000000000000;
	sram_mem[85587] = 16'b0000000000000000;
	sram_mem[85588] = 16'b0000000000000000;
	sram_mem[85589] = 16'b0000000000000000;
	sram_mem[85590] = 16'b0000000000000000;
	sram_mem[85591] = 16'b0000000000000000;
	sram_mem[85592] = 16'b0000000000000000;
	sram_mem[85593] = 16'b0000000000000000;
	sram_mem[85594] = 16'b0000000000000000;
	sram_mem[85595] = 16'b0000000000000000;
	sram_mem[85596] = 16'b0000000000000000;
	sram_mem[85597] = 16'b0000000000000000;
	sram_mem[85598] = 16'b0000000000000000;
	sram_mem[85599] = 16'b0000000000000000;
	sram_mem[85600] = 16'b0000000000000000;
	sram_mem[85601] = 16'b0000000000000000;
	sram_mem[85602] = 16'b0000000000000000;
	sram_mem[85603] = 16'b0000000000000000;
	sram_mem[85604] = 16'b0000000000000000;
	sram_mem[85605] = 16'b0000000000000000;
	sram_mem[85606] = 16'b0000000000000000;
	sram_mem[85607] = 16'b0000000000000000;
	sram_mem[85608] = 16'b0000000000000000;
	sram_mem[85609] = 16'b0000000000000000;
	sram_mem[85610] = 16'b0000000000000000;
	sram_mem[85611] = 16'b0000000000000000;
	sram_mem[85612] = 16'b0000000000000000;
	sram_mem[85613] = 16'b0000000000000000;
	sram_mem[85614] = 16'b0000000000000000;
	sram_mem[85615] = 16'b0000000000000000;
	sram_mem[85616] = 16'b0000000000000000;
	sram_mem[85617] = 16'b0000000000000000;
	sram_mem[85618] = 16'b0000000000000000;
	sram_mem[85619] = 16'b0000000000000000;
	sram_mem[85620] = 16'b0000000000000000;
	sram_mem[85621] = 16'b0000000000000000;
	sram_mem[85622] = 16'b0000000000000000;
	sram_mem[85623] = 16'b0000000000000000;
	sram_mem[85624] = 16'b0000000000000000;
	sram_mem[85625] = 16'b0000000000000000;
	sram_mem[85626] = 16'b0000000000000000;
	sram_mem[85627] = 16'b0000000000000000;
	sram_mem[85628] = 16'b0000000000000000;
	sram_mem[85629] = 16'b0000000000000000;
	sram_mem[85630] = 16'b0000000000000000;
	sram_mem[85631] = 16'b0000000000000000;
	sram_mem[85632] = 16'b0000000000000000;
	sram_mem[85633] = 16'b0000000000000000;
	sram_mem[85634] = 16'b0000000000000000;
	sram_mem[85635] = 16'b0000000000000000;
	sram_mem[85636] = 16'b0000000000000000;
	sram_mem[85637] = 16'b0000000000000000;
	sram_mem[85638] = 16'b0000000000000000;
	sram_mem[85639] = 16'b0000000000000000;
	sram_mem[85640] = 16'b0000000000000000;
	sram_mem[85641] = 16'b0000000000000000;
	sram_mem[85642] = 16'b0000000000000000;
	sram_mem[85643] = 16'b0000000000000000;
	sram_mem[85644] = 16'b0000000000000000;
	sram_mem[85645] = 16'b0000000000000000;
	sram_mem[85646] = 16'b0000000000000000;
	sram_mem[85647] = 16'b0000000000000000;
	sram_mem[85648] = 16'b0000000000000000;
	sram_mem[85649] = 16'b0000000000000000;
	sram_mem[85650] = 16'b0000000000000000;
	sram_mem[85651] = 16'b0000000000000000;
	sram_mem[85652] = 16'b0000000000000000;
	sram_mem[85653] = 16'b0000000000000000;
	sram_mem[85654] = 16'b0000000000000000;
	sram_mem[85655] = 16'b0000000000000000;
	sram_mem[85656] = 16'b0000000000000000;
	sram_mem[85657] = 16'b0000000000000000;
	sram_mem[85658] = 16'b0000000000000000;
	sram_mem[85659] = 16'b0000000000000000;
	sram_mem[85660] = 16'b0000000000000000;
	sram_mem[85661] = 16'b0000000000000000;
	sram_mem[85662] = 16'b0000000000000000;
	sram_mem[85663] = 16'b0000000000000000;
	sram_mem[85664] = 16'b0000000000000000;
	sram_mem[85665] = 16'b0000000000000000;
	sram_mem[85666] = 16'b0000000000000000;
	sram_mem[85667] = 16'b0000000000000000;
	sram_mem[85668] = 16'b0000000000000000;
	sram_mem[85669] = 16'b0000000000000000;
	sram_mem[85670] = 16'b0000000000000000;
	sram_mem[85671] = 16'b0000000000000000;
	sram_mem[85672] = 16'b0000000000000000;
	sram_mem[85673] = 16'b0000000000000000;
	sram_mem[85674] = 16'b0000000000000000;
	sram_mem[85675] = 16'b0000000000000000;
	sram_mem[85676] = 16'b0000000000000000;
	sram_mem[85677] = 16'b0000000000000000;
	sram_mem[85678] = 16'b0000000000000000;
	sram_mem[85679] = 16'b0000000000000000;
	sram_mem[85680] = 16'b0000000000000000;
	sram_mem[85681] = 16'b0000000000000000;
	sram_mem[85682] = 16'b0000000000000000;
	sram_mem[85683] = 16'b0000000000000000;
	sram_mem[85684] = 16'b0000000000000000;
	sram_mem[85685] = 16'b0000000000000000;
	sram_mem[85686] = 16'b0000000000000000;
	sram_mem[85687] = 16'b0000000000000000;
	sram_mem[85688] = 16'b0000000000000000;
	sram_mem[85689] = 16'b0000000000000000;
	sram_mem[85690] = 16'b0000000000000000;
	sram_mem[85691] = 16'b0000000000000000;
	sram_mem[85692] = 16'b0000000000000000;
	sram_mem[85693] = 16'b0000000000000000;
	sram_mem[85694] = 16'b0000000000000000;
	sram_mem[85695] = 16'b0000000000000000;
	sram_mem[85696] = 16'b0000000000000000;
	sram_mem[85697] = 16'b0000000000000000;
	sram_mem[85698] = 16'b0000000000000000;
	sram_mem[85699] = 16'b0000000000000000;
	sram_mem[85700] = 16'b0000000000000000;
	sram_mem[85701] = 16'b0000000000000000;
	sram_mem[85702] = 16'b0000000000000000;
	sram_mem[85703] = 16'b0000000000000000;
	sram_mem[85704] = 16'b0000000000000000;
	sram_mem[85705] = 16'b0000000000000000;
	sram_mem[85706] = 16'b0000000000000000;
	sram_mem[85707] = 16'b0000000000000000;
	sram_mem[85708] = 16'b0000000000000000;
	sram_mem[85709] = 16'b0000000000000000;
	sram_mem[85710] = 16'b0000000000000000;
	sram_mem[85711] = 16'b0000000000000000;
	sram_mem[85712] = 16'b0000000000000000;
	sram_mem[85713] = 16'b0000000000000000;
	sram_mem[85714] = 16'b0000000000000000;
	sram_mem[85715] = 16'b0000000000000000;
	sram_mem[85716] = 16'b0000000000000000;
	sram_mem[85717] = 16'b0000000000000000;
	sram_mem[85718] = 16'b0000000000000000;
	sram_mem[85719] = 16'b0000000000000000;
	sram_mem[85720] = 16'b0000000000000000;
	sram_mem[85721] = 16'b0000000000000000;
	sram_mem[85722] = 16'b0000000000000000;
	sram_mem[85723] = 16'b0000000000000000;
	sram_mem[85724] = 16'b0000000000000000;
	sram_mem[85725] = 16'b0000000000000000;
	sram_mem[85726] = 16'b0000000000000000;
	sram_mem[85727] = 16'b0000000000000000;
	sram_mem[85728] = 16'b0000000000000000;
	sram_mem[85729] = 16'b0000000000000000;
	sram_mem[85730] = 16'b0000000000000000;
	sram_mem[85731] = 16'b0000000000000000;
	sram_mem[85732] = 16'b0000000000000000;
	sram_mem[85733] = 16'b0000000000000000;
	sram_mem[85734] = 16'b0000000000000000;
	sram_mem[85735] = 16'b0000000000000000;
	sram_mem[85736] = 16'b0000000000000000;
	sram_mem[85737] = 16'b0000000000000000;
	sram_mem[85738] = 16'b0000000000000000;
	sram_mem[85739] = 16'b0000000000000000;
	sram_mem[85740] = 16'b0000000000000000;
	sram_mem[85741] = 16'b0000000000000000;
	sram_mem[85742] = 16'b0000000000000000;
	sram_mem[85743] = 16'b0000000000000000;
	sram_mem[85744] = 16'b0000000000000000;
	sram_mem[85745] = 16'b0000000000000000;
	sram_mem[85746] = 16'b0000000000000000;
	sram_mem[85747] = 16'b0000000000000000;
	sram_mem[85748] = 16'b0000000000000000;
	sram_mem[85749] = 16'b0000000000000000;
	sram_mem[85750] = 16'b0000000000000000;
	sram_mem[85751] = 16'b0000000000000000;
	sram_mem[85752] = 16'b0000000000000000;
	sram_mem[85753] = 16'b0000000000000000;
	sram_mem[85754] = 16'b0000000000000000;
	sram_mem[85755] = 16'b0000000000000000;
	sram_mem[85756] = 16'b0000000000000000;
	sram_mem[85757] = 16'b0000000000000000;
	sram_mem[85758] = 16'b0000000000000000;
	sram_mem[85759] = 16'b0000000000000000;
	sram_mem[85760] = 16'b0000000000000000;
	sram_mem[85761] = 16'b0000000000000000;
	sram_mem[85762] = 16'b0000000000000000;
	sram_mem[85763] = 16'b0000000000000000;
	sram_mem[85764] = 16'b0000000000000000;
	sram_mem[85765] = 16'b0000000000000000;
	sram_mem[85766] = 16'b0000000000000000;
	sram_mem[85767] = 16'b0000000000000000;
	sram_mem[85768] = 16'b0000000000000000;
	sram_mem[85769] = 16'b0000000000000000;
	sram_mem[85770] = 16'b0000000000000000;
	sram_mem[85771] = 16'b0000000000000000;
	sram_mem[85772] = 16'b0000000000000000;
	sram_mem[85773] = 16'b0000000000000000;
	sram_mem[85774] = 16'b0000000000000000;
	sram_mem[85775] = 16'b0000000000000000;
	sram_mem[85776] = 16'b0000000000000000;
	sram_mem[85777] = 16'b0000000000000000;
	sram_mem[85778] = 16'b0000000000000000;
	sram_mem[85779] = 16'b0000000000000000;
	sram_mem[85780] = 16'b0000000000000000;
	sram_mem[85781] = 16'b0000000000000000;
	sram_mem[85782] = 16'b0000000000000000;
	sram_mem[85783] = 16'b0000000000000000;
	sram_mem[85784] = 16'b0000000000000000;
	sram_mem[85785] = 16'b0000000000000000;
	sram_mem[85786] = 16'b0000000000000000;
	sram_mem[85787] = 16'b0000000000000000;
	sram_mem[85788] = 16'b0000000000000000;
	sram_mem[85789] = 16'b0000000000000000;
	sram_mem[85790] = 16'b0000000000000000;
	sram_mem[85791] = 16'b0000000000000000;
	sram_mem[85792] = 16'b0000000000000000;
	sram_mem[85793] = 16'b0000000000000000;
	sram_mem[85794] = 16'b0000000000000000;
	sram_mem[85795] = 16'b0000000000000000;
	sram_mem[85796] = 16'b0000000000000000;
	sram_mem[85797] = 16'b0000000000000000;
	sram_mem[85798] = 16'b0000000000000000;
	sram_mem[85799] = 16'b0000000000000000;
	sram_mem[85800] = 16'b0000000000000000;
	sram_mem[85801] = 16'b0000000000000000;
	sram_mem[85802] = 16'b0000000000000000;
	sram_mem[85803] = 16'b0000000000000000;
	sram_mem[85804] = 16'b0000000000000000;
	sram_mem[85805] = 16'b0000000000000000;
	sram_mem[85806] = 16'b0000000000000000;
	sram_mem[85807] = 16'b0000000000000000;
	sram_mem[85808] = 16'b0000000000000000;
	sram_mem[85809] = 16'b0000000000000000;
	sram_mem[85810] = 16'b0000000000000000;
	sram_mem[85811] = 16'b0000000000000000;
	sram_mem[85812] = 16'b0000000000000000;
	sram_mem[85813] = 16'b0000000000000000;
	sram_mem[85814] = 16'b0000000000000000;
	sram_mem[85815] = 16'b0000000000000000;
	sram_mem[85816] = 16'b0000000000000000;
	sram_mem[85817] = 16'b0000000000000000;
	sram_mem[85818] = 16'b0000000000000000;
	sram_mem[85819] = 16'b0000000000000000;
	sram_mem[85820] = 16'b0000000000000000;
	sram_mem[85821] = 16'b0000000000000000;
	sram_mem[85822] = 16'b0000000000000000;
	sram_mem[85823] = 16'b0000000000000000;
	sram_mem[85824] = 16'b0000000000000000;
	sram_mem[85825] = 16'b0000000000000000;
	sram_mem[85826] = 16'b0000000000000000;
	sram_mem[85827] = 16'b0000000000000000;
	sram_mem[85828] = 16'b0000000000000000;
	sram_mem[85829] = 16'b0000000000000000;
	sram_mem[85830] = 16'b0000000000000000;
	sram_mem[85831] = 16'b0000000000000000;
	sram_mem[85832] = 16'b0000000000000000;
	sram_mem[85833] = 16'b0000000000000000;
	sram_mem[85834] = 16'b0000000000000000;
	sram_mem[85835] = 16'b0000000000000000;
	sram_mem[85836] = 16'b0000000000000000;
	sram_mem[85837] = 16'b0000000000000000;
	sram_mem[85838] = 16'b0000000000000000;
	sram_mem[85839] = 16'b0000000000000000;
	sram_mem[85840] = 16'b0000000000000000;
	sram_mem[85841] = 16'b0000000000000000;
	sram_mem[85842] = 16'b0000000000000000;
	sram_mem[85843] = 16'b0000000000000000;
	sram_mem[85844] = 16'b0000000000000000;
	sram_mem[85845] = 16'b0000000000000000;
	sram_mem[85846] = 16'b0000000000000000;
	sram_mem[85847] = 16'b0000000000000000;
	sram_mem[85848] = 16'b0000000000000000;
	sram_mem[85849] = 16'b0000000000000000;
	sram_mem[85850] = 16'b0000000000000000;
	sram_mem[85851] = 16'b0000000000000000;
	sram_mem[85852] = 16'b0000000000000000;
	sram_mem[85853] = 16'b0000000000000000;
	sram_mem[85854] = 16'b0000000000000000;
	sram_mem[85855] = 16'b0000000000000000;
	sram_mem[85856] = 16'b0000000000000000;
	sram_mem[85857] = 16'b0000000000000000;
	sram_mem[85858] = 16'b0000000000000000;
	sram_mem[85859] = 16'b0000000000000000;
	sram_mem[85860] = 16'b0000000000000000;
	sram_mem[85861] = 16'b0000000000000000;
	sram_mem[85862] = 16'b0000000000000000;
	sram_mem[85863] = 16'b0000000000000000;
	sram_mem[85864] = 16'b0000000000000000;
	sram_mem[85865] = 16'b0000000000000000;
	sram_mem[85866] = 16'b0000000000000000;
	sram_mem[85867] = 16'b0000000000000000;
	sram_mem[85868] = 16'b0000000000000000;
	sram_mem[85869] = 16'b0000000000000000;
	sram_mem[85870] = 16'b0000000000000000;
	sram_mem[85871] = 16'b0000000000000000;
	sram_mem[85872] = 16'b0000000000000000;
	sram_mem[85873] = 16'b0000000000000000;
	sram_mem[85874] = 16'b0000000000000000;
	sram_mem[85875] = 16'b0000000000000000;
	sram_mem[85876] = 16'b0000000000000000;
	sram_mem[85877] = 16'b0000000000000000;
	sram_mem[85878] = 16'b0000000000000000;
	sram_mem[85879] = 16'b0000000000000000;
	sram_mem[85880] = 16'b0000000000000000;
	sram_mem[85881] = 16'b0000000000000000;
	sram_mem[85882] = 16'b0000000000000000;
	sram_mem[85883] = 16'b0000000000000000;
	sram_mem[85884] = 16'b0000000000000000;
	sram_mem[85885] = 16'b0000000000000000;
	sram_mem[85886] = 16'b0000000000000000;
	sram_mem[85887] = 16'b0000000000000000;
	sram_mem[85888] = 16'b0000000000000000;
	sram_mem[85889] = 16'b0000000000000000;
	sram_mem[85890] = 16'b0000000000000000;
	sram_mem[85891] = 16'b0000000000000000;
	sram_mem[85892] = 16'b0000000000000000;
	sram_mem[85893] = 16'b0000000000000000;
	sram_mem[85894] = 16'b0000000000000000;
	sram_mem[85895] = 16'b0000000000000000;
	sram_mem[85896] = 16'b0000000000000000;
	sram_mem[85897] = 16'b0000000000000000;
	sram_mem[85898] = 16'b0000000000000000;
	sram_mem[85899] = 16'b0000000000000000;
	sram_mem[85900] = 16'b0000000000000000;
	sram_mem[85901] = 16'b0000000000000000;
	sram_mem[85902] = 16'b0000000000000000;
	sram_mem[85903] = 16'b0000000000000000;
	sram_mem[85904] = 16'b0000000000000000;
	sram_mem[85905] = 16'b0000000000000000;
	sram_mem[85906] = 16'b0000000000000000;
	sram_mem[85907] = 16'b0000000000000000;
	sram_mem[85908] = 16'b0000000000000000;
	sram_mem[85909] = 16'b0000000000000000;
	sram_mem[85910] = 16'b0000000000000000;
	sram_mem[85911] = 16'b0000000000000000;
	sram_mem[85912] = 16'b0000000000000000;
	sram_mem[85913] = 16'b0000000000000000;
	sram_mem[85914] = 16'b0000000000000000;
	sram_mem[85915] = 16'b0000000000000000;
	sram_mem[85916] = 16'b0000000000000000;
	sram_mem[85917] = 16'b0000000000000000;
	sram_mem[85918] = 16'b0000000000000000;
	sram_mem[85919] = 16'b0000000000000000;
	sram_mem[85920] = 16'b0000000000000000;
	sram_mem[85921] = 16'b0000000000000000;
	sram_mem[85922] = 16'b0000000000000000;
	sram_mem[85923] = 16'b0000000000000000;
	sram_mem[85924] = 16'b0000000000000000;
	sram_mem[85925] = 16'b0000000000000000;
	sram_mem[85926] = 16'b0000000000000000;
	sram_mem[85927] = 16'b0000000000000000;
	sram_mem[85928] = 16'b0000000000000000;
	sram_mem[85929] = 16'b0000000000000000;
	sram_mem[85930] = 16'b0000000000000000;
	sram_mem[85931] = 16'b0000000000000000;
	sram_mem[85932] = 16'b0000000000000000;
	sram_mem[85933] = 16'b0000000000000000;
	sram_mem[85934] = 16'b0000000000000000;
	sram_mem[85935] = 16'b0000000000000000;
	sram_mem[85936] = 16'b0000000000000000;
	sram_mem[85937] = 16'b0000000000000000;
	sram_mem[85938] = 16'b0000000000000000;
	sram_mem[85939] = 16'b0000000000000000;
	sram_mem[85940] = 16'b0000000000000000;
	sram_mem[85941] = 16'b0000000000000000;
	sram_mem[85942] = 16'b0000000000000000;
	sram_mem[85943] = 16'b0000000000000000;
	sram_mem[85944] = 16'b0000000000000000;
	sram_mem[85945] = 16'b0000000000000000;
	sram_mem[85946] = 16'b0000000000000000;
	sram_mem[85947] = 16'b0000000000000000;
	sram_mem[85948] = 16'b0000000000000000;
	sram_mem[85949] = 16'b0000000000000000;
	sram_mem[85950] = 16'b0000000000000000;
	sram_mem[85951] = 16'b0000000000000000;
	sram_mem[85952] = 16'b0000000000000000;
	sram_mem[85953] = 16'b0000000000000000;
	sram_mem[85954] = 16'b0000000000000000;
	sram_mem[85955] = 16'b0000000000000000;
	sram_mem[85956] = 16'b0000000000000000;
	sram_mem[85957] = 16'b0000000000000000;
	sram_mem[85958] = 16'b0000000000000000;
	sram_mem[85959] = 16'b0000000000000000;
	sram_mem[85960] = 16'b0000000000000000;
	sram_mem[85961] = 16'b0000000000000000;
	sram_mem[85962] = 16'b0000000000000000;
	sram_mem[85963] = 16'b0000000000000000;
	sram_mem[85964] = 16'b0000000000000000;
	sram_mem[85965] = 16'b0000000000000000;
	sram_mem[85966] = 16'b0000000000000000;
	sram_mem[85967] = 16'b0000000000000000;
	sram_mem[85968] = 16'b0000000000000000;
	sram_mem[85969] = 16'b0000000000000000;
	sram_mem[85970] = 16'b0000000000000000;
	sram_mem[85971] = 16'b0000000000000000;
	sram_mem[85972] = 16'b0000000000000000;
	sram_mem[85973] = 16'b0000000000000000;
	sram_mem[85974] = 16'b0000000000000000;
	sram_mem[85975] = 16'b0000000000000000;
	sram_mem[85976] = 16'b0000000000000000;
	sram_mem[85977] = 16'b0000000000000000;
	sram_mem[85978] = 16'b0000000000000000;
	sram_mem[85979] = 16'b0000000000000000;
	sram_mem[85980] = 16'b0000000000000000;
	sram_mem[85981] = 16'b0000000000000000;
	sram_mem[85982] = 16'b0000000000000000;
	sram_mem[85983] = 16'b0000000000000000;
	sram_mem[85984] = 16'b0000000000000000;
	sram_mem[85985] = 16'b0000000000000000;
	sram_mem[85986] = 16'b0000000000000000;
	sram_mem[85987] = 16'b0000000000000000;
	sram_mem[85988] = 16'b0000000000000000;
	sram_mem[85989] = 16'b0000000000000000;
	sram_mem[85990] = 16'b0000000000000000;
	sram_mem[85991] = 16'b0000000000000000;
	sram_mem[85992] = 16'b0000000000000000;
	sram_mem[85993] = 16'b0000000000000000;
	sram_mem[85994] = 16'b0000000000000000;
	sram_mem[85995] = 16'b0000000000000000;
	sram_mem[85996] = 16'b0000000000000000;
	sram_mem[85997] = 16'b0000000000000000;
	sram_mem[85998] = 16'b0000000000000000;
	sram_mem[85999] = 16'b0000000000000000;
	sram_mem[86000] = 16'b0000000000000000;
	sram_mem[86001] = 16'b0000000000000000;
	sram_mem[86002] = 16'b0000000000000000;
	sram_mem[86003] = 16'b0000000000000000;
	sram_mem[86004] = 16'b0000000000000000;
	sram_mem[86005] = 16'b0000000000000000;
	sram_mem[86006] = 16'b0000000000000000;
	sram_mem[86007] = 16'b0000000000000000;
	sram_mem[86008] = 16'b0000000000000000;
	sram_mem[86009] = 16'b0000000000000000;
	sram_mem[86010] = 16'b0000000000000000;
	sram_mem[86011] = 16'b0000000000000000;
	sram_mem[86012] = 16'b0000000000000000;
	sram_mem[86013] = 16'b0000000000000000;
	sram_mem[86014] = 16'b0000000000000000;
	sram_mem[86015] = 16'b0000000000000000;
	sram_mem[86016] = 16'b0000000000000000;
	sram_mem[86017] = 16'b0000000000000000;
	sram_mem[86018] = 16'b0000000000000000;
	sram_mem[86019] = 16'b0000000000000000;
	sram_mem[86020] = 16'b0000000000000000;
	sram_mem[86021] = 16'b0000000000000000;
	sram_mem[86022] = 16'b0000000000000000;
	sram_mem[86023] = 16'b0000000000000000;
	sram_mem[86024] = 16'b0000000000000000;
	sram_mem[86025] = 16'b0000000000000000;
	sram_mem[86026] = 16'b0000000000000000;
	sram_mem[86027] = 16'b0000000000000000;
	sram_mem[86028] = 16'b0000000000000000;
	sram_mem[86029] = 16'b0000000000000000;
	sram_mem[86030] = 16'b0000000000000000;
	sram_mem[86031] = 16'b0000000000000000;
	sram_mem[86032] = 16'b0000000000000000;
	sram_mem[86033] = 16'b0000000000000000;
	sram_mem[86034] = 16'b0000000000000000;
	sram_mem[86035] = 16'b0000000000000000;
	sram_mem[86036] = 16'b0000000000000000;
	sram_mem[86037] = 16'b0000000000000000;
	sram_mem[86038] = 16'b0000000000000000;
	sram_mem[86039] = 16'b0000000000000000;
	sram_mem[86040] = 16'b0000000000000000;
	sram_mem[86041] = 16'b0000000000000000;
	sram_mem[86042] = 16'b0000000000000000;
	sram_mem[86043] = 16'b0000000000000000;
	sram_mem[86044] = 16'b0000000000000000;
	sram_mem[86045] = 16'b0000000000000000;
	sram_mem[86046] = 16'b0000000000000000;
	sram_mem[86047] = 16'b0000000000000000;
	sram_mem[86048] = 16'b0000000000000000;
	sram_mem[86049] = 16'b0000000000000000;
	sram_mem[86050] = 16'b0000000000000000;
	sram_mem[86051] = 16'b0000000000000000;
	sram_mem[86052] = 16'b0000000000000000;
	sram_mem[86053] = 16'b0000000000000000;
	sram_mem[86054] = 16'b0000000000000000;
	sram_mem[86055] = 16'b0000000000000000;
	sram_mem[86056] = 16'b0000000000000000;
	sram_mem[86057] = 16'b0000000000000000;
	sram_mem[86058] = 16'b0000000000000000;
	sram_mem[86059] = 16'b0000000000000000;
	sram_mem[86060] = 16'b0000000000000000;
	sram_mem[86061] = 16'b0000000000000000;
	sram_mem[86062] = 16'b0000000000000000;
	sram_mem[86063] = 16'b0000000000000000;
	sram_mem[86064] = 16'b0000000000000000;
	sram_mem[86065] = 16'b0000000000000000;
	sram_mem[86066] = 16'b0000000000000000;
	sram_mem[86067] = 16'b0000000000000000;
	sram_mem[86068] = 16'b0000000000000000;
	sram_mem[86069] = 16'b0000000000000000;
	sram_mem[86070] = 16'b0000000000000000;
	sram_mem[86071] = 16'b0000000000000000;
	sram_mem[86072] = 16'b0000000000000000;
	sram_mem[86073] = 16'b0000000000000000;
	sram_mem[86074] = 16'b0000000000000000;
	sram_mem[86075] = 16'b0000000000000000;
	sram_mem[86076] = 16'b0000000000000000;
	sram_mem[86077] = 16'b0000000000000000;
	sram_mem[86078] = 16'b0000000000000000;
	sram_mem[86079] = 16'b0000000000000000;
	sram_mem[86080] = 16'b0000000000000000;
	sram_mem[86081] = 16'b0000000000000000;
	sram_mem[86082] = 16'b0000000000000000;
	sram_mem[86083] = 16'b0000000000000000;
	sram_mem[86084] = 16'b0000000000000000;
	sram_mem[86085] = 16'b0000000000000000;
	sram_mem[86086] = 16'b0000000000000000;
	sram_mem[86087] = 16'b0000000000000000;
	sram_mem[86088] = 16'b0000000000000000;
	sram_mem[86089] = 16'b0000000000000000;
	sram_mem[86090] = 16'b0000000000000000;
	sram_mem[86091] = 16'b0000000000000000;
	sram_mem[86092] = 16'b0000000000000000;
	sram_mem[86093] = 16'b0000000000000000;
	sram_mem[86094] = 16'b0000000000000000;
	sram_mem[86095] = 16'b0000000000000000;
	sram_mem[86096] = 16'b0000000000000000;
	sram_mem[86097] = 16'b0000000000000000;
	sram_mem[86098] = 16'b0000000000000000;
	sram_mem[86099] = 16'b0000000000000000;
	sram_mem[86100] = 16'b0000000000000000;
	sram_mem[86101] = 16'b0000000000000000;
	sram_mem[86102] = 16'b0000000000000000;
	sram_mem[86103] = 16'b0000000000000000;
	sram_mem[86104] = 16'b0000000000000000;
	sram_mem[86105] = 16'b0000000000000000;
	sram_mem[86106] = 16'b0000000000000000;
	sram_mem[86107] = 16'b0000000000000000;
	sram_mem[86108] = 16'b0000000000000000;
	sram_mem[86109] = 16'b0000000000000000;
	sram_mem[86110] = 16'b0000000000000000;
	sram_mem[86111] = 16'b0000000000000000;
	sram_mem[86112] = 16'b0000000000000000;
	sram_mem[86113] = 16'b0000000000000000;
	sram_mem[86114] = 16'b0000000000000000;
	sram_mem[86115] = 16'b0000000000000000;
	sram_mem[86116] = 16'b0000000000000000;
	sram_mem[86117] = 16'b0000000000000000;
	sram_mem[86118] = 16'b0000000000000000;
	sram_mem[86119] = 16'b0000000000000000;
	sram_mem[86120] = 16'b0000000000000000;
	sram_mem[86121] = 16'b0000000000000000;
	sram_mem[86122] = 16'b0000000000000000;
	sram_mem[86123] = 16'b0000000000000000;
	sram_mem[86124] = 16'b0000000000000000;
	sram_mem[86125] = 16'b0000000000000000;
	sram_mem[86126] = 16'b0000000000000000;
	sram_mem[86127] = 16'b0000000000000000;
	sram_mem[86128] = 16'b0000000000000000;
	sram_mem[86129] = 16'b0000000000000000;
	sram_mem[86130] = 16'b0000000000000000;
	sram_mem[86131] = 16'b0000000000000000;
	sram_mem[86132] = 16'b0000000000000000;
	sram_mem[86133] = 16'b0000000000000000;
	sram_mem[86134] = 16'b0000000000000000;
	sram_mem[86135] = 16'b0000000000000000;
	sram_mem[86136] = 16'b0000000000000000;
	sram_mem[86137] = 16'b0000000000000000;
	sram_mem[86138] = 16'b0000000000000000;
	sram_mem[86139] = 16'b0000000000000000;
	sram_mem[86140] = 16'b0000000000000000;
	sram_mem[86141] = 16'b0000000000000000;
	sram_mem[86142] = 16'b0000000000000000;
	sram_mem[86143] = 16'b0000000000000000;
	sram_mem[86144] = 16'b0000000000000000;
	sram_mem[86145] = 16'b0000000000000000;
	sram_mem[86146] = 16'b0000000000000000;
	sram_mem[86147] = 16'b0000000000000000;
	sram_mem[86148] = 16'b0000000000000000;
	sram_mem[86149] = 16'b0000000000000000;
	sram_mem[86150] = 16'b0000000000000000;
	sram_mem[86151] = 16'b0000000000000000;
	sram_mem[86152] = 16'b0000000000000000;
	sram_mem[86153] = 16'b0000000000000000;
	sram_mem[86154] = 16'b0000000000000000;
	sram_mem[86155] = 16'b0000000000000000;
	sram_mem[86156] = 16'b0000000000000000;
	sram_mem[86157] = 16'b0000000000000000;
	sram_mem[86158] = 16'b0000000000000000;
	sram_mem[86159] = 16'b0000000000000000;
	sram_mem[86160] = 16'b0000000000000000;
	sram_mem[86161] = 16'b0000000000000000;
	sram_mem[86162] = 16'b0000000000000000;
	sram_mem[86163] = 16'b0000000000000000;
	sram_mem[86164] = 16'b0000000000000000;
	sram_mem[86165] = 16'b0000000000000000;
	sram_mem[86166] = 16'b0000000000000000;
	sram_mem[86167] = 16'b0000000000000000;
	sram_mem[86168] = 16'b0000000000000000;
	sram_mem[86169] = 16'b0000000000000000;
	sram_mem[86170] = 16'b0000000000000000;
	sram_mem[86171] = 16'b0000000000000000;
	sram_mem[86172] = 16'b0000000000000000;
	sram_mem[86173] = 16'b0000000000000000;
	sram_mem[86174] = 16'b0000000000000000;
	sram_mem[86175] = 16'b0000000000000000;
	sram_mem[86176] = 16'b0000000000000000;
	sram_mem[86177] = 16'b0000000000000000;
	sram_mem[86178] = 16'b0000000000000000;
	sram_mem[86179] = 16'b0000000000000000;
	sram_mem[86180] = 16'b0000000000000000;
	sram_mem[86181] = 16'b0000000000000000;
	sram_mem[86182] = 16'b0000000000000000;
	sram_mem[86183] = 16'b0000000000000000;
	sram_mem[86184] = 16'b0000000000000000;
	sram_mem[86185] = 16'b0000000000000000;
	sram_mem[86186] = 16'b0000000000000000;
	sram_mem[86187] = 16'b0000000000000000;
	sram_mem[86188] = 16'b0000000000000000;
	sram_mem[86189] = 16'b0000000000000000;
	sram_mem[86190] = 16'b0000000000000000;
	sram_mem[86191] = 16'b0000000000000000;
	sram_mem[86192] = 16'b0000000000000000;
	sram_mem[86193] = 16'b0000000000000000;
	sram_mem[86194] = 16'b0000000000000000;
	sram_mem[86195] = 16'b0000000000000000;
	sram_mem[86196] = 16'b0000000000000000;
	sram_mem[86197] = 16'b0000000000000000;
	sram_mem[86198] = 16'b0000000000000000;
	sram_mem[86199] = 16'b0000000000000000;
	sram_mem[86200] = 16'b0000000000000000;
	sram_mem[86201] = 16'b0000000000000000;
	sram_mem[86202] = 16'b0000000000000000;
	sram_mem[86203] = 16'b0000000000000000;
	sram_mem[86204] = 16'b0000000000000000;
	sram_mem[86205] = 16'b0000000000000000;
	sram_mem[86206] = 16'b0000000000000000;
	sram_mem[86207] = 16'b0000000000000000;
	sram_mem[86208] = 16'b0000000000000000;
	sram_mem[86209] = 16'b0000000000000000;
	sram_mem[86210] = 16'b0000000000000000;
	sram_mem[86211] = 16'b0000000000000000;
	sram_mem[86212] = 16'b0000000000000000;
	sram_mem[86213] = 16'b0000000000000000;
	sram_mem[86214] = 16'b0000000000000000;
	sram_mem[86215] = 16'b0000000000000000;
	sram_mem[86216] = 16'b0000000000000000;
	sram_mem[86217] = 16'b0000000000000000;
	sram_mem[86218] = 16'b0000000000000000;
	sram_mem[86219] = 16'b0000000000000000;
	sram_mem[86220] = 16'b0000000000000000;
	sram_mem[86221] = 16'b0000000000000000;
	sram_mem[86222] = 16'b0000000000000000;
	sram_mem[86223] = 16'b0000000000000000;
	sram_mem[86224] = 16'b0000000000000000;
	sram_mem[86225] = 16'b0000000000000000;
	sram_mem[86226] = 16'b0000000000000000;
	sram_mem[86227] = 16'b0000000000000000;
	sram_mem[86228] = 16'b0000000000000000;
	sram_mem[86229] = 16'b0000000000000000;
	sram_mem[86230] = 16'b0000000000000000;
	sram_mem[86231] = 16'b0000000000000000;
	sram_mem[86232] = 16'b0000000000000000;
	sram_mem[86233] = 16'b0000000000000000;
	sram_mem[86234] = 16'b0000000000000000;
	sram_mem[86235] = 16'b0000000000000000;
	sram_mem[86236] = 16'b0000000000000000;
	sram_mem[86237] = 16'b0000000000000000;
	sram_mem[86238] = 16'b0000000000000000;
	sram_mem[86239] = 16'b0000000000000000;
	sram_mem[86240] = 16'b0000000000000000;
	sram_mem[86241] = 16'b0000000000000000;
	sram_mem[86242] = 16'b0000000000000000;
	sram_mem[86243] = 16'b0000000000000000;
	sram_mem[86244] = 16'b0000000000000000;
	sram_mem[86245] = 16'b0000000000000000;
	sram_mem[86246] = 16'b0000000000000000;
	sram_mem[86247] = 16'b0000000000000000;
	sram_mem[86248] = 16'b0000000000000000;
	sram_mem[86249] = 16'b0000000000000000;
	sram_mem[86250] = 16'b0000000000000000;
	sram_mem[86251] = 16'b0000000000000000;
	sram_mem[86252] = 16'b0000000000000000;
	sram_mem[86253] = 16'b0000000000000000;
	sram_mem[86254] = 16'b0000000000000000;
	sram_mem[86255] = 16'b0000000000000000;
	sram_mem[86256] = 16'b0000000000000000;
	sram_mem[86257] = 16'b0000000000000000;
	sram_mem[86258] = 16'b0000000000000000;
	sram_mem[86259] = 16'b0000000000000000;
	sram_mem[86260] = 16'b0000000000000000;
	sram_mem[86261] = 16'b0000000000000000;
	sram_mem[86262] = 16'b0000000000000000;
	sram_mem[86263] = 16'b0000000000000000;
	sram_mem[86264] = 16'b0000000000000000;
	sram_mem[86265] = 16'b0000000000000000;
	sram_mem[86266] = 16'b0000000000000000;
	sram_mem[86267] = 16'b0000000000000000;
	sram_mem[86268] = 16'b0000000000000000;
	sram_mem[86269] = 16'b0000000000000000;
	sram_mem[86270] = 16'b0000000000000000;
	sram_mem[86271] = 16'b0000000000000000;
	sram_mem[86272] = 16'b0000000000000000;
	sram_mem[86273] = 16'b0000000000000000;
	sram_mem[86274] = 16'b0000000000000000;
	sram_mem[86275] = 16'b0000000000000000;
	sram_mem[86276] = 16'b0000000000000000;
	sram_mem[86277] = 16'b0000000000000000;
	sram_mem[86278] = 16'b0000000000000000;
	sram_mem[86279] = 16'b0000000000000000;
	sram_mem[86280] = 16'b0000000000000000;
	sram_mem[86281] = 16'b0000000000000000;
	sram_mem[86282] = 16'b0000000000000000;
	sram_mem[86283] = 16'b0000000000000000;
	sram_mem[86284] = 16'b0000000000000000;
	sram_mem[86285] = 16'b0000000000000000;
	sram_mem[86286] = 16'b0000000000000000;
	sram_mem[86287] = 16'b0000000000000000;
	sram_mem[86288] = 16'b0000000000000000;
	sram_mem[86289] = 16'b0000000000000000;
	sram_mem[86290] = 16'b0000000000000000;
	sram_mem[86291] = 16'b0000000000000000;
	sram_mem[86292] = 16'b0000000000000000;
	sram_mem[86293] = 16'b0000000000000000;
	sram_mem[86294] = 16'b0000000000000000;
	sram_mem[86295] = 16'b0000000000000000;
	sram_mem[86296] = 16'b0000000000000000;
	sram_mem[86297] = 16'b0000000000000000;
	sram_mem[86298] = 16'b0000000000000000;
	sram_mem[86299] = 16'b0000000000000000;
	sram_mem[86300] = 16'b0000000000000000;
	sram_mem[86301] = 16'b0000000000000000;
	sram_mem[86302] = 16'b0000000000000000;
	sram_mem[86303] = 16'b0000000000000000;
	sram_mem[86304] = 16'b0000000000000000;
	sram_mem[86305] = 16'b0000000000000000;
	sram_mem[86306] = 16'b0000000000000000;
	sram_mem[86307] = 16'b0000000000000000;
	sram_mem[86308] = 16'b0000000000000000;
	sram_mem[86309] = 16'b0000000000000000;
	sram_mem[86310] = 16'b0000000000000000;
	sram_mem[86311] = 16'b0000000000000000;
	sram_mem[86312] = 16'b0000000000000000;
	sram_mem[86313] = 16'b0000000000000000;
	sram_mem[86314] = 16'b0000000000000000;
	sram_mem[86315] = 16'b0000000000000000;
	sram_mem[86316] = 16'b0000000000000000;
	sram_mem[86317] = 16'b0000000000000000;
	sram_mem[86318] = 16'b0000000000000000;
	sram_mem[86319] = 16'b0000000000000000;
	sram_mem[86320] = 16'b0000000000000000;
	sram_mem[86321] = 16'b0000000000000000;
	sram_mem[86322] = 16'b0000000000000000;
	sram_mem[86323] = 16'b0000000000000000;
	sram_mem[86324] = 16'b0000000000000000;
	sram_mem[86325] = 16'b0000000000000000;
	sram_mem[86326] = 16'b0000000000000000;
	sram_mem[86327] = 16'b0000000000000000;
	sram_mem[86328] = 16'b0000000000000000;
	sram_mem[86329] = 16'b0000000000000000;
	sram_mem[86330] = 16'b0000000000000000;
	sram_mem[86331] = 16'b0000000000000000;
	sram_mem[86332] = 16'b0000000000000000;
	sram_mem[86333] = 16'b0000000000000000;
	sram_mem[86334] = 16'b0000000000000000;
	sram_mem[86335] = 16'b0000000000000000;
	sram_mem[86336] = 16'b0000000000000000;
	sram_mem[86337] = 16'b0000000000000000;
	sram_mem[86338] = 16'b0000000000000000;
	sram_mem[86339] = 16'b0000000000000000;
	sram_mem[86340] = 16'b0000000000000000;
	sram_mem[86341] = 16'b0000000000000000;
	sram_mem[86342] = 16'b0000000000000000;
	sram_mem[86343] = 16'b0000000000000000;
	sram_mem[86344] = 16'b0000000000000000;
	sram_mem[86345] = 16'b0000000000000000;
	sram_mem[86346] = 16'b0000000000000000;
	sram_mem[86347] = 16'b0000000000000000;
	sram_mem[86348] = 16'b0000000000000000;
	sram_mem[86349] = 16'b0000000000000000;
	sram_mem[86350] = 16'b0000000000000000;
	sram_mem[86351] = 16'b0000000000000000;
	sram_mem[86352] = 16'b0000000000000000;
	sram_mem[86353] = 16'b0000000000000000;
	sram_mem[86354] = 16'b0000000000000000;
	sram_mem[86355] = 16'b0000000000000000;
	sram_mem[86356] = 16'b0000000000000000;
	sram_mem[86357] = 16'b0000000000000000;
	sram_mem[86358] = 16'b0000000000000000;
	sram_mem[86359] = 16'b0000000000000000;
	sram_mem[86360] = 16'b0000000000000000;
	sram_mem[86361] = 16'b0000000000000000;
	sram_mem[86362] = 16'b0000000000000000;
	sram_mem[86363] = 16'b0000000000000000;
	sram_mem[86364] = 16'b0000000000000000;
	sram_mem[86365] = 16'b0000000000000000;
	sram_mem[86366] = 16'b0000000000000000;
	sram_mem[86367] = 16'b0000000000000000;
	sram_mem[86368] = 16'b0000000000000000;
	sram_mem[86369] = 16'b0000000000000000;
	sram_mem[86370] = 16'b0000000000000000;
	sram_mem[86371] = 16'b0000000000000000;
	sram_mem[86372] = 16'b0000000000000000;
	sram_mem[86373] = 16'b0000000000000000;
	sram_mem[86374] = 16'b0000000000000000;
	sram_mem[86375] = 16'b0000000000000000;
	sram_mem[86376] = 16'b0000000000000000;
	sram_mem[86377] = 16'b0000000000000000;
	sram_mem[86378] = 16'b0000000000000000;
	sram_mem[86379] = 16'b0000000000000000;
	sram_mem[86380] = 16'b0000000000000000;
	sram_mem[86381] = 16'b0000000000000000;
	sram_mem[86382] = 16'b0000000000000000;
	sram_mem[86383] = 16'b0000000000000000;
	sram_mem[86384] = 16'b0000000000000000;
	sram_mem[86385] = 16'b0000000000000000;
	sram_mem[86386] = 16'b0000000000000000;
	sram_mem[86387] = 16'b0000000000000000;
	sram_mem[86388] = 16'b0000000000000000;
	sram_mem[86389] = 16'b0000000000000000;
	sram_mem[86390] = 16'b0000000000000000;
	sram_mem[86391] = 16'b0000000000000000;
	sram_mem[86392] = 16'b0000000000000000;
	sram_mem[86393] = 16'b0000000000000000;
	sram_mem[86394] = 16'b0000000000000000;
	sram_mem[86395] = 16'b0000000000000000;
	sram_mem[86396] = 16'b0000000000000000;
	sram_mem[86397] = 16'b0000000000000000;
	sram_mem[86398] = 16'b0000000000000000;
	sram_mem[86399] = 16'b0000000000000000;
	sram_mem[86400] = 16'b0000000000000000;
	sram_mem[86401] = 16'b0000000000000000;
	sram_mem[86402] = 16'b0000000000000000;
	sram_mem[86403] = 16'b0000000000000000;
	sram_mem[86404] = 16'b0000000000000000;
	sram_mem[86405] = 16'b0000000000000000;
	sram_mem[86406] = 16'b0000000000000000;
	sram_mem[86407] = 16'b0000000000000000;
	sram_mem[86408] = 16'b0000000000000000;
	sram_mem[86409] = 16'b0000000000000000;
	sram_mem[86410] = 16'b0000000000000000;
	sram_mem[86411] = 16'b0000000000000000;
	sram_mem[86412] = 16'b0000000000000000;
	sram_mem[86413] = 16'b0000000000000000;
	sram_mem[86414] = 16'b0000000000000000;
	sram_mem[86415] = 16'b0000000000000000;
	sram_mem[86416] = 16'b0000000000000000;
	sram_mem[86417] = 16'b0000000000000000;
	sram_mem[86418] = 16'b0000000000000000;
	sram_mem[86419] = 16'b0000000000000000;
	sram_mem[86420] = 16'b0000000000000000;
	sram_mem[86421] = 16'b0000000000000000;
	sram_mem[86422] = 16'b0000000000000000;
	sram_mem[86423] = 16'b0000000000000000;
	sram_mem[86424] = 16'b0000000000000000;
	sram_mem[86425] = 16'b0000000000000000;
	sram_mem[86426] = 16'b0000000000000000;
	sram_mem[86427] = 16'b0000000000000000;
	sram_mem[86428] = 16'b0000000000000000;
	sram_mem[86429] = 16'b0000000000000000;
	sram_mem[86430] = 16'b0000000000000000;
	sram_mem[86431] = 16'b0000000000000000;
	sram_mem[86432] = 16'b0000000000000000;
	sram_mem[86433] = 16'b0000000000000000;
	sram_mem[86434] = 16'b0000000000000000;
	sram_mem[86435] = 16'b0000000000000000;
	sram_mem[86436] = 16'b0000000000000000;
	sram_mem[86437] = 16'b0000000000000000;
	sram_mem[86438] = 16'b0000000000000000;
	sram_mem[86439] = 16'b0000000000000000;
	sram_mem[86440] = 16'b0000000000000000;
	sram_mem[86441] = 16'b0000000000000000;
	sram_mem[86442] = 16'b0000000000000000;
	sram_mem[86443] = 16'b0000000000000000;
	sram_mem[86444] = 16'b0000000000000000;
	sram_mem[86445] = 16'b0000000000000000;
	sram_mem[86446] = 16'b0000000000000000;
	sram_mem[86447] = 16'b0000000000000000;
	sram_mem[86448] = 16'b0000000000000000;
	sram_mem[86449] = 16'b0000000000000000;
	sram_mem[86450] = 16'b0000000000000000;
	sram_mem[86451] = 16'b0000000000000000;
	sram_mem[86452] = 16'b0000000000000000;
	sram_mem[86453] = 16'b0000000000000000;
	sram_mem[86454] = 16'b0000000000000000;
	sram_mem[86455] = 16'b0000000000000000;
	sram_mem[86456] = 16'b0000000000000000;
	sram_mem[86457] = 16'b0000000000000000;
	sram_mem[86458] = 16'b0000000000000000;
	sram_mem[86459] = 16'b0000000000000000;
	sram_mem[86460] = 16'b0000000000000000;
	sram_mem[86461] = 16'b0000000000000000;
	sram_mem[86462] = 16'b0000000000000000;
	sram_mem[86463] = 16'b0000000000000000;
	sram_mem[86464] = 16'b0000000000000000;
	sram_mem[86465] = 16'b0000000000000000;
	sram_mem[86466] = 16'b0000000000000000;
	sram_mem[86467] = 16'b0000000000000000;
	sram_mem[86468] = 16'b0000000000000000;
	sram_mem[86469] = 16'b0000000000000000;
	sram_mem[86470] = 16'b0000000000000000;
	sram_mem[86471] = 16'b0000000000000000;
	sram_mem[86472] = 16'b0000000000000000;
	sram_mem[86473] = 16'b0000000000000000;
	sram_mem[86474] = 16'b0000000000000000;
	sram_mem[86475] = 16'b0000000000000000;
	sram_mem[86476] = 16'b0000000000000000;
	sram_mem[86477] = 16'b0000000000000000;
	sram_mem[86478] = 16'b0000000000000000;
	sram_mem[86479] = 16'b0000000000000000;
	sram_mem[86480] = 16'b0000000000000000;
	sram_mem[86481] = 16'b0000000000000000;
	sram_mem[86482] = 16'b0000000000000000;
	sram_mem[86483] = 16'b0000000000000000;
	sram_mem[86484] = 16'b0000000000000000;
	sram_mem[86485] = 16'b0000000000000000;
	sram_mem[86486] = 16'b0000000000000000;
	sram_mem[86487] = 16'b0000000000000000;
	sram_mem[86488] = 16'b0000000000000000;
	sram_mem[86489] = 16'b0000000000000000;
	sram_mem[86490] = 16'b0000000000000000;
	sram_mem[86491] = 16'b0000000000000000;
	sram_mem[86492] = 16'b0000000000000000;
	sram_mem[86493] = 16'b0000000000000000;
	sram_mem[86494] = 16'b0000000000000000;
	sram_mem[86495] = 16'b0000000000000000;
	sram_mem[86496] = 16'b0000000000000000;
	sram_mem[86497] = 16'b0000000000000000;
	sram_mem[86498] = 16'b0000000000000000;
	sram_mem[86499] = 16'b0000000000000000;
	sram_mem[86500] = 16'b0000000000000000;
	sram_mem[86501] = 16'b0000000000000000;
	sram_mem[86502] = 16'b0000000000000000;
	sram_mem[86503] = 16'b0000000000000000;
	sram_mem[86504] = 16'b0000000000000000;
	sram_mem[86505] = 16'b0000000000000000;
	sram_mem[86506] = 16'b0000000000000000;
	sram_mem[86507] = 16'b0000000000000000;
	sram_mem[86508] = 16'b0000000000000000;
	sram_mem[86509] = 16'b0000000000000000;
	sram_mem[86510] = 16'b0000000000000000;
	sram_mem[86511] = 16'b0000000000000000;
	sram_mem[86512] = 16'b0000000000000000;
	sram_mem[86513] = 16'b0000000000000000;
	sram_mem[86514] = 16'b0000000000000000;
	sram_mem[86515] = 16'b0000000000000000;
	sram_mem[86516] = 16'b0000000000000000;
	sram_mem[86517] = 16'b0000000000000000;
	sram_mem[86518] = 16'b0000000000000000;
	sram_mem[86519] = 16'b0000000000000000;
	sram_mem[86520] = 16'b0000000000000000;
	sram_mem[86521] = 16'b0000000000000000;
	sram_mem[86522] = 16'b0000000000000000;
	sram_mem[86523] = 16'b0000000000000000;
	sram_mem[86524] = 16'b0000000000000000;
	sram_mem[86525] = 16'b0000000000000000;
	sram_mem[86526] = 16'b0000000000000000;
	sram_mem[86527] = 16'b0000000000000000;
	sram_mem[86528] = 16'b0000000000000000;
	sram_mem[86529] = 16'b0000000000000000;
	sram_mem[86530] = 16'b0000000000000000;
	sram_mem[86531] = 16'b0000000000000000;
	sram_mem[86532] = 16'b0000000000000000;
	sram_mem[86533] = 16'b0000000000000000;
	sram_mem[86534] = 16'b0000000000000000;
	sram_mem[86535] = 16'b0000000000000000;
	sram_mem[86536] = 16'b0000000000000000;
	sram_mem[86537] = 16'b0000000000000000;
	sram_mem[86538] = 16'b0000000000000000;
	sram_mem[86539] = 16'b0000000000000000;
	sram_mem[86540] = 16'b0000000000000000;
	sram_mem[86541] = 16'b0000000000000000;
	sram_mem[86542] = 16'b0000000000000000;
	sram_mem[86543] = 16'b0000000000000000;
	sram_mem[86544] = 16'b0000000000000000;
	sram_mem[86545] = 16'b0000000000000000;
	sram_mem[86546] = 16'b0000000000000000;
	sram_mem[86547] = 16'b0000000000000000;
	sram_mem[86548] = 16'b0000000000000000;
	sram_mem[86549] = 16'b0000000000000000;
	sram_mem[86550] = 16'b0000000000000000;
	sram_mem[86551] = 16'b0000000000000000;
	sram_mem[86552] = 16'b0000000000000000;
	sram_mem[86553] = 16'b0000000000000000;
	sram_mem[86554] = 16'b0000000000000000;
	sram_mem[86555] = 16'b0000000000000000;
	sram_mem[86556] = 16'b0000000000000000;
	sram_mem[86557] = 16'b0000000000000000;
	sram_mem[86558] = 16'b0000000000000000;
	sram_mem[86559] = 16'b0000000000000000;
	sram_mem[86560] = 16'b0000000000000000;
	sram_mem[86561] = 16'b0000000000000000;
	sram_mem[86562] = 16'b0000000000000000;
	sram_mem[86563] = 16'b0000000000000000;
	sram_mem[86564] = 16'b0000000000000000;
	sram_mem[86565] = 16'b0000000000000000;
	sram_mem[86566] = 16'b0000000000000000;
	sram_mem[86567] = 16'b0000000000000000;
	sram_mem[86568] = 16'b0000000000000000;
	sram_mem[86569] = 16'b0000000000000000;
	sram_mem[86570] = 16'b0000000000000000;
	sram_mem[86571] = 16'b0000000000000000;
	sram_mem[86572] = 16'b0000000000000000;
	sram_mem[86573] = 16'b0000000000000000;
	sram_mem[86574] = 16'b0000000000000000;
	sram_mem[86575] = 16'b0000000000000000;
	sram_mem[86576] = 16'b0000000000000000;
	sram_mem[86577] = 16'b0000000000000000;
	sram_mem[86578] = 16'b0000000000000000;
	sram_mem[86579] = 16'b0000000000000000;
	sram_mem[86580] = 16'b0000000000000000;
	sram_mem[86581] = 16'b0000000000000000;
	sram_mem[86582] = 16'b0000000000000000;
	sram_mem[86583] = 16'b0000000000000000;
	sram_mem[86584] = 16'b0000000000000000;
	sram_mem[86585] = 16'b0000000000000000;
	sram_mem[86586] = 16'b0000000000000000;
	sram_mem[86587] = 16'b0000000000000000;
	sram_mem[86588] = 16'b0000000000000000;
	sram_mem[86589] = 16'b0000000000000000;
	sram_mem[86590] = 16'b0000000000000000;
	sram_mem[86591] = 16'b0000000000000000;
	sram_mem[86592] = 16'b0000000000000000;
	sram_mem[86593] = 16'b0000000000000000;
	sram_mem[86594] = 16'b0000000000000000;
	sram_mem[86595] = 16'b0000000000000000;
	sram_mem[86596] = 16'b0000000000000000;
	sram_mem[86597] = 16'b0000000000000000;
	sram_mem[86598] = 16'b0000000000000000;
	sram_mem[86599] = 16'b0000000000000000;
	sram_mem[86600] = 16'b0000000000000000;
	sram_mem[86601] = 16'b0000000000000000;
	sram_mem[86602] = 16'b0000000000000000;
	sram_mem[86603] = 16'b0000000000000000;
	sram_mem[86604] = 16'b0000000000000000;
	sram_mem[86605] = 16'b0000000000000000;
	sram_mem[86606] = 16'b0000000000000000;
	sram_mem[86607] = 16'b0000000000000000;
	sram_mem[86608] = 16'b0000000000000000;
	sram_mem[86609] = 16'b0000000000000000;
	sram_mem[86610] = 16'b0000000000000000;
	sram_mem[86611] = 16'b0000000000000000;
	sram_mem[86612] = 16'b0000000000000000;
	sram_mem[86613] = 16'b0000000000000000;
	sram_mem[86614] = 16'b0000000000000000;
	sram_mem[86615] = 16'b0000000000000000;
	sram_mem[86616] = 16'b0000000000000000;
	sram_mem[86617] = 16'b0000000000000000;
	sram_mem[86618] = 16'b0000000000000000;
	sram_mem[86619] = 16'b0000000000000000;
	sram_mem[86620] = 16'b0000000000000000;
	sram_mem[86621] = 16'b0000000000000000;
	sram_mem[86622] = 16'b0000000000000000;
	sram_mem[86623] = 16'b0000000000000000;
	sram_mem[86624] = 16'b0000000000000000;
	sram_mem[86625] = 16'b0000000000000000;
	sram_mem[86626] = 16'b0000000000000000;
	sram_mem[86627] = 16'b0000000000000000;
	sram_mem[86628] = 16'b0000000000000000;
	sram_mem[86629] = 16'b0000000000000000;
	sram_mem[86630] = 16'b0000000000000000;
	sram_mem[86631] = 16'b0000000000000000;
	sram_mem[86632] = 16'b0000000000000000;
	sram_mem[86633] = 16'b0000000000000000;
	sram_mem[86634] = 16'b0000000000000000;
	sram_mem[86635] = 16'b0000000000000000;
	sram_mem[86636] = 16'b0000000000000000;
	sram_mem[86637] = 16'b0000000000000000;
	sram_mem[86638] = 16'b0000000000000000;
	sram_mem[86639] = 16'b0000000000000000;
	sram_mem[86640] = 16'b0000000000000000;
	sram_mem[86641] = 16'b0000000000000000;
	sram_mem[86642] = 16'b0000000000000000;
	sram_mem[86643] = 16'b0000000000000000;
	sram_mem[86644] = 16'b0000000000000000;
	sram_mem[86645] = 16'b0000000000000000;
	sram_mem[86646] = 16'b0000000000000000;
	sram_mem[86647] = 16'b0000000000000000;
	sram_mem[86648] = 16'b0000000000000000;
	sram_mem[86649] = 16'b0000000000000000;
	sram_mem[86650] = 16'b0000000000000000;
	sram_mem[86651] = 16'b0000000000000000;
	sram_mem[86652] = 16'b0000000000000000;
	sram_mem[86653] = 16'b0000000000000000;
	sram_mem[86654] = 16'b0000000000000000;
	sram_mem[86655] = 16'b0000000000000000;
	sram_mem[86656] = 16'b0000000000000000;
	sram_mem[86657] = 16'b0000000000000000;
	sram_mem[86658] = 16'b0000000000000000;
	sram_mem[86659] = 16'b0000000000000000;
	sram_mem[86660] = 16'b0000000000000000;
	sram_mem[86661] = 16'b0000000000000000;
	sram_mem[86662] = 16'b0000000000000000;
	sram_mem[86663] = 16'b0000000000000000;
	sram_mem[86664] = 16'b0000000000000000;
	sram_mem[86665] = 16'b0000000000000000;
	sram_mem[86666] = 16'b0000000000000000;
	sram_mem[86667] = 16'b0000000000000000;
	sram_mem[86668] = 16'b0000000000000000;
	sram_mem[86669] = 16'b0000000000000000;
	sram_mem[86670] = 16'b0000000000000000;
	sram_mem[86671] = 16'b0000000000000000;
	sram_mem[86672] = 16'b0000000000000000;
	sram_mem[86673] = 16'b0000000000000000;
	sram_mem[86674] = 16'b0000000000000000;
	sram_mem[86675] = 16'b0000000000000000;
	sram_mem[86676] = 16'b0000000000000000;
	sram_mem[86677] = 16'b0000000000000000;
	sram_mem[86678] = 16'b0000000000000000;
	sram_mem[86679] = 16'b0000000000000000;
	sram_mem[86680] = 16'b0000000000000000;
	sram_mem[86681] = 16'b0000000000000000;
	sram_mem[86682] = 16'b0000000000000000;
	sram_mem[86683] = 16'b0000000000000000;
	sram_mem[86684] = 16'b0000000000000000;
	sram_mem[86685] = 16'b0000000000000000;
	sram_mem[86686] = 16'b0000000000000000;
	sram_mem[86687] = 16'b0000000000000000;
	sram_mem[86688] = 16'b0000000000000000;
	sram_mem[86689] = 16'b0000000000000000;
	sram_mem[86690] = 16'b0000000000000000;
	sram_mem[86691] = 16'b0000000000000000;
	sram_mem[86692] = 16'b0000000000000000;
	sram_mem[86693] = 16'b0000000000000000;
	sram_mem[86694] = 16'b0000000000000000;
	sram_mem[86695] = 16'b0000000000000000;
	sram_mem[86696] = 16'b0000000000000000;
	sram_mem[86697] = 16'b0000000000000000;
	sram_mem[86698] = 16'b0000000000000000;
	sram_mem[86699] = 16'b0000000000000000;
	sram_mem[86700] = 16'b0000000000000000;
	sram_mem[86701] = 16'b0000000000000000;
	sram_mem[86702] = 16'b0000000000000000;
	sram_mem[86703] = 16'b0000000000000000;
	sram_mem[86704] = 16'b0000000000000000;
	sram_mem[86705] = 16'b0000000000000000;
	sram_mem[86706] = 16'b0000000000000000;
	sram_mem[86707] = 16'b0000000000000000;
	sram_mem[86708] = 16'b0000000000000000;
	sram_mem[86709] = 16'b0000000000000000;
	sram_mem[86710] = 16'b0000000000000000;
	sram_mem[86711] = 16'b0000000000000000;
	sram_mem[86712] = 16'b0000000000000000;
	sram_mem[86713] = 16'b0000000000000000;
	sram_mem[86714] = 16'b0000000000000000;
	sram_mem[86715] = 16'b0000000000000000;
	sram_mem[86716] = 16'b0000000000000000;
	sram_mem[86717] = 16'b0000000000000000;
	sram_mem[86718] = 16'b0000000000000000;
	sram_mem[86719] = 16'b0000000000000000;
	sram_mem[86720] = 16'b0000000000000000;
	sram_mem[86721] = 16'b0000000000000000;
	sram_mem[86722] = 16'b0000000000000000;
	sram_mem[86723] = 16'b0000000000000000;
	sram_mem[86724] = 16'b0000000000000000;
	sram_mem[86725] = 16'b0000000000000000;
	sram_mem[86726] = 16'b0000000000000000;
	sram_mem[86727] = 16'b0000000000000000;
	sram_mem[86728] = 16'b0000000000000000;
	sram_mem[86729] = 16'b0000000000000000;
	sram_mem[86730] = 16'b0000000000000000;
	sram_mem[86731] = 16'b0000000000000000;
	sram_mem[86732] = 16'b0000000000000000;
	sram_mem[86733] = 16'b0000000000000000;
	sram_mem[86734] = 16'b0000000000000000;
	sram_mem[86735] = 16'b0000000000000000;
	sram_mem[86736] = 16'b0000000000000000;
	sram_mem[86737] = 16'b0000000000000000;
	sram_mem[86738] = 16'b0000000000000000;
	sram_mem[86739] = 16'b0000000000000000;
	sram_mem[86740] = 16'b0000000000000000;
	sram_mem[86741] = 16'b0000000000000000;
	sram_mem[86742] = 16'b0000000000000000;
	sram_mem[86743] = 16'b0000000000000000;
	sram_mem[86744] = 16'b0000000000000000;
	sram_mem[86745] = 16'b0000000000000000;
	sram_mem[86746] = 16'b0000000000000000;
	sram_mem[86747] = 16'b0000000000000000;
	sram_mem[86748] = 16'b0000000000000000;
	sram_mem[86749] = 16'b0000000000000000;
	sram_mem[86750] = 16'b0000000000000000;
	sram_mem[86751] = 16'b0000000000000000;
	sram_mem[86752] = 16'b0000000000000000;
	sram_mem[86753] = 16'b0000000000000000;
	sram_mem[86754] = 16'b0000000000000000;
	sram_mem[86755] = 16'b0000000000000000;
	sram_mem[86756] = 16'b0000000000000000;
	sram_mem[86757] = 16'b0000000000000000;
	sram_mem[86758] = 16'b0000000000000000;
	sram_mem[86759] = 16'b0000000000000000;
	sram_mem[86760] = 16'b0000000000000000;
	sram_mem[86761] = 16'b0000000000000000;
	sram_mem[86762] = 16'b0000000000000000;
	sram_mem[86763] = 16'b0000000000000000;
	sram_mem[86764] = 16'b0000000000000000;
	sram_mem[86765] = 16'b0000000000000000;
	sram_mem[86766] = 16'b0000000000000000;
	sram_mem[86767] = 16'b0000000000000000;
	sram_mem[86768] = 16'b0000000000000000;
	sram_mem[86769] = 16'b0000000000000000;
	sram_mem[86770] = 16'b0000000000000000;
	sram_mem[86771] = 16'b0000000000000000;
	sram_mem[86772] = 16'b0000000000000000;
	sram_mem[86773] = 16'b0000000000000000;
	sram_mem[86774] = 16'b0000000000000000;
	sram_mem[86775] = 16'b0000000000000000;
	sram_mem[86776] = 16'b0000000000000000;
	sram_mem[86777] = 16'b0000000000000000;
	sram_mem[86778] = 16'b0000000000000000;
	sram_mem[86779] = 16'b0000000000000000;
	sram_mem[86780] = 16'b0000000000000000;
	sram_mem[86781] = 16'b0000000000000000;
	sram_mem[86782] = 16'b0000000000000000;
	sram_mem[86783] = 16'b0000000000000000;
	sram_mem[86784] = 16'b0000000000000000;
	sram_mem[86785] = 16'b0000000000000000;
	sram_mem[86786] = 16'b0000000000000000;
	sram_mem[86787] = 16'b0000000000000000;
	sram_mem[86788] = 16'b0000000000000000;
	sram_mem[86789] = 16'b0000000000000000;
	sram_mem[86790] = 16'b0000000000000000;
	sram_mem[86791] = 16'b0000000000000000;
	sram_mem[86792] = 16'b0000000000000000;
	sram_mem[86793] = 16'b0000000000000000;
	sram_mem[86794] = 16'b0000000000000000;
	sram_mem[86795] = 16'b0000000000000000;
	sram_mem[86796] = 16'b0000000000000000;
	sram_mem[86797] = 16'b0000000000000000;
	sram_mem[86798] = 16'b0000000000000000;
	sram_mem[86799] = 16'b0000000000000000;
	sram_mem[86800] = 16'b0000000000000000;
	sram_mem[86801] = 16'b0000000000000000;
	sram_mem[86802] = 16'b0000000000000000;
	sram_mem[86803] = 16'b0000000000000000;
	sram_mem[86804] = 16'b0000000000000000;
	sram_mem[86805] = 16'b0000000000000000;
	sram_mem[86806] = 16'b0000000000000000;
	sram_mem[86807] = 16'b0000000000000000;
	sram_mem[86808] = 16'b0000000000000000;
	sram_mem[86809] = 16'b0000000000000000;
	sram_mem[86810] = 16'b0000000000000000;
	sram_mem[86811] = 16'b0000000000000000;
	sram_mem[86812] = 16'b0000000000000000;
	sram_mem[86813] = 16'b0000000000000000;
	sram_mem[86814] = 16'b0000000000000000;
	sram_mem[86815] = 16'b0000000000000000;
	sram_mem[86816] = 16'b0000000000000000;
	sram_mem[86817] = 16'b0000000000000000;
	sram_mem[86818] = 16'b0000000000000000;
	sram_mem[86819] = 16'b0000000000000000;
	sram_mem[86820] = 16'b0000000000000000;
	sram_mem[86821] = 16'b0000000000000000;
	sram_mem[86822] = 16'b0000000000000000;
	sram_mem[86823] = 16'b0000000000000000;
	sram_mem[86824] = 16'b0000000000000000;
	sram_mem[86825] = 16'b0000000000000000;
	sram_mem[86826] = 16'b0000000000000000;
	sram_mem[86827] = 16'b0000000000000000;
	sram_mem[86828] = 16'b0000000000000000;
	sram_mem[86829] = 16'b0000000000000000;
	sram_mem[86830] = 16'b0000000000000000;
	sram_mem[86831] = 16'b0000000000000000;
	sram_mem[86832] = 16'b0000000000000000;
	sram_mem[86833] = 16'b0000000000000000;
	sram_mem[86834] = 16'b0000000000000000;
	sram_mem[86835] = 16'b0000000000000000;
	sram_mem[86836] = 16'b0000000000000000;
	sram_mem[86837] = 16'b0000000000000000;
	sram_mem[86838] = 16'b0000000000000000;
	sram_mem[86839] = 16'b0000000000000000;
	sram_mem[86840] = 16'b0000000000000000;
	sram_mem[86841] = 16'b0000000000000000;
	sram_mem[86842] = 16'b0000000000000000;
	sram_mem[86843] = 16'b0000000000000000;
	sram_mem[86844] = 16'b0000000000000000;
	sram_mem[86845] = 16'b0000000000000000;
	sram_mem[86846] = 16'b0000000000000000;
	sram_mem[86847] = 16'b0000000000000000;
	sram_mem[86848] = 16'b0000000000000000;
	sram_mem[86849] = 16'b0000000000000000;
	sram_mem[86850] = 16'b0000000000000000;
	sram_mem[86851] = 16'b0000000000000000;
	sram_mem[86852] = 16'b0000000000000000;
	sram_mem[86853] = 16'b0000000000000000;
	sram_mem[86854] = 16'b0000000000000000;
	sram_mem[86855] = 16'b0000000000000000;
	sram_mem[86856] = 16'b0000000000000000;
	sram_mem[86857] = 16'b0000000000000000;
	sram_mem[86858] = 16'b0000000000000000;
	sram_mem[86859] = 16'b0000000000000000;
	sram_mem[86860] = 16'b0000000000000000;
	sram_mem[86861] = 16'b0000000000000000;
	sram_mem[86862] = 16'b0000000000000000;
	sram_mem[86863] = 16'b0000000000000000;
	sram_mem[86864] = 16'b0000000000000000;
	sram_mem[86865] = 16'b0000000000000000;
	sram_mem[86866] = 16'b0000000000000000;
	sram_mem[86867] = 16'b0000000000000000;
	sram_mem[86868] = 16'b0000000000000000;
	sram_mem[86869] = 16'b0000000000000000;
	sram_mem[86870] = 16'b0000000000000000;
	sram_mem[86871] = 16'b0000000000000000;
	sram_mem[86872] = 16'b0000000000000000;
	sram_mem[86873] = 16'b0000000000000000;
	sram_mem[86874] = 16'b0000000000000000;
	sram_mem[86875] = 16'b0000000000000000;
	sram_mem[86876] = 16'b0000000000000000;
	sram_mem[86877] = 16'b0000000000000000;
	sram_mem[86878] = 16'b0000000000000000;
	sram_mem[86879] = 16'b0000000000000000;
	sram_mem[86880] = 16'b0000000000000000;
	sram_mem[86881] = 16'b0000000000000000;
	sram_mem[86882] = 16'b0000000000000000;
	sram_mem[86883] = 16'b0000000000000000;
	sram_mem[86884] = 16'b0000000000000000;
	sram_mem[86885] = 16'b0000000000000000;
	sram_mem[86886] = 16'b0000000000000000;
	sram_mem[86887] = 16'b0000000000000000;
	sram_mem[86888] = 16'b0000000000000000;
	sram_mem[86889] = 16'b0000000000000000;
	sram_mem[86890] = 16'b0000000000000000;
	sram_mem[86891] = 16'b0000000000000000;
	sram_mem[86892] = 16'b0000000000000000;
	sram_mem[86893] = 16'b0000000000000000;
	sram_mem[86894] = 16'b0000000000000000;
	sram_mem[86895] = 16'b0000000000000000;
	sram_mem[86896] = 16'b0000000000000000;
	sram_mem[86897] = 16'b0000000000000000;
	sram_mem[86898] = 16'b0000000000000000;
	sram_mem[86899] = 16'b0000000000000000;
	sram_mem[86900] = 16'b0000000000000000;
	sram_mem[86901] = 16'b0000000000000000;
	sram_mem[86902] = 16'b0000000000000000;
	sram_mem[86903] = 16'b0000000000000000;
	sram_mem[86904] = 16'b0000000000000000;
	sram_mem[86905] = 16'b0000000000000000;
	sram_mem[86906] = 16'b0000000000000000;
	sram_mem[86907] = 16'b0000000000000000;
	sram_mem[86908] = 16'b0000000000000000;
	sram_mem[86909] = 16'b0000000000000000;
	sram_mem[86910] = 16'b0000000000000000;
	sram_mem[86911] = 16'b0000000000000000;
	sram_mem[86912] = 16'b0000000000000000;
	sram_mem[86913] = 16'b0000000000000000;
	sram_mem[86914] = 16'b0000000000000000;
	sram_mem[86915] = 16'b0000000000000000;
	sram_mem[86916] = 16'b0000000000000000;
	sram_mem[86917] = 16'b0000000000000000;
	sram_mem[86918] = 16'b0000000000000000;
	sram_mem[86919] = 16'b0000000000000000;
	sram_mem[86920] = 16'b0000000000000000;
	sram_mem[86921] = 16'b0000000000000000;
	sram_mem[86922] = 16'b0000000000000000;
	sram_mem[86923] = 16'b0000000000000000;
	sram_mem[86924] = 16'b0000000000000000;
	sram_mem[86925] = 16'b0000000000000000;
	sram_mem[86926] = 16'b0000000000000000;
	sram_mem[86927] = 16'b0000000000000000;
	sram_mem[86928] = 16'b0000000000000000;
	sram_mem[86929] = 16'b0000000000000000;
	sram_mem[86930] = 16'b0000000000000000;
	sram_mem[86931] = 16'b0000000000000000;
	sram_mem[86932] = 16'b0000000000000000;
	sram_mem[86933] = 16'b0000000000000000;
	sram_mem[86934] = 16'b0000000000000000;
	sram_mem[86935] = 16'b0000000000000000;
	sram_mem[86936] = 16'b0000000000000000;
	sram_mem[86937] = 16'b0000000000000000;
	sram_mem[86938] = 16'b0000000000000000;
	sram_mem[86939] = 16'b0000000000000000;
	sram_mem[86940] = 16'b0000000000000000;
	sram_mem[86941] = 16'b0000000000000000;
	sram_mem[86942] = 16'b0000000000000000;
	sram_mem[86943] = 16'b0000000000000000;
	sram_mem[86944] = 16'b0000000000000000;
	sram_mem[86945] = 16'b0000000000000000;
	sram_mem[86946] = 16'b0000000000000000;
	sram_mem[86947] = 16'b0000000000000000;
	sram_mem[86948] = 16'b0000000000000000;
	sram_mem[86949] = 16'b0000000000000000;
	sram_mem[86950] = 16'b0000000000000000;
	sram_mem[86951] = 16'b0000000000000000;
	sram_mem[86952] = 16'b0000000000000000;
	sram_mem[86953] = 16'b0000000000000000;
	sram_mem[86954] = 16'b0000000000000000;
	sram_mem[86955] = 16'b0000000000000000;
	sram_mem[86956] = 16'b0000000000000000;
	sram_mem[86957] = 16'b0000000000000000;
	sram_mem[86958] = 16'b0000000000000000;
	sram_mem[86959] = 16'b0000000000000000;
	sram_mem[86960] = 16'b0000000000000000;
	sram_mem[86961] = 16'b0000000000000000;
	sram_mem[86962] = 16'b0000000000000000;
	sram_mem[86963] = 16'b0000000000000000;
	sram_mem[86964] = 16'b0000000000000000;
	sram_mem[86965] = 16'b0000000000000000;
	sram_mem[86966] = 16'b0000000000000000;
	sram_mem[86967] = 16'b0000000000000000;
	sram_mem[86968] = 16'b0000000000000000;
	sram_mem[86969] = 16'b0000000000000000;
	sram_mem[86970] = 16'b0000000000000000;
	sram_mem[86971] = 16'b0000000000000000;
	sram_mem[86972] = 16'b0000000000000000;
	sram_mem[86973] = 16'b0000000000000000;
	sram_mem[86974] = 16'b0000000000000000;
	sram_mem[86975] = 16'b0000000000000000;
	sram_mem[86976] = 16'b0000000000000000;
	sram_mem[86977] = 16'b0000000000000000;
	sram_mem[86978] = 16'b0000000000000000;
	sram_mem[86979] = 16'b0000000000000000;
	sram_mem[86980] = 16'b0000000000000000;
	sram_mem[86981] = 16'b0000000000000000;
	sram_mem[86982] = 16'b0000000000000000;
	sram_mem[86983] = 16'b0000000000000000;
	sram_mem[86984] = 16'b0000000000000000;
	sram_mem[86985] = 16'b0000000000000000;
	sram_mem[86986] = 16'b0000000000000000;
	sram_mem[86987] = 16'b0000000000000000;
	sram_mem[86988] = 16'b0000000000000000;
	sram_mem[86989] = 16'b0000000000000000;
	sram_mem[86990] = 16'b0000000000000000;
	sram_mem[86991] = 16'b0000000000000000;
	sram_mem[86992] = 16'b0000000000000000;
	sram_mem[86993] = 16'b0000000000000000;
	sram_mem[86994] = 16'b0000000000000000;
	sram_mem[86995] = 16'b0000000000000000;
	sram_mem[86996] = 16'b0000000000000000;
	sram_mem[86997] = 16'b0000000000000000;
	sram_mem[86998] = 16'b0000000000000000;
	sram_mem[86999] = 16'b0000000000000000;
	sram_mem[87000] = 16'b0000000000000000;
	sram_mem[87001] = 16'b0000000000000000;
	sram_mem[87002] = 16'b0000000000000000;
	sram_mem[87003] = 16'b0000000000000000;
	sram_mem[87004] = 16'b0000000000000000;
	sram_mem[87005] = 16'b0000000000000000;
	sram_mem[87006] = 16'b0000000000000000;
	sram_mem[87007] = 16'b0000000000000000;
	sram_mem[87008] = 16'b0000000000000000;
	sram_mem[87009] = 16'b0000000000000000;
	sram_mem[87010] = 16'b0000000000000000;
	sram_mem[87011] = 16'b0000000000000000;
	sram_mem[87012] = 16'b0000000000000000;
	sram_mem[87013] = 16'b0000000000000000;
	sram_mem[87014] = 16'b0000000000000000;
	sram_mem[87015] = 16'b0000000000000000;
	sram_mem[87016] = 16'b0000000000000000;
	sram_mem[87017] = 16'b0000000000000000;
	sram_mem[87018] = 16'b0000000000000000;
	sram_mem[87019] = 16'b0000000000000000;
	sram_mem[87020] = 16'b0000000000000000;
	sram_mem[87021] = 16'b0000000000000000;
	sram_mem[87022] = 16'b0000000000000000;
	sram_mem[87023] = 16'b0000000000000000;
	sram_mem[87024] = 16'b0000000000000000;
	sram_mem[87025] = 16'b0000000000000000;
	sram_mem[87026] = 16'b0000000000000000;
	sram_mem[87027] = 16'b0000000000000000;
	sram_mem[87028] = 16'b0000000000000000;
	sram_mem[87029] = 16'b0000000000000000;
	sram_mem[87030] = 16'b0000000000000000;
	sram_mem[87031] = 16'b0000000000000000;
	sram_mem[87032] = 16'b0000000000000000;
	sram_mem[87033] = 16'b0000000000000000;
	sram_mem[87034] = 16'b0000000000000000;
	sram_mem[87035] = 16'b0000000000000000;
	sram_mem[87036] = 16'b0000000000000000;
	sram_mem[87037] = 16'b0000000000000000;
	sram_mem[87038] = 16'b0000000000000000;
	sram_mem[87039] = 16'b0000000000000000;
	sram_mem[87040] = 16'b0000000000000000;
	sram_mem[87041] = 16'b0000000000000000;
	sram_mem[87042] = 16'b0000000000000000;
	sram_mem[87043] = 16'b0000000000000000;
	sram_mem[87044] = 16'b0000000000000000;
	sram_mem[87045] = 16'b0000000000000000;
	sram_mem[87046] = 16'b0000000000000000;
	sram_mem[87047] = 16'b0000000000000000;
	sram_mem[87048] = 16'b0000000000000000;
	sram_mem[87049] = 16'b0000000000000000;
	sram_mem[87050] = 16'b0000000000000000;
	sram_mem[87051] = 16'b0000000000000000;
	sram_mem[87052] = 16'b0000000000000000;
	sram_mem[87053] = 16'b0000000000000000;
	sram_mem[87054] = 16'b0000000000000000;
	sram_mem[87055] = 16'b0000000000000000;
	sram_mem[87056] = 16'b0000000000000000;
	sram_mem[87057] = 16'b0000000000000000;
	sram_mem[87058] = 16'b0000000000000000;
	sram_mem[87059] = 16'b0000000000000000;
	sram_mem[87060] = 16'b0000000000000000;
	sram_mem[87061] = 16'b0000000000000000;
	sram_mem[87062] = 16'b0000000000000000;
	sram_mem[87063] = 16'b0000000000000000;
	sram_mem[87064] = 16'b0000000000000000;
	sram_mem[87065] = 16'b0000000000000000;
	sram_mem[87066] = 16'b0000000000000000;
	sram_mem[87067] = 16'b0000000000000000;
	sram_mem[87068] = 16'b0000000000000000;
	sram_mem[87069] = 16'b0000000000000000;
	sram_mem[87070] = 16'b0000000000000000;
	sram_mem[87071] = 16'b0000000000000000;
	sram_mem[87072] = 16'b0000000000000000;
	sram_mem[87073] = 16'b0000000000000000;
	sram_mem[87074] = 16'b0000000000000000;
	sram_mem[87075] = 16'b0000000000000000;
	sram_mem[87076] = 16'b0000000000000000;
	sram_mem[87077] = 16'b0000000000000000;
	sram_mem[87078] = 16'b0000000000000000;
	sram_mem[87079] = 16'b0000000000000000;
	sram_mem[87080] = 16'b0000000000000000;
	sram_mem[87081] = 16'b0000000000000000;
	sram_mem[87082] = 16'b0000000000000000;
	sram_mem[87083] = 16'b0000000000000000;
	sram_mem[87084] = 16'b0000000000000000;
	sram_mem[87085] = 16'b0000000000000000;
	sram_mem[87086] = 16'b0000000000000000;
	sram_mem[87087] = 16'b0000000000000000;
	sram_mem[87088] = 16'b0000000000000000;
	sram_mem[87089] = 16'b0000000000000000;
	sram_mem[87090] = 16'b0000000000000000;
	sram_mem[87091] = 16'b0000000000000000;
	sram_mem[87092] = 16'b0000000000000000;
	sram_mem[87093] = 16'b0000000000000000;
	sram_mem[87094] = 16'b0000000000000000;
	sram_mem[87095] = 16'b0000000000000000;
	sram_mem[87096] = 16'b0000000000000000;
	sram_mem[87097] = 16'b0000000000000000;
	sram_mem[87098] = 16'b0000000000000000;
	sram_mem[87099] = 16'b0000000000000000;
	sram_mem[87100] = 16'b0000000000000000;
	sram_mem[87101] = 16'b0000000000000000;
	sram_mem[87102] = 16'b0000000000000000;
	sram_mem[87103] = 16'b0000000000000000;
	sram_mem[87104] = 16'b0000000000000000;
	sram_mem[87105] = 16'b0000000000000000;
	sram_mem[87106] = 16'b0000000000000000;
	sram_mem[87107] = 16'b0000000000000000;
	sram_mem[87108] = 16'b0000000000000000;
	sram_mem[87109] = 16'b0000000000000000;
	sram_mem[87110] = 16'b0000000000000000;
	sram_mem[87111] = 16'b0000000000000000;
	sram_mem[87112] = 16'b0000000000000000;
	sram_mem[87113] = 16'b0000000000000000;
	sram_mem[87114] = 16'b0000000000000000;
	sram_mem[87115] = 16'b0000000000000000;
	sram_mem[87116] = 16'b0000000000000000;
	sram_mem[87117] = 16'b0000000000000000;
	sram_mem[87118] = 16'b0000000000000000;
	sram_mem[87119] = 16'b0000000000000000;
	sram_mem[87120] = 16'b0000000000000000;
	sram_mem[87121] = 16'b0000000000000000;
	sram_mem[87122] = 16'b0000000000000000;
	sram_mem[87123] = 16'b0000000000000000;
	sram_mem[87124] = 16'b0000000000000000;
	sram_mem[87125] = 16'b0000000000000000;
	sram_mem[87126] = 16'b0000000000000000;
	sram_mem[87127] = 16'b0000000000000000;
	sram_mem[87128] = 16'b0000000000000000;
	sram_mem[87129] = 16'b0000000000000000;
	sram_mem[87130] = 16'b0000000000000000;
	sram_mem[87131] = 16'b0000000000000000;
	sram_mem[87132] = 16'b0000000000000000;
	sram_mem[87133] = 16'b0000000000000000;
	sram_mem[87134] = 16'b0000000000000000;
	sram_mem[87135] = 16'b0000000000000000;
	sram_mem[87136] = 16'b0000000000000000;
	sram_mem[87137] = 16'b0000000000000000;
	sram_mem[87138] = 16'b0000000000000000;
	sram_mem[87139] = 16'b0000000000000000;
	sram_mem[87140] = 16'b0000000000000000;
	sram_mem[87141] = 16'b0000000000000000;
	sram_mem[87142] = 16'b0000000000000000;
	sram_mem[87143] = 16'b0000000000000000;
	sram_mem[87144] = 16'b0000000000000000;
	sram_mem[87145] = 16'b0000000000000000;
	sram_mem[87146] = 16'b0000000000000000;
	sram_mem[87147] = 16'b0000000000000000;
	sram_mem[87148] = 16'b0000000000000000;
	sram_mem[87149] = 16'b0000000000000000;
	sram_mem[87150] = 16'b0000000000000000;
	sram_mem[87151] = 16'b0000000000000000;
	sram_mem[87152] = 16'b0000000000000000;
	sram_mem[87153] = 16'b0000000000000000;
	sram_mem[87154] = 16'b0000000000000000;
	sram_mem[87155] = 16'b0000000000000000;
	sram_mem[87156] = 16'b0000000000000000;
	sram_mem[87157] = 16'b0000000000000000;
	sram_mem[87158] = 16'b0000000000000000;
	sram_mem[87159] = 16'b0000000000000000;
	sram_mem[87160] = 16'b0000000000000000;
	sram_mem[87161] = 16'b0000000000000000;
	sram_mem[87162] = 16'b0000000000000000;
	sram_mem[87163] = 16'b0000000000000000;
	sram_mem[87164] = 16'b0000000000000000;
	sram_mem[87165] = 16'b0000000000000000;
	sram_mem[87166] = 16'b0000000000000000;
	sram_mem[87167] = 16'b0000000000000000;
	sram_mem[87168] = 16'b0000000000000000;
	sram_mem[87169] = 16'b0000000000000000;
	sram_mem[87170] = 16'b0000000000000000;
	sram_mem[87171] = 16'b0000000000000000;
	sram_mem[87172] = 16'b0000000000000000;
	sram_mem[87173] = 16'b0000000000000000;
	sram_mem[87174] = 16'b0000000000000000;
	sram_mem[87175] = 16'b0000000000000000;
	sram_mem[87176] = 16'b0000000000000000;
	sram_mem[87177] = 16'b0000000000000000;
	sram_mem[87178] = 16'b0000000000000000;
	sram_mem[87179] = 16'b0000000000000000;
	sram_mem[87180] = 16'b0000000000000000;
	sram_mem[87181] = 16'b0000000000000000;
	sram_mem[87182] = 16'b0000000000000000;
	sram_mem[87183] = 16'b0000000000000000;
	sram_mem[87184] = 16'b0000000000000000;
	sram_mem[87185] = 16'b0000000000000000;
	sram_mem[87186] = 16'b0000000000000000;
	sram_mem[87187] = 16'b0000000000000000;
	sram_mem[87188] = 16'b0000000000000000;
	sram_mem[87189] = 16'b0000000000000000;
	sram_mem[87190] = 16'b0000000000000000;
	sram_mem[87191] = 16'b0000000000000000;
	sram_mem[87192] = 16'b0000000000000000;
	sram_mem[87193] = 16'b0000000000000000;
	sram_mem[87194] = 16'b0000000000000000;
	sram_mem[87195] = 16'b0000000000000000;
	sram_mem[87196] = 16'b0000000000000000;
	sram_mem[87197] = 16'b0000000000000000;
	sram_mem[87198] = 16'b0000000000000000;
	sram_mem[87199] = 16'b0000000000000000;
	sram_mem[87200] = 16'b0000000000000000;
	sram_mem[87201] = 16'b0000000000000000;
	sram_mem[87202] = 16'b0000000000000000;
	sram_mem[87203] = 16'b0000000000000000;
	sram_mem[87204] = 16'b0000000000000000;
	sram_mem[87205] = 16'b0000000000000000;
	sram_mem[87206] = 16'b0000000000000000;
	sram_mem[87207] = 16'b0000000000000000;
	sram_mem[87208] = 16'b0000000000000000;
	sram_mem[87209] = 16'b0000000000000000;
	sram_mem[87210] = 16'b0000000000000000;
	sram_mem[87211] = 16'b0000000000000000;
	sram_mem[87212] = 16'b0000000000000000;
	sram_mem[87213] = 16'b0000000000000000;
	sram_mem[87214] = 16'b0000000000000000;
	sram_mem[87215] = 16'b0000000000000000;
	sram_mem[87216] = 16'b0000000000000000;
	sram_mem[87217] = 16'b0000000000000000;
	sram_mem[87218] = 16'b0000000000000000;
	sram_mem[87219] = 16'b0000000000000000;
	sram_mem[87220] = 16'b0000000000000000;
	sram_mem[87221] = 16'b0000000000000000;
	sram_mem[87222] = 16'b0000000000000000;
	sram_mem[87223] = 16'b0000000000000000;
	sram_mem[87224] = 16'b0000000000000000;
	sram_mem[87225] = 16'b0000000000000000;
	sram_mem[87226] = 16'b0000000000000000;
	sram_mem[87227] = 16'b0000000000000000;
	sram_mem[87228] = 16'b0000000000000000;
	sram_mem[87229] = 16'b0000000000000000;
	sram_mem[87230] = 16'b0000000000000000;
	sram_mem[87231] = 16'b0000000000000000;
	sram_mem[87232] = 16'b0000000000000000;
	sram_mem[87233] = 16'b0000000000000000;
	sram_mem[87234] = 16'b0000000000000000;
	sram_mem[87235] = 16'b0000000000000000;
	sram_mem[87236] = 16'b0000000000000000;
	sram_mem[87237] = 16'b0000000000000000;
	sram_mem[87238] = 16'b0000000000000000;
	sram_mem[87239] = 16'b0000000000000000;
	sram_mem[87240] = 16'b0000000000000000;
	sram_mem[87241] = 16'b0000000000000000;
	sram_mem[87242] = 16'b0000000000000000;
	sram_mem[87243] = 16'b0000000000000000;
	sram_mem[87244] = 16'b0000000000000000;
	sram_mem[87245] = 16'b0000000000000000;
	sram_mem[87246] = 16'b0000000000000000;
	sram_mem[87247] = 16'b0000000000000000;
	sram_mem[87248] = 16'b0000000000000000;
	sram_mem[87249] = 16'b0000000000000000;
	sram_mem[87250] = 16'b0000000000000000;
	sram_mem[87251] = 16'b0000000000000000;
	sram_mem[87252] = 16'b0000000000000000;
	sram_mem[87253] = 16'b0000000000000000;
	sram_mem[87254] = 16'b0000000000000000;
	sram_mem[87255] = 16'b0000000000000000;
	sram_mem[87256] = 16'b0000000000000000;
	sram_mem[87257] = 16'b0000000000000000;
	sram_mem[87258] = 16'b0000000000000000;
	sram_mem[87259] = 16'b0000000000000000;
	sram_mem[87260] = 16'b0000000000000000;
	sram_mem[87261] = 16'b0000000000000000;
	sram_mem[87262] = 16'b0000000000000000;
	sram_mem[87263] = 16'b0000000000000000;
	sram_mem[87264] = 16'b0000000000000000;
	sram_mem[87265] = 16'b0000000000000000;
	sram_mem[87266] = 16'b0000000000000000;
	sram_mem[87267] = 16'b0000000000000000;
	sram_mem[87268] = 16'b0000000000000000;
	sram_mem[87269] = 16'b0000000000000000;
	sram_mem[87270] = 16'b0000000000000000;
	sram_mem[87271] = 16'b0000000000000000;
	sram_mem[87272] = 16'b0000000000000000;
	sram_mem[87273] = 16'b0000000000000000;
	sram_mem[87274] = 16'b0000000000000000;
	sram_mem[87275] = 16'b0000000000000000;
	sram_mem[87276] = 16'b0000000000000000;
	sram_mem[87277] = 16'b0000000000000000;
	sram_mem[87278] = 16'b0000000000000000;
	sram_mem[87279] = 16'b0000000000000000;
	sram_mem[87280] = 16'b0000000000000000;
	sram_mem[87281] = 16'b0000000000000000;
	sram_mem[87282] = 16'b0000000000000000;
	sram_mem[87283] = 16'b0000000000000000;
	sram_mem[87284] = 16'b0000000000000000;
	sram_mem[87285] = 16'b0000000000000000;
	sram_mem[87286] = 16'b0000000000000000;
	sram_mem[87287] = 16'b0000000000000000;
	sram_mem[87288] = 16'b0000000000000000;
	sram_mem[87289] = 16'b0000000000000000;
	sram_mem[87290] = 16'b0000000000000000;
	sram_mem[87291] = 16'b0000000000000000;
	sram_mem[87292] = 16'b0000000000000000;
	sram_mem[87293] = 16'b0000000000000000;
	sram_mem[87294] = 16'b0000000000000000;
	sram_mem[87295] = 16'b0000000000000000;
	sram_mem[87296] = 16'b0000000000000000;
	sram_mem[87297] = 16'b0000000000000000;
	sram_mem[87298] = 16'b0000000000000000;
	sram_mem[87299] = 16'b0000000000000000;
	sram_mem[87300] = 16'b0000000000000000;
	sram_mem[87301] = 16'b0000000000000000;
	sram_mem[87302] = 16'b0000000000000000;
	sram_mem[87303] = 16'b0000000000000000;
	sram_mem[87304] = 16'b0000000000000000;
	sram_mem[87305] = 16'b0000000000000000;
	sram_mem[87306] = 16'b0000000000000000;
	sram_mem[87307] = 16'b0000000000000000;
	sram_mem[87308] = 16'b0000000000000000;
	sram_mem[87309] = 16'b0000000000000000;
	sram_mem[87310] = 16'b0000000000000000;
	sram_mem[87311] = 16'b0000000000000000;
	sram_mem[87312] = 16'b0000000000000000;
	sram_mem[87313] = 16'b0000000000000000;
	sram_mem[87314] = 16'b0000000000000000;
	sram_mem[87315] = 16'b0000000000000000;
	sram_mem[87316] = 16'b0000000000000000;
	sram_mem[87317] = 16'b0000000000000000;
	sram_mem[87318] = 16'b0000000000000000;
	sram_mem[87319] = 16'b0000000000000000;
	sram_mem[87320] = 16'b0000000000000000;
	sram_mem[87321] = 16'b0000000000000000;
	sram_mem[87322] = 16'b0000000000000000;
	sram_mem[87323] = 16'b0000000000000000;
	sram_mem[87324] = 16'b0000000000000000;
	sram_mem[87325] = 16'b0000000000000000;
	sram_mem[87326] = 16'b0000000000000000;
	sram_mem[87327] = 16'b0000000000000000;
	sram_mem[87328] = 16'b0000000000000000;
	sram_mem[87329] = 16'b0000000000000000;
	sram_mem[87330] = 16'b0000000000000000;
	sram_mem[87331] = 16'b0000000000000000;
	sram_mem[87332] = 16'b0000000000000000;
	sram_mem[87333] = 16'b0000000000000000;
	sram_mem[87334] = 16'b0000000000000000;
	sram_mem[87335] = 16'b0000000000000000;
	sram_mem[87336] = 16'b0000000000000000;
	sram_mem[87337] = 16'b0000000000000000;
	sram_mem[87338] = 16'b0000000000000000;
	sram_mem[87339] = 16'b0000000000000000;
	sram_mem[87340] = 16'b0000000000000000;
	sram_mem[87341] = 16'b0000000000000000;
	sram_mem[87342] = 16'b0000000000000000;
	sram_mem[87343] = 16'b0000000000000000;
	sram_mem[87344] = 16'b0000000000000000;
	sram_mem[87345] = 16'b0000000000000000;
	sram_mem[87346] = 16'b0000000000000000;
	sram_mem[87347] = 16'b0000000000000000;
	sram_mem[87348] = 16'b0000000000000000;
	sram_mem[87349] = 16'b0000000000000000;
	sram_mem[87350] = 16'b0000000000000000;
	sram_mem[87351] = 16'b0000000000000000;
	sram_mem[87352] = 16'b0000000000000000;
	sram_mem[87353] = 16'b0000000000000000;
	sram_mem[87354] = 16'b0000000000000000;
	sram_mem[87355] = 16'b0000000000000000;
	sram_mem[87356] = 16'b0000000000000000;
	sram_mem[87357] = 16'b0000000000000000;
	sram_mem[87358] = 16'b0000000000000000;
	sram_mem[87359] = 16'b0000000000000000;
	sram_mem[87360] = 16'b0000000000000000;
	sram_mem[87361] = 16'b0000000000000000;
	sram_mem[87362] = 16'b0000000000000000;
	sram_mem[87363] = 16'b0000000000000000;
	sram_mem[87364] = 16'b0000000000000000;
	sram_mem[87365] = 16'b0000000000000000;
	sram_mem[87366] = 16'b0000000000000000;
	sram_mem[87367] = 16'b0000000000000000;
	sram_mem[87368] = 16'b0000000000000000;
	sram_mem[87369] = 16'b0000000000000000;
	sram_mem[87370] = 16'b0000000000000000;
	sram_mem[87371] = 16'b0000000000000000;
	sram_mem[87372] = 16'b0000000000000000;
	sram_mem[87373] = 16'b0000000000000000;
	sram_mem[87374] = 16'b0000000000000000;
	sram_mem[87375] = 16'b0000000000000000;
	sram_mem[87376] = 16'b0000000000000000;
	sram_mem[87377] = 16'b0000000000000000;
	sram_mem[87378] = 16'b0000000000000000;
	sram_mem[87379] = 16'b0000000000000000;
	sram_mem[87380] = 16'b0000000000000000;
	sram_mem[87381] = 16'b0000000000000000;
	sram_mem[87382] = 16'b0000000000000000;
	sram_mem[87383] = 16'b0000000000000000;
	sram_mem[87384] = 16'b0000000000000000;
	sram_mem[87385] = 16'b0000000000000000;
	sram_mem[87386] = 16'b0000000000000000;
	sram_mem[87387] = 16'b0000000000000000;
	sram_mem[87388] = 16'b0000000000000000;
	sram_mem[87389] = 16'b0000000000000000;
	sram_mem[87390] = 16'b0000000000000000;
	sram_mem[87391] = 16'b0000000000000000;
	sram_mem[87392] = 16'b0000000000000000;
	sram_mem[87393] = 16'b0000000000000000;
	sram_mem[87394] = 16'b0000000000000000;
	sram_mem[87395] = 16'b0000000000000000;
	sram_mem[87396] = 16'b0000000000000000;
	sram_mem[87397] = 16'b0000000000000000;
	sram_mem[87398] = 16'b0000000000000000;
	sram_mem[87399] = 16'b0000000000000000;
	sram_mem[87400] = 16'b0000000000000000;
	sram_mem[87401] = 16'b0000000000000000;
	sram_mem[87402] = 16'b0000000000000000;
	sram_mem[87403] = 16'b0000000000000000;
	sram_mem[87404] = 16'b0000000000000000;
	sram_mem[87405] = 16'b0000000000000000;
	sram_mem[87406] = 16'b0000000000000000;
	sram_mem[87407] = 16'b0000000000000000;
	sram_mem[87408] = 16'b0000000000000000;
	sram_mem[87409] = 16'b0000000000000000;
	sram_mem[87410] = 16'b0000000000000000;
	sram_mem[87411] = 16'b0000000000000000;
	sram_mem[87412] = 16'b0000000000000000;
	sram_mem[87413] = 16'b0000000000000000;
	sram_mem[87414] = 16'b0000000000000000;
	sram_mem[87415] = 16'b0000000000000000;
	sram_mem[87416] = 16'b0000000000000000;
	sram_mem[87417] = 16'b0000000000000000;
	sram_mem[87418] = 16'b0000000000000000;
	sram_mem[87419] = 16'b0000000000000000;
	sram_mem[87420] = 16'b0000000000000000;
	sram_mem[87421] = 16'b0000000000000000;
	sram_mem[87422] = 16'b0000000000000000;
	sram_mem[87423] = 16'b0000000000000000;
	sram_mem[87424] = 16'b0000000000000000;
	sram_mem[87425] = 16'b0000000000000000;
	sram_mem[87426] = 16'b0000000000000000;
	sram_mem[87427] = 16'b0000000000000000;
	sram_mem[87428] = 16'b0000000000000000;
	sram_mem[87429] = 16'b0000000000000000;
	sram_mem[87430] = 16'b0000000000000000;
	sram_mem[87431] = 16'b0000000000000000;
	sram_mem[87432] = 16'b0000000000000000;
	sram_mem[87433] = 16'b0000000000000000;
	sram_mem[87434] = 16'b0000000000000000;
	sram_mem[87435] = 16'b0000000000000000;
	sram_mem[87436] = 16'b0000000000000000;
	sram_mem[87437] = 16'b0000000000000000;
	sram_mem[87438] = 16'b0000000000000000;
	sram_mem[87439] = 16'b0000000000000000;
	sram_mem[87440] = 16'b0000000000000000;
	sram_mem[87441] = 16'b0000000000000000;
	sram_mem[87442] = 16'b0000000000000000;
	sram_mem[87443] = 16'b0000000000000000;
	sram_mem[87444] = 16'b0000000000000000;
	sram_mem[87445] = 16'b0000000000000000;
	sram_mem[87446] = 16'b0000000000000000;
	sram_mem[87447] = 16'b0000000000000000;
	sram_mem[87448] = 16'b0000000000000000;
	sram_mem[87449] = 16'b0000000000000000;
	sram_mem[87450] = 16'b0000000000000000;
	sram_mem[87451] = 16'b0000000000000000;
	sram_mem[87452] = 16'b0000000000000000;
	sram_mem[87453] = 16'b0000000000000000;
	sram_mem[87454] = 16'b0000000000000000;
	sram_mem[87455] = 16'b0000000000000000;
	sram_mem[87456] = 16'b0000000000000000;
	sram_mem[87457] = 16'b0000000000000000;
	sram_mem[87458] = 16'b0000000000000000;
	sram_mem[87459] = 16'b0000000000000000;
	sram_mem[87460] = 16'b0000000000000000;
	sram_mem[87461] = 16'b0000000000000000;
	sram_mem[87462] = 16'b0000000000000000;
	sram_mem[87463] = 16'b0000000000000000;
	sram_mem[87464] = 16'b0000000000000000;
	sram_mem[87465] = 16'b0000000000000000;
	sram_mem[87466] = 16'b0000000000000000;
	sram_mem[87467] = 16'b0000000000000000;
	sram_mem[87468] = 16'b0000000000000000;
	sram_mem[87469] = 16'b0000000000000000;
	sram_mem[87470] = 16'b0000000000000000;
	sram_mem[87471] = 16'b0000000000000000;
	sram_mem[87472] = 16'b0000000000000000;
	sram_mem[87473] = 16'b0000000000000000;
	sram_mem[87474] = 16'b0000000000000000;
	sram_mem[87475] = 16'b0000000000000000;
	sram_mem[87476] = 16'b0000000000000000;
	sram_mem[87477] = 16'b0000000000000000;
	sram_mem[87478] = 16'b0000000000000000;
	sram_mem[87479] = 16'b0000000000000000;
	sram_mem[87480] = 16'b0000000000000000;
	sram_mem[87481] = 16'b0000000000000000;
	sram_mem[87482] = 16'b0000000000000000;
	sram_mem[87483] = 16'b0000000000000000;
	sram_mem[87484] = 16'b0000000000000000;
	sram_mem[87485] = 16'b0000000000000000;
	sram_mem[87486] = 16'b0000000000000000;
	sram_mem[87487] = 16'b0000000000000000;
	sram_mem[87488] = 16'b0000000000000000;
	sram_mem[87489] = 16'b0000000000000000;
	sram_mem[87490] = 16'b0000000000000000;
	sram_mem[87491] = 16'b0000000000000000;
	sram_mem[87492] = 16'b0000000000000000;
	sram_mem[87493] = 16'b0000000000000000;
	sram_mem[87494] = 16'b0000000000000000;
	sram_mem[87495] = 16'b0000000000000000;
	sram_mem[87496] = 16'b0000000000000000;
	sram_mem[87497] = 16'b0000000000000000;
	sram_mem[87498] = 16'b0000000000000000;
	sram_mem[87499] = 16'b0000000000000000;
	sram_mem[87500] = 16'b0000000000000000;
	sram_mem[87501] = 16'b0000000000000000;
	sram_mem[87502] = 16'b0000000000000000;
	sram_mem[87503] = 16'b0000000000000000;
	sram_mem[87504] = 16'b0000000000000000;
	sram_mem[87505] = 16'b0000000000000000;
	sram_mem[87506] = 16'b0000000000000000;
	sram_mem[87507] = 16'b0000000000000000;
	sram_mem[87508] = 16'b0000000000000000;
	sram_mem[87509] = 16'b0000000000000000;
	sram_mem[87510] = 16'b0000000000000000;
	sram_mem[87511] = 16'b0000000000000000;
	sram_mem[87512] = 16'b0000000000000000;
	sram_mem[87513] = 16'b0000000000000000;
	sram_mem[87514] = 16'b0000000000000000;
	sram_mem[87515] = 16'b0000000000000000;
	sram_mem[87516] = 16'b0000000000000000;
	sram_mem[87517] = 16'b0000000000000000;
	sram_mem[87518] = 16'b0000000000000000;
	sram_mem[87519] = 16'b0000000000000000;
	sram_mem[87520] = 16'b0000000000000000;
	sram_mem[87521] = 16'b0000000000000000;
	sram_mem[87522] = 16'b0000000000000000;
	sram_mem[87523] = 16'b0000000000000000;
	sram_mem[87524] = 16'b0000000000000000;
	sram_mem[87525] = 16'b0000000000000000;
	sram_mem[87526] = 16'b0000000000000000;
	sram_mem[87527] = 16'b0000000000000000;
	sram_mem[87528] = 16'b0000000000000000;
	sram_mem[87529] = 16'b0000000000000000;
	sram_mem[87530] = 16'b0000000000000000;
	sram_mem[87531] = 16'b0000000000000000;
	sram_mem[87532] = 16'b0000000000000000;
	sram_mem[87533] = 16'b0000000000000000;
	sram_mem[87534] = 16'b0000000000000000;
	sram_mem[87535] = 16'b0000000000000000;
	sram_mem[87536] = 16'b0000000000000000;
	sram_mem[87537] = 16'b0000000000000000;
	sram_mem[87538] = 16'b0000000000000000;
	sram_mem[87539] = 16'b0000000000000000;
	sram_mem[87540] = 16'b0000000000000000;
	sram_mem[87541] = 16'b0000000000000000;
	sram_mem[87542] = 16'b0000000000000000;
	sram_mem[87543] = 16'b0000000000000000;
	sram_mem[87544] = 16'b0000000000000000;
	sram_mem[87545] = 16'b0000000000000000;
	sram_mem[87546] = 16'b0000000000000000;
	sram_mem[87547] = 16'b0000000000000000;
	sram_mem[87548] = 16'b0000000000000000;
	sram_mem[87549] = 16'b0000000000000000;
	sram_mem[87550] = 16'b0000000000000000;
	sram_mem[87551] = 16'b0000000000000000;
	sram_mem[87552] = 16'b0000000000000000;
	sram_mem[87553] = 16'b0000000000000000;
	sram_mem[87554] = 16'b0000000000000000;
	sram_mem[87555] = 16'b0000000000000000;
	sram_mem[87556] = 16'b0000000000000000;
	sram_mem[87557] = 16'b0000000000000000;
	sram_mem[87558] = 16'b0000000000000000;
	sram_mem[87559] = 16'b0000000000000000;
	sram_mem[87560] = 16'b0000000000000000;
	sram_mem[87561] = 16'b0000000000000000;
	sram_mem[87562] = 16'b0000000000000000;
	sram_mem[87563] = 16'b0000000000000000;
	sram_mem[87564] = 16'b0000000000000000;
	sram_mem[87565] = 16'b0000000000000000;
	sram_mem[87566] = 16'b0000000000000000;
	sram_mem[87567] = 16'b0000000000000000;
	sram_mem[87568] = 16'b0000000000000000;
	sram_mem[87569] = 16'b0000000000000000;
	sram_mem[87570] = 16'b0000000000000000;
	sram_mem[87571] = 16'b0000000000000000;
	sram_mem[87572] = 16'b0000000000000000;
	sram_mem[87573] = 16'b0000000000000000;
	sram_mem[87574] = 16'b0000000000000000;
	sram_mem[87575] = 16'b0000000000000000;
	sram_mem[87576] = 16'b0000000000000000;
	sram_mem[87577] = 16'b0000000000000000;
	sram_mem[87578] = 16'b0000000000000000;
	sram_mem[87579] = 16'b0000000000000000;
	sram_mem[87580] = 16'b0000000000000000;
	sram_mem[87581] = 16'b0000000000000000;
	sram_mem[87582] = 16'b0000000000000000;
	sram_mem[87583] = 16'b0000000000000000;
	sram_mem[87584] = 16'b0000000000000000;
	sram_mem[87585] = 16'b0000000000000000;
	sram_mem[87586] = 16'b0000000000000000;
	sram_mem[87587] = 16'b0000000000000000;
	sram_mem[87588] = 16'b0000000000000000;
	sram_mem[87589] = 16'b0000000000000000;
	sram_mem[87590] = 16'b0000000000000000;
	sram_mem[87591] = 16'b0000000000000000;
	sram_mem[87592] = 16'b0000000000000000;
	sram_mem[87593] = 16'b0000000000000000;
	sram_mem[87594] = 16'b0000000000000000;
	sram_mem[87595] = 16'b0000000000000000;
	sram_mem[87596] = 16'b0000000000000000;
	sram_mem[87597] = 16'b0000000000000000;
	sram_mem[87598] = 16'b0000000000000000;
	sram_mem[87599] = 16'b0000000000000000;
	sram_mem[87600] = 16'b0000000000000000;
	sram_mem[87601] = 16'b0000000000000000;
	sram_mem[87602] = 16'b0000000000000000;
	sram_mem[87603] = 16'b0000000000000000;
	sram_mem[87604] = 16'b0000000000000000;
	sram_mem[87605] = 16'b0000000000000000;
	sram_mem[87606] = 16'b0000000000000000;
	sram_mem[87607] = 16'b0000000000000000;
	sram_mem[87608] = 16'b0000000000000000;
	sram_mem[87609] = 16'b0000000000000000;
	sram_mem[87610] = 16'b0000000000000000;
	sram_mem[87611] = 16'b0000000000000000;
	sram_mem[87612] = 16'b0000000000000000;
	sram_mem[87613] = 16'b0000000000000000;
	sram_mem[87614] = 16'b0000000000000000;
	sram_mem[87615] = 16'b0000000000000000;
	sram_mem[87616] = 16'b0000000000000000;
	sram_mem[87617] = 16'b0000000000000000;
	sram_mem[87618] = 16'b0000000000000000;
	sram_mem[87619] = 16'b0000000000000000;
	sram_mem[87620] = 16'b0000000000000000;
	sram_mem[87621] = 16'b0000000000000000;
	sram_mem[87622] = 16'b0000000000000000;
	sram_mem[87623] = 16'b0000000000000000;
	sram_mem[87624] = 16'b0000000000000000;
	sram_mem[87625] = 16'b0000000000000000;
	sram_mem[87626] = 16'b0000000000000000;
	sram_mem[87627] = 16'b0000000000000000;
	sram_mem[87628] = 16'b0000000000000000;
	sram_mem[87629] = 16'b0000000000000000;
	sram_mem[87630] = 16'b0000000000000000;
	sram_mem[87631] = 16'b0000000000000000;
	sram_mem[87632] = 16'b0000000000000000;
	sram_mem[87633] = 16'b0000000000000000;
	sram_mem[87634] = 16'b0000000000000000;
	sram_mem[87635] = 16'b0000000000000000;
	sram_mem[87636] = 16'b0000000000000000;
	sram_mem[87637] = 16'b0000000000000000;
	sram_mem[87638] = 16'b0000000000000000;
	sram_mem[87639] = 16'b0000000000000000;
	sram_mem[87640] = 16'b0000000000000000;
	sram_mem[87641] = 16'b0000000000000000;
	sram_mem[87642] = 16'b0000000000000000;
	sram_mem[87643] = 16'b0000000000000000;
	sram_mem[87644] = 16'b0000000000000000;
	sram_mem[87645] = 16'b0000000000000000;
	sram_mem[87646] = 16'b0000000000000000;
	sram_mem[87647] = 16'b0000000000000000;
	sram_mem[87648] = 16'b0000000000000000;
	sram_mem[87649] = 16'b0000000000000000;
	sram_mem[87650] = 16'b0000000000000000;
	sram_mem[87651] = 16'b0000000000000000;
	sram_mem[87652] = 16'b0000000000000000;
	sram_mem[87653] = 16'b0000000000000000;
	sram_mem[87654] = 16'b0000000000000000;
	sram_mem[87655] = 16'b0000000000000000;
	sram_mem[87656] = 16'b0000000000000000;
	sram_mem[87657] = 16'b0000000000000000;
	sram_mem[87658] = 16'b0000000000000000;
	sram_mem[87659] = 16'b0000000000000000;
	sram_mem[87660] = 16'b0000000000000000;
	sram_mem[87661] = 16'b0000000000000000;
	sram_mem[87662] = 16'b0000000000000000;
	sram_mem[87663] = 16'b0000000000000000;
	sram_mem[87664] = 16'b0000000000000000;
	sram_mem[87665] = 16'b0000000000000000;
	sram_mem[87666] = 16'b0000000000000000;
	sram_mem[87667] = 16'b0000000000000000;
	sram_mem[87668] = 16'b0000000000000000;
	sram_mem[87669] = 16'b0000000000000000;
	sram_mem[87670] = 16'b0000000000000000;
	sram_mem[87671] = 16'b0000000000000000;
	sram_mem[87672] = 16'b0000000000000000;
	sram_mem[87673] = 16'b0000000000000000;
	sram_mem[87674] = 16'b0000000000000000;
	sram_mem[87675] = 16'b0000000000000000;
	sram_mem[87676] = 16'b0000000000000000;
	sram_mem[87677] = 16'b0000000000000000;
	sram_mem[87678] = 16'b0000000000000000;
	sram_mem[87679] = 16'b0000000000000000;
	sram_mem[87680] = 16'b0000000000000000;
	sram_mem[87681] = 16'b0000000000000000;
	sram_mem[87682] = 16'b0000000000000000;
	sram_mem[87683] = 16'b0000000000000000;
	sram_mem[87684] = 16'b0000000000000000;
	sram_mem[87685] = 16'b0000000000000000;
	sram_mem[87686] = 16'b0000000000000000;
	sram_mem[87687] = 16'b0000000000000000;
	sram_mem[87688] = 16'b0000000000000000;
	sram_mem[87689] = 16'b0000000000000000;
	sram_mem[87690] = 16'b0000000000000000;
	sram_mem[87691] = 16'b0000000000000000;
	sram_mem[87692] = 16'b0000000000000000;
	sram_mem[87693] = 16'b0000000000000000;
	sram_mem[87694] = 16'b0000000000000000;
	sram_mem[87695] = 16'b0000000000000000;
	sram_mem[87696] = 16'b0000000000000000;
	sram_mem[87697] = 16'b0000000000000000;
	sram_mem[87698] = 16'b0000000000000000;
	sram_mem[87699] = 16'b0000000000000000;
	sram_mem[87700] = 16'b0000000000000000;
	sram_mem[87701] = 16'b0000000000000000;
	sram_mem[87702] = 16'b0000000000000000;
	sram_mem[87703] = 16'b0000000000000000;
	sram_mem[87704] = 16'b0000000000000000;
	sram_mem[87705] = 16'b0000000000000000;
	sram_mem[87706] = 16'b0000000000000000;
	sram_mem[87707] = 16'b0000000000000000;
	sram_mem[87708] = 16'b0000000000000000;
	sram_mem[87709] = 16'b0000000000000000;
	sram_mem[87710] = 16'b0000000000000000;
	sram_mem[87711] = 16'b0000000000000000;
	sram_mem[87712] = 16'b0000000000000000;
	sram_mem[87713] = 16'b0000000000000000;
	sram_mem[87714] = 16'b0000000000000000;
	sram_mem[87715] = 16'b0000000000000000;
	sram_mem[87716] = 16'b0000000000000000;
	sram_mem[87717] = 16'b0000000000000000;
	sram_mem[87718] = 16'b0000000000000000;
	sram_mem[87719] = 16'b0000000000000000;
	sram_mem[87720] = 16'b0000000000000000;
	sram_mem[87721] = 16'b0000000000000000;
	sram_mem[87722] = 16'b0000000000000000;
	sram_mem[87723] = 16'b0000000000000000;
	sram_mem[87724] = 16'b0000000000000000;
	sram_mem[87725] = 16'b0000000000000000;
	sram_mem[87726] = 16'b0000000000000000;
	sram_mem[87727] = 16'b0000000000000000;
	sram_mem[87728] = 16'b0000000000000000;
	sram_mem[87729] = 16'b0000000000000000;
	sram_mem[87730] = 16'b0000000000000000;
	sram_mem[87731] = 16'b0000000000000000;
	sram_mem[87732] = 16'b0000000000000000;
	sram_mem[87733] = 16'b0000000000000000;
	sram_mem[87734] = 16'b0000000000000000;
	sram_mem[87735] = 16'b0000000000000000;
	sram_mem[87736] = 16'b0000000000000000;
	sram_mem[87737] = 16'b0000000000000000;
	sram_mem[87738] = 16'b0000000000000000;
	sram_mem[87739] = 16'b0000000000000000;
	sram_mem[87740] = 16'b0000000000000000;
	sram_mem[87741] = 16'b0000000000000000;
	sram_mem[87742] = 16'b0000000000000000;
	sram_mem[87743] = 16'b0000000000000000;
	sram_mem[87744] = 16'b0000000000000000;
	sram_mem[87745] = 16'b0000000000000000;
	sram_mem[87746] = 16'b0000000000000000;
	sram_mem[87747] = 16'b0000000000000000;
	sram_mem[87748] = 16'b0000000000000000;
	sram_mem[87749] = 16'b0000000000000000;
	sram_mem[87750] = 16'b0000000000000000;
	sram_mem[87751] = 16'b0000000000000000;
	sram_mem[87752] = 16'b0000000000000000;
	sram_mem[87753] = 16'b0000000000000000;
	sram_mem[87754] = 16'b0000000000000000;
	sram_mem[87755] = 16'b0000000000000000;
	sram_mem[87756] = 16'b0000000000000000;
	sram_mem[87757] = 16'b0000000000000000;
	sram_mem[87758] = 16'b0000000000000000;
	sram_mem[87759] = 16'b0000000000000000;
	sram_mem[87760] = 16'b0000000000000000;
	sram_mem[87761] = 16'b0000000000000000;
	sram_mem[87762] = 16'b0000000000000000;
	sram_mem[87763] = 16'b0000000000000000;
	sram_mem[87764] = 16'b0000000000000000;
	sram_mem[87765] = 16'b0000000000000000;
	sram_mem[87766] = 16'b0000000000000000;
	sram_mem[87767] = 16'b0000000000000000;
	sram_mem[87768] = 16'b0000000000000000;
	sram_mem[87769] = 16'b0000000000000000;
	sram_mem[87770] = 16'b0000000000000000;
	sram_mem[87771] = 16'b0000000000000000;
	sram_mem[87772] = 16'b0000000000000000;
	sram_mem[87773] = 16'b0000000000000000;
	sram_mem[87774] = 16'b0000000000000000;
	sram_mem[87775] = 16'b0000000000000000;
	sram_mem[87776] = 16'b0000000000000000;
	sram_mem[87777] = 16'b0000000000000000;
	sram_mem[87778] = 16'b0000000000000000;
	sram_mem[87779] = 16'b0000000000000000;
	sram_mem[87780] = 16'b0000000000000000;
	sram_mem[87781] = 16'b0000000000000000;
	sram_mem[87782] = 16'b0000000000000000;
	sram_mem[87783] = 16'b0000000000000000;
	sram_mem[87784] = 16'b0000000000000000;
	sram_mem[87785] = 16'b0000000000000000;
	sram_mem[87786] = 16'b0000000000000000;
	sram_mem[87787] = 16'b0000000000000000;
	sram_mem[87788] = 16'b0000000000000000;
	sram_mem[87789] = 16'b0000000000000000;
	sram_mem[87790] = 16'b0000000000000000;
	sram_mem[87791] = 16'b0000000000000000;
	sram_mem[87792] = 16'b0000000000000000;
	sram_mem[87793] = 16'b0000000000000000;
	sram_mem[87794] = 16'b0000000000000000;
	sram_mem[87795] = 16'b0000000000000000;
	sram_mem[87796] = 16'b0000000000000000;
	sram_mem[87797] = 16'b0000000000000000;
	sram_mem[87798] = 16'b0000000000000000;
	sram_mem[87799] = 16'b0000000000000000;
	sram_mem[87800] = 16'b0000000000000000;
	sram_mem[87801] = 16'b0000000000000000;
	sram_mem[87802] = 16'b0000000000000000;
	sram_mem[87803] = 16'b0000000000000000;
	sram_mem[87804] = 16'b0000000000000000;
	sram_mem[87805] = 16'b0000000000000000;
	sram_mem[87806] = 16'b0000000000000000;
	sram_mem[87807] = 16'b0000000000000000;
	sram_mem[87808] = 16'b0000000000000000;
	sram_mem[87809] = 16'b0000000000000000;
	sram_mem[87810] = 16'b0000000000000000;
	sram_mem[87811] = 16'b0000000000000000;
	sram_mem[87812] = 16'b0000000000000000;
	sram_mem[87813] = 16'b0000000000000000;
	sram_mem[87814] = 16'b0000000000000000;
	sram_mem[87815] = 16'b0000000000000000;
	sram_mem[87816] = 16'b0000000000000000;
	sram_mem[87817] = 16'b0000000000000000;
	sram_mem[87818] = 16'b0000000000000000;
	sram_mem[87819] = 16'b0000000000000000;
	sram_mem[87820] = 16'b0000000000000000;
	sram_mem[87821] = 16'b0000000000000000;
	sram_mem[87822] = 16'b0000000000000000;
	sram_mem[87823] = 16'b0000000000000000;
	sram_mem[87824] = 16'b0000000000000000;
	sram_mem[87825] = 16'b0000000000000000;
	sram_mem[87826] = 16'b0000000000000000;
	sram_mem[87827] = 16'b0000000000000000;
	sram_mem[87828] = 16'b0000000000000000;
	sram_mem[87829] = 16'b0000000000000000;
	sram_mem[87830] = 16'b0000000000000000;
	sram_mem[87831] = 16'b0000000000000000;
	sram_mem[87832] = 16'b0000000000000000;
	sram_mem[87833] = 16'b0000000000000000;
	sram_mem[87834] = 16'b0000000000000000;
	sram_mem[87835] = 16'b0000000000000000;
	sram_mem[87836] = 16'b0000000000000000;
	sram_mem[87837] = 16'b0000000000000000;
	sram_mem[87838] = 16'b0000000000000000;
	sram_mem[87839] = 16'b0000000000000000;
	sram_mem[87840] = 16'b0000000000000000;
	sram_mem[87841] = 16'b0000000000000000;
	sram_mem[87842] = 16'b0000000000000000;
	sram_mem[87843] = 16'b0000000000000000;
	sram_mem[87844] = 16'b0000000000000000;
	sram_mem[87845] = 16'b0000000000000000;
	sram_mem[87846] = 16'b0000000000000000;
	sram_mem[87847] = 16'b0000000000000000;
	sram_mem[87848] = 16'b0000000000000000;
	sram_mem[87849] = 16'b0000000000000000;
	sram_mem[87850] = 16'b0000000000000000;
	sram_mem[87851] = 16'b0000000000000000;
	sram_mem[87852] = 16'b0000000000000000;
	sram_mem[87853] = 16'b0000000000000000;
	sram_mem[87854] = 16'b0000000000000000;
	sram_mem[87855] = 16'b0000000000000000;
	sram_mem[87856] = 16'b0000000000000000;
	sram_mem[87857] = 16'b0000000000000000;
	sram_mem[87858] = 16'b0000000000000000;
	sram_mem[87859] = 16'b0000000000000000;
	sram_mem[87860] = 16'b0000000000000000;
	sram_mem[87861] = 16'b0000000000000000;
	sram_mem[87862] = 16'b0000000000000000;
	sram_mem[87863] = 16'b0000000000000000;
	sram_mem[87864] = 16'b0000000000000000;
	sram_mem[87865] = 16'b0000000000000000;
	sram_mem[87866] = 16'b0000000000000000;
	sram_mem[87867] = 16'b0000000000000000;
	sram_mem[87868] = 16'b0000000000000000;
	sram_mem[87869] = 16'b0000000000000000;
	sram_mem[87870] = 16'b0000000000000000;
	sram_mem[87871] = 16'b0000000000000000;
	sram_mem[87872] = 16'b0000000000000000;
	sram_mem[87873] = 16'b0000000000000000;
	sram_mem[87874] = 16'b0000000000000000;
	sram_mem[87875] = 16'b0000000000000000;
	sram_mem[87876] = 16'b0000000000000000;
	sram_mem[87877] = 16'b0000000000000000;
	sram_mem[87878] = 16'b0000000000000000;
	sram_mem[87879] = 16'b0000000000000000;
	sram_mem[87880] = 16'b0000000000000000;
	sram_mem[87881] = 16'b0000000000000000;
	sram_mem[87882] = 16'b0000000000000000;
	sram_mem[87883] = 16'b0000000000000000;
	sram_mem[87884] = 16'b0000000000000000;
	sram_mem[87885] = 16'b0000000000000000;
	sram_mem[87886] = 16'b0000000000000000;
	sram_mem[87887] = 16'b0000000000000000;
	sram_mem[87888] = 16'b0000000000000000;
	sram_mem[87889] = 16'b0000000000000000;
	sram_mem[87890] = 16'b0000000000000000;
	sram_mem[87891] = 16'b0000000000000000;
	sram_mem[87892] = 16'b0000000000000000;
	sram_mem[87893] = 16'b0000000000000000;
	sram_mem[87894] = 16'b0000000000000000;
	sram_mem[87895] = 16'b0000000000000000;
	sram_mem[87896] = 16'b0000000000000000;
	sram_mem[87897] = 16'b0000000000000000;
	sram_mem[87898] = 16'b0000000000000000;
	sram_mem[87899] = 16'b0000000000000000;
	sram_mem[87900] = 16'b0000000000000000;
	sram_mem[87901] = 16'b0000000000000000;
	sram_mem[87902] = 16'b0000000000000000;
	sram_mem[87903] = 16'b0000000000000000;
	sram_mem[87904] = 16'b0000000000000000;
	sram_mem[87905] = 16'b0000000000000000;
	sram_mem[87906] = 16'b0000000000000000;
	sram_mem[87907] = 16'b0000000000000000;
	sram_mem[87908] = 16'b0000000000000000;
	sram_mem[87909] = 16'b0000000000000000;
	sram_mem[87910] = 16'b0000000000000000;
	sram_mem[87911] = 16'b0000000000000000;
	sram_mem[87912] = 16'b0000000000000000;
	sram_mem[87913] = 16'b0000000000000000;
	sram_mem[87914] = 16'b0000000000000000;
	sram_mem[87915] = 16'b0000000000000000;
	sram_mem[87916] = 16'b0000000000000000;
	sram_mem[87917] = 16'b0000000000000000;
	sram_mem[87918] = 16'b0000000000000000;
	sram_mem[87919] = 16'b0000000000000000;
	sram_mem[87920] = 16'b0000000000000000;
	sram_mem[87921] = 16'b0000000000000000;
	sram_mem[87922] = 16'b0000000000000000;
	sram_mem[87923] = 16'b0000000000000000;
	sram_mem[87924] = 16'b0000000000000000;
	sram_mem[87925] = 16'b0000000000000000;
	sram_mem[87926] = 16'b0000000000000000;
	sram_mem[87927] = 16'b0000000000000000;
	sram_mem[87928] = 16'b0000000000000000;
	sram_mem[87929] = 16'b0000000000000000;
	sram_mem[87930] = 16'b0000000000000000;
	sram_mem[87931] = 16'b0000000000000000;
	sram_mem[87932] = 16'b0000000000000000;
	sram_mem[87933] = 16'b0000000000000000;
	sram_mem[87934] = 16'b0000000000000000;
	sram_mem[87935] = 16'b0000000000000000;
	sram_mem[87936] = 16'b0000000000000000;
	sram_mem[87937] = 16'b0000000000000000;
	sram_mem[87938] = 16'b0000000000000000;
	sram_mem[87939] = 16'b0000000000000000;
	sram_mem[87940] = 16'b0000000000000000;
	sram_mem[87941] = 16'b0000000000000000;
	sram_mem[87942] = 16'b0000000000000000;
	sram_mem[87943] = 16'b0000000000000000;
	sram_mem[87944] = 16'b0000000000000000;
	sram_mem[87945] = 16'b0000000000000000;
	sram_mem[87946] = 16'b0000000000000000;
	sram_mem[87947] = 16'b0000000000000000;
	sram_mem[87948] = 16'b0000000000000000;
	sram_mem[87949] = 16'b0000000000000000;
	sram_mem[87950] = 16'b0000000000000000;
	sram_mem[87951] = 16'b0000000000000000;
	sram_mem[87952] = 16'b0000000000000000;
	sram_mem[87953] = 16'b0000000000000000;
	sram_mem[87954] = 16'b0000000000000000;
	sram_mem[87955] = 16'b0000000000000000;
	sram_mem[87956] = 16'b0000000000000000;
	sram_mem[87957] = 16'b0000000000000000;
	sram_mem[87958] = 16'b0000000000000000;
	sram_mem[87959] = 16'b0000000000000000;
	sram_mem[87960] = 16'b0000000000000000;
	sram_mem[87961] = 16'b0000000000000000;
	sram_mem[87962] = 16'b0000000000000000;
	sram_mem[87963] = 16'b0000000000000000;
	sram_mem[87964] = 16'b0000000000000000;
	sram_mem[87965] = 16'b0000000000000000;
	sram_mem[87966] = 16'b0000000000000000;
	sram_mem[87967] = 16'b0000000000000000;
	sram_mem[87968] = 16'b0000000000000000;
	sram_mem[87969] = 16'b0000000000000000;
	sram_mem[87970] = 16'b0000000000000000;
	sram_mem[87971] = 16'b0000000000000000;
	sram_mem[87972] = 16'b0000000000000000;
	sram_mem[87973] = 16'b0000000000000000;
	sram_mem[87974] = 16'b0000000000000000;
	sram_mem[87975] = 16'b0000000000000000;
	sram_mem[87976] = 16'b0000000000000000;
	sram_mem[87977] = 16'b0000000000000000;
	sram_mem[87978] = 16'b0000000000000000;
	sram_mem[87979] = 16'b0000000000000000;
	sram_mem[87980] = 16'b0000000000000000;
	sram_mem[87981] = 16'b0000000000000000;
	sram_mem[87982] = 16'b0000000000000000;
	sram_mem[87983] = 16'b0000000000000000;
	sram_mem[87984] = 16'b0000000000000000;
	sram_mem[87985] = 16'b0000000000000000;
	sram_mem[87986] = 16'b0000000000000000;
	sram_mem[87987] = 16'b0000000000000000;
	sram_mem[87988] = 16'b0000000000000000;
	sram_mem[87989] = 16'b0000000000000000;
	sram_mem[87990] = 16'b0000000000000000;
	sram_mem[87991] = 16'b0000000000000000;
	sram_mem[87992] = 16'b0000000000000000;
	sram_mem[87993] = 16'b0000000000000000;
	sram_mem[87994] = 16'b0000000000000000;
	sram_mem[87995] = 16'b0000000000000000;
	sram_mem[87996] = 16'b0000000000000000;
	sram_mem[87997] = 16'b0000000000000000;
	sram_mem[87998] = 16'b0000000000000000;
	sram_mem[87999] = 16'b0000000000000000;
	sram_mem[88000] = 16'b0000000000000000;
	sram_mem[88001] = 16'b0000000000000000;
	sram_mem[88002] = 16'b0000000000000000;
	sram_mem[88003] = 16'b0000000000000000;
	sram_mem[88004] = 16'b0000000000000000;
	sram_mem[88005] = 16'b0000000000000000;
	sram_mem[88006] = 16'b0000000000000000;
	sram_mem[88007] = 16'b0000000000000000;
	sram_mem[88008] = 16'b0000000000000000;
	sram_mem[88009] = 16'b0000000000000000;
	sram_mem[88010] = 16'b0000000000000000;
	sram_mem[88011] = 16'b0000000000000000;
	sram_mem[88012] = 16'b0000000000000000;
	sram_mem[88013] = 16'b0000000000000000;
	sram_mem[88014] = 16'b0000000000000000;
	sram_mem[88015] = 16'b0000000000000000;
	sram_mem[88016] = 16'b0000000000000000;
	sram_mem[88017] = 16'b0000000000000000;
	sram_mem[88018] = 16'b0000000000000000;
	sram_mem[88019] = 16'b0000000000000000;
	sram_mem[88020] = 16'b0000000000000000;
	sram_mem[88021] = 16'b0000000000000000;
	sram_mem[88022] = 16'b0000000000000000;
	sram_mem[88023] = 16'b0000000000000000;
	sram_mem[88024] = 16'b0000000000000000;
	sram_mem[88025] = 16'b0000000000000000;
	sram_mem[88026] = 16'b0000000000000000;
	sram_mem[88027] = 16'b0000000000000000;
	sram_mem[88028] = 16'b0000000000000000;
	sram_mem[88029] = 16'b0000000000000000;
	sram_mem[88030] = 16'b0000000000000000;
	sram_mem[88031] = 16'b0000000000000000;
	sram_mem[88032] = 16'b0000000000000000;
	sram_mem[88033] = 16'b0000000000000000;
	sram_mem[88034] = 16'b0000000000000000;
	sram_mem[88035] = 16'b0000000000000000;
	sram_mem[88036] = 16'b0000000000000000;
	sram_mem[88037] = 16'b0000000000000000;
	sram_mem[88038] = 16'b0000000000000000;
	sram_mem[88039] = 16'b0000000000000000;
	sram_mem[88040] = 16'b0000000000000000;
	sram_mem[88041] = 16'b0000000000000000;
	sram_mem[88042] = 16'b0000000000000000;
	sram_mem[88043] = 16'b0000000000000000;
	sram_mem[88044] = 16'b0000000000000000;
	sram_mem[88045] = 16'b0000000000000000;
	sram_mem[88046] = 16'b0000000000000000;
	sram_mem[88047] = 16'b0000000000000000;
	sram_mem[88048] = 16'b0000000000000000;
	sram_mem[88049] = 16'b0000000000000000;
	sram_mem[88050] = 16'b0000000000000000;
	sram_mem[88051] = 16'b0000000000000000;
	sram_mem[88052] = 16'b0000000000000000;
	sram_mem[88053] = 16'b0000000000000000;
	sram_mem[88054] = 16'b0000000000000000;
	sram_mem[88055] = 16'b0000000000000000;
	sram_mem[88056] = 16'b0000000000000000;
	sram_mem[88057] = 16'b0000000000000000;
	sram_mem[88058] = 16'b0000000000000000;
	sram_mem[88059] = 16'b0000000000000000;
	sram_mem[88060] = 16'b0000000000000000;
	sram_mem[88061] = 16'b0000000000000000;
	sram_mem[88062] = 16'b0000000000000000;
	sram_mem[88063] = 16'b0000000000000000;
	sram_mem[88064] = 16'b0000000000000000;
	sram_mem[88065] = 16'b0000000000000000;
	sram_mem[88066] = 16'b0000000000000000;
	sram_mem[88067] = 16'b0000000000000000;
	sram_mem[88068] = 16'b0000000000000000;
	sram_mem[88069] = 16'b0000000000000000;
	sram_mem[88070] = 16'b0000000000000000;
	sram_mem[88071] = 16'b0000000000000000;
	sram_mem[88072] = 16'b0000000000000000;
	sram_mem[88073] = 16'b0000000000000000;
	sram_mem[88074] = 16'b0000000000000000;
	sram_mem[88075] = 16'b0000000000000000;
	sram_mem[88076] = 16'b0000000000000000;
	sram_mem[88077] = 16'b0000000000000000;
	sram_mem[88078] = 16'b0000000000000000;
	sram_mem[88079] = 16'b0000000000000000;
	sram_mem[88080] = 16'b0000000000000000;
	sram_mem[88081] = 16'b0000000000000000;
	sram_mem[88082] = 16'b0000000000000000;
	sram_mem[88083] = 16'b0000000000000000;
	sram_mem[88084] = 16'b0000000000000000;
	sram_mem[88085] = 16'b0000000000000000;
	sram_mem[88086] = 16'b0000000000000000;
	sram_mem[88087] = 16'b0000000000000000;
	sram_mem[88088] = 16'b0000000000000000;
	sram_mem[88089] = 16'b0000000000000000;
	sram_mem[88090] = 16'b0000000000000000;
	sram_mem[88091] = 16'b0000000000000000;
	sram_mem[88092] = 16'b0000000000000000;
	sram_mem[88093] = 16'b0000000000000000;
	sram_mem[88094] = 16'b0000000000000000;
	sram_mem[88095] = 16'b0000000000000000;
	sram_mem[88096] = 16'b0000000000000000;
	sram_mem[88097] = 16'b0000000000000000;
	sram_mem[88098] = 16'b0000000000000000;
	sram_mem[88099] = 16'b0000000000000000;
	sram_mem[88100] = 16'b0000000000000000;
	sram_mem[88101] = 16'b0000000000000000;
	sram_mem[88102] = 16'b0000000000000000;
	sram_mem[88103] = 16'b0000000000000000;
	sram_mem[88104] = 16'b0000000000000000;
	sram_mem[88105] = 16'b0000000000000000;
	sram_mem[88106] = 16'b0000000000000000;
	sram_mem[88107] = 16'b0000000000000000;
	sram_mem[88108] = 16'b0000000000000000;
	sram_mem[88109] = 16'b0000000000000000;
	sram_mem[88110] = 16'b0000000000000000;
	sram_mem[88111] = 16'b0000000000000000;
	sram_mem[88112] = 16'b0000000000000000;
	sram_mem[88113] = 16'b0000000000000000;
	sram_mem[88114] = 16'b0000000000000000;
	sram_mem[88115] = 16'b0000000000000000;
	sram_mem[88116] = 16'b0000000000000000;
	sram_mem[88117] = 16'b0000000000000000;
	sram_mem[88118] = 16'b0000000000000000;
	sram_mem[88119] = 16'b0000000000000000;
	sram_mem[88120] = 16'b0000000000000000;
	sram_mem[88121] = 16'b0000000000000000;
	sram_mem[88122] = 16'b0000000000000000;
	sram_mem[88123] = 16'b0000000000000000;
	sram_mem[88124] = 16'b0000000000000000;
	sram_mem[88125] = 16'b0000000000000000;
	sram_mem[88126] = 16'b0000000000000000;
	sram_mem[88127] = 16'b0000000000000000;
	sram_mem[88128] = 16'b0000000000000000;
	sram_mem[88129] = 16'b0000000000000000;
	sram_mem[88130] = 16'b0000000000000000;
	sram_mem[88131] = 16'b0000000000000000;
	sram_mem[88132] = 16'b0000000000000000;
	sram_mem[88133] = 16'b0000000000000000;
	sram_mem[88134] = 16'b0000000000000000;
	sram_mem[88135] = 16'b0000000000000000;
	sram_mem[88136] = 16'b0000000000000000;
	sram_mem[88137] = 16'b0000000000000000;
	sram_mem[88138] = 16'b0000000000000000;
	sram_mem[88139] = 16'b0000000000000000;
	sram_mem[88140] = 16'b0000000000000000;
	sram_mem[88141] = 16'b0000000000000000;
	sram_mem[88142] = 16'b0000000000000000;
	sram_mem[88143] = 16'b0000000000000000;
	sram_mem[88144] = 16'b0000000000000000;
	sram_mem[88145] = 16'b0000000000000000;
	sram_mem[88146] = 16'b0000000000000000;
	sram_mem[88147] = 16'b0000000000000000;
	sram_mem[88148] = 16'b0000000000000000;
	sram_mem[88149] = 16'b0000000000000000;
	sram_mem[88150] = 16'b0000000000000000;
	sram_mem[88151] = 16'b0000000000000000;
	sram_mem[88152] = 16'b0000000000000000;
	sram_mem[88153] = 16'b0000000000000000;
	sram_mem[88154] = 16'b0000000000000000;
	sram_mem[88155] = 16'b0000000000000000;
	sram_mem[88156] = 16'b0000000000000000;
	sram_mem[88157] = 16'b0000000000000000;
	sram_mem[88158] = 16'b0000000000000000;
	sram_mem[88159] = 16'b0000000000000000;
	sram_mem[88160] = 16'b0000000000000000;
	sram_mem[88161] = 16'b0000000000000000;
	sram_mem[88162] = 16'b0000000000000000;
	sram_mem[88163] = 16'b0000000000000000;
	sram_mem[88164] = 16'b0000000000000000;
	sram_mem[88165] = 16'b0000000000000000;
	sram_mem[88166] = 16'b0000000000000000;
	sram_mem[88167] = 16'b0000000000000000;
	sram_mem[88168] = 16'b0000000000000000;
	sram_mem[88169] = 16'b0000000000000000;
	sram_mem[88170] = 16'b0000000000000000;
	sram_mem[88171] = 16'b0000000000000000;
	sram_mem[88172] = 16'b0000000000000000;
	sram_mem[88173] = 16'b0000000000000000;
	sram_mem[88174] = 16'b0000000000000000;
	sram_mem[88175] = 16'b0000000000000000;
	sram_mem[88176] = 16'b0000000000000000;
	sram_mem[88177] = 16'b0000000000000000;
	sram_mem[88178] = 16'b0000000000000000;
	sram_mem[88179] = 16'b0000000000000000;
	sram_mem[88180] = 16'b0000000000000000;
	sram_mem[88181] = 16'b0000000000000000;
	sram_mem[88182] = 16'b0000000000000000;
	sram_mem[88183] = 16'b0000000000000000;
	sram_mem[88184] = 16'b0000000000000000;
	sram_mem[88185] = 16'b0000000000000000;
	sram_mem[88186] = 16'b0000000000000000;
	sram_mem[88187] = 16'b0000000000000000;
	sram_mem[88188] = 16'b0000000000000000;
	sram_mem[88189] = 16'b0000000000000000;
	sram_mem[88190] = 16'b0000000000000000;
	sram_mem[88191] = 16'b0000000000000000;
	sram_mem[88192] = 16'b0000000000000000;
	sram_mem[88193] = 16'b0000000000000000;
	sram_mem[88194] = 16'b0000000000000000;
	sram_mem[88195] = 16'b0000000000000000;
	sram_mem[88196] = 16'b0000000000000000;
	sram_mem[88197] = 16'b0000000000000000;
	sram_mem[88198] = 16'b0000000000000000;
	sram_mem[88199] = 16'b0000000000000000;
	sram_mem[88200] = 16'b0000000000000000;
	sram_mem[88201] = 16'b0000000000000000;
	sram_mem[88202] = 16'b0000000000000000;
	sram_mem[88203] = 16'b0000000000000000;
	sram_mem[88204] = 16'b0000000000000000;
	sram_mem[88205] = 16'b0000000000000000;
	sram_mem[88206] = 16'b0000000000000000;
	sram_mem[88207] = 16'b0000000000000000;
	sram_mem[88208] = 16'b0000000000000000;
	sram_mem[88209] = 16'b0000000000000000;
	sram_mem[88210] = 16'b0000000000000000;
	sram_mem[88211] = 16'b0000000000000000;
	sram_mem[88212] = 16'b0000000000000000;
	sram_mem[88213] = 16'b0000000000000000;
	sram_mem[88214] = 16'b0000000000000000;
	sram_mem[88215] = 16'b0000000000000000;
	sram_mem[88216] = 16'b0000000000000000;
	sram_mem[88217] = 16'b0000000000000000;
	sram_mem[88218] = 16'b0000000000000000;
	sram_mem[88219] = 16'b0000000000000000;
	sram_mem[88220] = 16'b0000000000000000;
	sram_mem[88221] = 16'b0000000000000000;
	sram_mem[88222] = 16'b0000000000000000;
	sram_mem[88223] = 16'b0000000000000000;
	sram_mem[88224] = 16'b0000000000000000;
	sram_mem[88225] = 16'b0000000000000000;
	sram_mem[88226] = 16'b0000000000000000;
	sram_mem[88227] = 16'b0000000000000000;
	sram_mem[88228] = 16'b0000000000000000;
	sram_mem[88229] = 16'b0000000000000000;
	sram_mem[88230] = 16'b0000000000000000;
	sram_mem[88231] = 16'b0000000000000000;
	sram_mem[88232] = 16'b0000000000000000;
	sram_mem[88233] = 16'b0000000000000000;
	sram_mem[88234] = 16'b0000000000000000;
	sram_mem[88235] = 16'b0000000000000000;
	sram_mem[88236] = 16'b0000000000000000;
	sram_mem[88237] = 16'b0000000000000000;
	sram_mem[88238] = 16'b0000000000000000;
	sram_mem[88239] = 16'b0000000000000000;
	sram_mem[88240] = 16'b0000000000000000;
	sram_mem[88241] = 16'b0000000000000000;
	sram_mem[88242] = 16'b0000000000000000;
	sram_mem[88243] = 16'b0000000000000000;
	sram_mem[88244] = 16'b0000000000000000;
	sram_mem[88245] = 16'b0000000000000000;
	sram_mem[88246] = 16'b0000000000000000;
	sram_mem[88247] = 16'b0000000000000000;
	sram_mem[88248] = 16'b0000000000000000;
	sram_mem[88249] = 16'b0000000000000000;
	sram_mem[88250] = 16'b0000000000000000;
	sram_mem[88251] = 16'b0000000000000000;
	sram_mem[88252] = 16'b0000000000000000;
	sram_mem[88253] = 16'b0000000000000000;
	sram_mem[88254] = 16'b0000000000000000;
	sram_mem[88255] = 16'b0000000000000000;
	sram_mem[88256] = 16'b0000000000000000;
	sram_mem[88257] = 16'b0000000000000000;
	sram_mem[88258] = 16'b0000000000000000;
	sram_mem[88259] = 16'b0000000000000000;
	sram_mem[88260] = 16'b0000000000000000;
	sram_mem[88261] = 16'b0000000000000000;
	sram_mem[88262] = 16'b0000000000000000;
	sram_mem[88263] = 16'b0000000000000000;
	sram_mem[88264] = 16'b0000000000000000;
	sram_mem[88265] = 16'b0000000000000000;
	sram_mem[88266] = 16'b0000000000000000;
	sram_mem[88267] = 16'b0000000000000000;
	sram_mem[88268] = 16'b0000000000000000;
	sram_mem[88269] = 16'b0000000000000000;
	sram_mem[88270] = 16'b0000000000000000;
	sram_mem[88271] = 16'b0000000000000000;
	sram_mem[88272] = 16'b0000000000000000;
	sram_mem[88273] = 16'b0000000000000000;
	sram_mem[88274] = 16'b0000000000000000;
	sram_mem[88275] = 16'b0000000000000000;
	sram_mem[88276] = 16'b0000000000000000;
	sram_mem[88277] = 16'b0000000000000000;
	sram_mem[88278] = 16'b0000000000000000;
	sram_mem[88279] = 16'b0000000000000000;
	sram_mem[88280] = 16'b0000000000000000;
	sram_mem[88281] = 16'b0000000000000000;
	sram_mem[88282] = 16'b0000000000000000;
	sram_mem[88283] = 16'b0000000000000000;
	sram_mem[88284] = 16'b0000000000000000;
	sram_mem[88285] = 16'b0000000000000000;
	sram_mem[88286] = 16'b0000000000000000;
	sram_mem[88287] = 16'b0000000000000000;
	sram_mem[88288] = 16'b0000000000000000;
	sram_mem[88289] = 16'b0000000000000000;
	sram_mem[88290] = 16'b0000000000000000;
	sram_mem[88291] = 16'b0000000000000000;
	sram_mem[88292] = 16'b0000000000000000;
	sram_mem[88293] = 16'b0000000000000000;
	sram_mem[88294] = 16'b0000000000000000;
	sram_mem[88295] = 16'b0000000000000000;
	sram_mem[88296] = 16'b0000000000000000;
	sram_mem[88297] = 16'b0000000000000000;
	sram_mem[88298] = 16'b0000000000000000;
	sram_mem[88299] = 16'b0000000000000000;
	sram_mem[88300] = 16'b0000000000000000;
	sram_mem[88301] = 16'b0000000000000000;
	sram_mem[88302] = 16'b0000000000000000;
	sram_mem[88303] = 16'b0000000000000000;
	sram_mem[88304] = 16'b0000000000000000;
	sram_mem[88305] = 16'b0000000000000000;
	sram_mem[88306] = 16'b0000000000000000;
	sram_mem[88307] = 16'b0000000000000000;
	sram_mem[88308] = 16'b0000000000000000;
	sram_mem[88309] = 16'b0000000000000000;
	sram_mem[88310] = 16'b0000000000000000;
	sram_mem[88311] = 16'b0000000000000000;
	sram_mem[88312] = 16'b0000000000000000;
	sram_mem[88313] = 16'b0000000000000000;
	sram_mem[88314] = 16'b0000000000000000;
	sram_mem[88315] = 16'b0000000000000000;
	sram_mem[88316] = 16'b0000000000000000;
	sram_mem[88317] = 16'b0000000000000000;
	sram_mem[88318] = 16'b0000000000000000;
	sram_mem[88319] = 16'b0000000000000000;
	sram_mem[88320] = 16'b0000000000000000;
	sram_mem[88321] = 16'b0000000000000000;
	sram_mem[88322] = 16'b0000000000000000;
	sram_mem[88323] = 16'b0000000000000000;
	sram_mem[88324] = 16'b0000000000000000;
	sram_mem[88325] = 16'b0000000000000000;
	sram_mem[88326] = 16'b0000000000000000;
	sram_mem[88327] = 16'b0000000000000000;
	sram_mem[88328] = 16'b0000000000000000;
	sram_mem[88329] = 16'b0000000000000000;
	sram_mem[88330] = 16'b0000000000000000;
	sram_mem[88331] = 16'b0000000000000000;
	sram_mem[88332] = 16'b0000000000000000;
	sram_mem[88333] = 16'b0000000000000000;
	sram_mem[88334] = 16'b0000000000000000;
	sram_mem[88335] = 16'b0000000000000000;
	sram_mem[88336] = 16'b0000000000000000;
	sram_mem[88337] = 16'b0000000000000000;
	sram_mem[88338] = 16'b0000000000000000;
	sram_mem[88339] = 16'b0000000000000000;
	sram_mem[88340] = 16'b0000000000000000;
	sram_mem[88341] = 16'b0000000000000000;
	sram_mem[88342] = 16'b0000000000000000;
	sram_mem[88343] = 16'b0000000000000000;
	sram_mem[88344] = 16'b0000000000000000;
	sram_mem[88345] = 16'b0000000000000000;
	sram_mem[88346] = 16'b0000000000000000;
	sram_mem[88347] = 16'b0000000000000000;
	sram_mem[88348] = 16'b0000000000000000;
	sram_mem[88349] = 16'b0000000000000000;
	sram_mem[88350] = 16'b0000000000000000;
	sram_mem[88351] = 16'b0000000000000000;
	sram_mem[88352] = 16'b0000000000000000;
	sram_mem[88353] = 16'b0000000000000000;
	sram_mem[88354] = 16'b0000000000000000;
	sram_mem[88355] = 16'b0000000000000000;
	sram_mem[88356] = 16'b0000000000000000;
	sram_mem[88357] = 16'b0000000000000000;
	sram_mem[88358] = 16'b0000000000000000;
	sram_mem[88359] = 16'b0000000000000000;
	sram_mem[88360] = 16'b0000000000000000;
	sram_mem[88361] = 16'b0000000000000000;
	sram_mem[88362] = 16'b0000000000000000;
	sram_mem[88363] = 16'b0000000000000000;
	sram_mem[88364] = 16'b0000000000000000;
	sram_mem[88365] = 16'b0000000000000000;
	sram_mem[88366] = 16'b0000000000000000;
	sram_mem[88367] = 16'b0000000000000000;
	sram_mem[88368] = 16'b0000000000000000;
	sram_mem[88369] = 16'b0000000000000000;
	sram_mem[88370] = 16'b0000000000000000;
	sram_mem[88371] = 16'b0000000000000000;
	sram_mem[88372] = 16'b0000000000000000;
	sram_mem[88373] = 16'b0000000000000000;
	sram_mem[88374] = 16'b0000000000000000;
	sram_mem[88375] = 16'b0000000000000000;
	sram_mem[88376] = 16'b0000000000000000;
	sram_mem[88377] = 16'b0000000000000000;
	sram_mem[88378] = 16'b0000000000000000;
	sram_mem[88379] = 16'b0000000000000000;
	sram_mem[88380] = 16'b0000000000000000;
	sram_mem[88381] = 16'b0000000000000000;
	sram_mem[88382] = 16'b0000000000000000;
	sram_mem[88383] = 16'b0000000000000000;
	sram_mem[88384] = 16'b0000000000000000;
	sram_mem[88385] = 16'b0000000000000000;
	sram_mem[88386] = 16'b0000000000000000;
	sram_mem[88387] = 16'b0000000000000000;
	sram_mem[88388] = 16'b0000000000000000;
	sram_mem[88389] = 16'b0000000000000000;
	sram_mem[88390] = 16'b0000000000000000;
	sram_mem[88391] = 16'b0000000000000000;
	sram_mem[88392] = 16'b0000000000000000;
	sram_mem[88393] = 16'b0000000000000000;
	sram_mem[88394] = 16'b0000000000000000;
	sram_mem[88395] = 16'b0000000000000000;
	sram_mem[88396] = 16'b0000000000000000;
	sram_mem[88397] = 16'b0000000000000000;
	sram_mem[88398] = 16'b0000000000000000;
	sram_mem[88399] = 16'b0000000000000000;
	sram_mem[88400] = 16'b0000000000000000;
	sram_mem[88401] = 16'b0000000000000000;
	sram_mem[88402] = 16'b0000000000000000;
	sram_mem[88403] = 16'b0000000000000000;
	sram_mem[88404] = 16'b0000000000000000;
	sram_mem[88405] = 16'b0000000000000000;
	sram_mem[88406] = 16'b0000000000000000;
	sram_mem[88407] = 16'b0000000000000000;
	sram_mem[88408] = 16'b0000000000000000;
	sram_mem[88409] = 16'b0000000000000000;
	sram_mem[88410] = 16'b0000000000000000;
	sram_mem[88411] = 16'b0000000000000000;
	sram_mem[88412] = 16'b0000000000000000;
	sram_mem[88413] = 16'b0000000000000000;
	sram_mem[88414] = 16'b0000000000000000;
	sram_mem[88415] = 16'b0000000000000000;
	sram_mem[88416] = 16'b0000000000000000;
	sram_mem[88417] = 16'b0000000000000000;
	sram_mem[88418] = 16'b0000000000000000;
	sram_mem[88419] = 16'b0000000000000000;
	sram_mem[88420] = 16'b0000000000000000;
	sram_mem[88421] = 16'b0000000000000000;
	sram_mem[88422] = 16'b0000000000000000;
	sram_mem[88423] = 16'b0000000000000000;
	sram_mem[88424] = 16'b0000000000000000;
	sram_mem[88425] = 16'b0000000000000000;
	sram_mem[88426] = 16'b0000000000000000;
	sram_mem[88427] = 16'b0000000000000000;
	sram_mem[88428] = 16'b0000000000000000;
	sram_mem[88429] = 16'b0000000000000000;
	sram_mem[88430] = 16'b0000000000000000;
	sram_mem[88431] = 16'b0000000000000000;
	sram_mem[88432] = 16'b0000000000000000;
	sram_mem[88433] = 16'b0000000000000000;
	sram_mem[88434] = 16'b0000000000000000;
	sram_mem[88435] = 16'b0000000000000000;
	sram_mem[88436] = 16'b0000000000000000;
	sram_mem[88437] = 16'b0000000000000000;
	sram_mem[88438] = 16'b0000000000000000;
	sram_mem[88439] = 16'b0000000000000000;
	sram_mem[88440] = 16'b0000000000000000;
	sram_mem[88441] = 16'b0000000000000000;
	sram_mem[88442] = 16'b0000000000000000;
	sram_mem[88443] = 16'b0000000000000000;
	sram_mem[88444] = 16'b0000000000000000;
	sram_mem[88445] = 16'b0000000000000000;
	sram_mem[88446] = 16'b0000000000000000;
	sram_mem[88447] = 16'b0000000000000000;
	sram_mem[88448] = 16'b0000000000000000;
	sram_mem[88449] = 16'b0000000000000000;
	sram_mem[88450] = 16'b0000000000000000;
	sram_mem[88451] = 16'b0000000000000000;
	sram_mem[88452] = 16'b0000000000000000;
	sram_mem[88453] = 16'b0000000000000000;
	sram_mem[88454] = 16'b0000000000000000;
	sram_mem[88455] = 16'b0000000000000000;
	sram_mem[88456] = 16'b0000000000000000;
	sram_mem[88457] = 16'b0000000000000000;
	sram_mem[88458] = 16'b0000000000000000;
	sram_mem[88459] = 16'b0000000000000000;
	sram_mem[88460] = 16'b0000000000000000;
	sram_mem[88461] = 16'b0000000000000000;
	sram_mem[88462] = 16'b0000000000000000;
	sram_mem[88463] = 16'b0000000000000000;
	sram_mem[88464] = 16'b0000000000000000;
	sram_mem[88465] = 16'b0000000000000000;
	sram_mem[88466] = 16'b0000000000000000;
	sram_mem[88467] = 16'b0000000000000000;
	sram_mem[88468] = 16'b0000000000000000;
	sram_mem[88469] = 16'b0000000000000000;
	sram_mem[88470] = 16'b0000000000000000;
	sram_mem[88471] = 16'b0000000000000000;
	sram_mem[88472] = 16'b0000000000000000;
	sram_mem[88473] = 16'b0000000000000000;
	sram_mem[88474] = 16'b0000000000000000;
	sram_mem[88475] = 16'b0000000000000000;
	sram_mem[88476] = 16'b0000000000000000;
	sram_mem[88477] = 16'b0000000000000000;
	sram_mem[88478] = 16'b0000000000000000;
	sram_mem[88479] = 16'b0000000000000000;
	sram_mem[88480] = 16'b0000000000000000;
	sram_mem[88481] = 16'b0000000000000000;
	sram_mem[88482] = 16'b0000000000000000;
	sram_mem[88483] = 16'b0000000000000000;
	sram_mem[88484] = 16'b0000000000000000;
	sram_mem[88485] = 16'b0000000000000000;
	sram_mem[88486] = 16'b0000000000000000;
	sram_mem[88487] = 16'b0000000000000000;
	sram_mem[88488] = 16'b0000000000000000;
	sram_mem[88489] = 16'b0000000000000000;
	sram_mem[88490] = 16'b0000000000000000;
	sram_mem[88491] = 16'b0000000000000000;
	sram_mem[88492] = 16'b0000000000000000;
	sram_mem[88493] = 16'b0000000000000000;
	sram_mem[88494] = 16'b0000000000000000;
	sram_mem[88495] = 16'b0000000000000000;
	sram_mem[88496] = 16'b0000000000000000;
	sram_mem[88497] = 16'b0000000000000000;
	sram_mem[88498] = 16'b0000000000000000;
	sram_mem[88499] = 16'b0000000000000000;
	sram_mem[88500] = 16'b0000000000000000;
	sram_mem[88501] = 16'b0000000000000000;
	sram_mem[88502] = 16'b0000000000000000;
	sram_mem[88503] = 16'b0000000000000000;
	sram_mem[88504] = 16'b0000000000000000;
	sram_mem[88505] = 16'b0000000000000000;
	sram_mem[88506] = 16'b0000000000000000;
	sram_mem[88507] = 16'b0000000000000000;
	sram_mem[88508] = 16'b0000000000000000;
	sram_mem[88509] = 16'b0000000000000000;
	sram_mem[88510] = 16'b0000000000000000;
	sram_mem[88511] = 16'b0000000000000000;
	sram_mem[88512] = 16'b0000000000000000;
	sram_mem[88513] = 16'b0000000000000000;
	sram_mem[88514] = 16'b0000000000000000;
	sram_mem[88515] = 16'b0000000000000000;
	sram_mem[88516] = 16'b0000000000000000;
	sram_mem[88517] = 16'b0000000000000000;
	sram_mem[88518] = 16'b0000000000000000;
	sram_mem[88519] = 16'b0000000000000000;
	sram_mem[88520] = 16'b0000000000000000;
	sram_mem[88521] = 16'b0000000000000000;
	sram_mem[88522] = 16'b0000000000000000;
	sram_mem[88523] = 16'b0000000000000000;
	sram_mem[88524] = 16'b0000000000000000;
	sram_mem[88525] = 16'b0000000000000000;
	sram_mem[88526] = 16'b0000000000000000;
	sram_mem[88527] = 16'b0000000000000000;
	sram_mem[88528] = 16'b0000000000000000;
	sram_mem[88529] = 16'b0000000000000000;
	sram_mem[88530] = 16'b0000000000000000;
	sram_mem[88531] = 16'b0000000000000000;
	sram_mem[88532] = 16'b0000000000000000;
	sram_mem[88533] = 16'b0000000000000000;
	sram_mem[88534] = 16'b0000000000000000;
	sram_mem[88535] = 16'b0000000000000000;
	sram_mem[88536] = 16'b0000000000000000;
	sram_mem[88537] = 16'b0000000000000000;
	sram_mem[88538] = 16'b0000000000000000;
	sram_mem[88539] = 16'b0000000000000000;
	sram_mem[88540] = 16'b0000000000000000;
	sram_mem[88541] = 16'b0000000000000000;
	sram_mem[88542] = 16'b0000000000000000;
	sram_mem[88543] = 16'b0000000000000000;
	sram_mem[88544] = 16'b0000000000000000;
	sram_mem[88545] = 16'b0000000000000000;
	sram_mem[88546] = 16'b0000000000000000;
	sram_mem[88547] = 16'b0000000000000000;
	sram_mem[88548] = 16'b0000000000000000;
	sram_mem[88549] = 16'b0000000000000000;
	sram_mem[88550] = 16'b0000000000000000;
	sram_mem[88551] = 16'b0000000000000000;
	sram_mem[88552] = 16'b0000000000000000;
	sram_mem[88553] = 16'b0000000000000000;
	sram_mem[88554] = 16'b0000000000000000;
	sram_mem[88555] = 16'b0000000000000000;
	sram_mem[88556] = 16'b0000000000000000;
	sram_mem[88557] = 16'b0000000000000000;
	sram_mem[88558] = 16'b0000000000000000;
	sram_mem[88559] = 16'b0000000000000000;
	sram_mem[88560] = 16'b0000000000000000;
	sram_mem[88561] = 16'b0000000000000000;
	sram_mem[88562] = 16'b0000000000000000;
	sram_mem[88563] = 16'b0000000000000000;
	sram_mem[88564] = 16'b0000000000000000;
	sram_mem[88565] = 16'b0000000000000000;
	sram_mem[88566] = 16'b0000000000000000;
	sram_mem[88567] = 16'b0000000000000000;
	sram_mem[88568] = 16'b0000000000000000;
	sram_mem[88569] = 16'b0000000000000000;
	sram_mem[88570] = 16'b0000000000000000;
	sram_mem[88571] = 16'b0000000000000000;
	sram_mem[88572] = 16'b0000000000000000;
	sram_mem[88573] = 16'b0000000000000000;
	sram_mem[88574] = 16'b0000000000000000;
	sram_mem[88575] = 16'b0000000000000000;
	sram_mem[88576] = 16'b0000000000000000;
	sram_mem[88577] = 16'b0000000000000000;
	sram_mem[88578] = 16'b0000000000000000;
	sram_mem[88579] = 16'b0000000000000000;
	sram_mem[88580] = 16'b0000000000000000;
	sram_mem[88581] = 16'b0000000000000000;
	sram_mem[88582] = 16'b0000000000000000;
	sram_mem[88583] = 16'b0000000000000000;
	sram_mem[88584] = 16'b0000000000000000;
	sram_mem[88585] = 16'b0000000000000000;
	sram_mem[88586] = 16'b0000000000000000;
	sram_mem[88587] = 16'b0000000000000000;
	sram_mem[88588] = 16'b0000000000000000;
	sram_mem[88589] = 16'b0000000000000000;
	sram_mem[88590] = 16'b0000000000000000;
	sram_mem[88591] = 16'b0000000000000000;
	sram_mem[88592] = 16'b0000000000000000;
	sram_mem[88593] = 16'b0000000000000000;
	sram_mem[88594] = 16'b0000000000000000;
	sram_mem[88595] = 16'b0000000000000000;
	sram_mem[88596] = 16'b0000000000000000;
	sram_mem[88597] = 16'b0000000000000000;
	sram_mem[88598] = 16'b0000000000000000;
	sram_mem[88599] = 16'b0000000000000000;
	sram_mem[88600] = 16'b0000000000000000;
	sram_mem[88601] = 16'b0000000000000000;
	sram_mem[88602] = 16'b0000000000000000;
	sram_mem[88603] = 16'b0000000000000000;
	sram_mem[88604] = 16'b0000000000000000;
	sram_mem[88605] = 16'b0000000000000000;
	sram_mem[88606] = 16'b0000000000000000;
	sram_mem[88607] = 16'b0000000000000000;
	sram_mem[88608] = 16'b0000000000000000;
	sram_mem[88609] = 16'b0000000000000000;
	sram_mem[88610] = 16'b0000000000000000;
	sram_mem[88611] = 16'b0000000000000000;
	sram_mem[88612] = 16'b0000000000000000;
	sram_mem[88613] = 16'b0000000000000000;
	sram_mem[88614] = 16'b0000000000000000;
	sram_mem[88615] = 16'b0000000000000000;
	sram_mem[88616] = 16'b0000000000000000;
	sram_mem[88617] = 16'b0000000000000000;
	sram_mem[88618] = 16'b0000000000000000;
	sram_mem[88619] = 16'b0000000000000000;
	sram_mem[88620] = 16'b0000000000000000;
	sram_mem[88621] = 16'b0000000000000000;
	sram_mem[88622] = 16'b0000000000000000;
	sram_mem[88623] = 16'b0000000000000000;
	sram_mem[88624] = 16'b0000000000000000;
	sram_mem[88625] = 16'b0000000000000000;
	sram_mem[88626] = 16'b0000000000000000;
	sram_mem[88627] = 16'b0000000000000000;
	sram_mem[88628] = 16'b0000000000000000;
	sram_mem[88629] = 16'b0000000000000000;
	sram_mem[88630] = 16'b0000000000000000;
	sram_mem[88631] = 16'b0000000000000000;
	sram_mem[88632] = 16'b0000000000000000;
	sram_mem[88633] = 16'b0000000000000000;
	sram_mem[88634] = 16'b0000000000000000;
	sram_mem[88635] = 16'b0000000000000000;
	sram_mem[88636] = 16'b0000000000000000;
	sram_mem[88637] = 16'b0000000000000000;
	sram_mem[88638] = 16'b0000000000000000;
	sram_mem[88639] = 16'b0000000000000000;
	sram_mem[88640] = 16'b0000000000000000;
	sram_mem[88641] = 16'b0000000000000000;
	sram_mem[88642] = 16'b0000000000000000;
	sram_mem[88643] = 16'b0000000000000000;
	sram_mem[88644] = 16'b0000000000000000;
	sram_mem[88645] = 16'b0000000000000000;
	sram_mem[88646] = 16'b0000000000000000;
	sram_mem[88647] = 16'b0000000000000000;
	sram_mem[88648] = 16'b0000000000000000;
	sram_mem[88649] = 16'b0000000000000000;
	sram_mem[88650] = 16'b0000000000000000;
	sram_mem[88651] = 16'b0000000000000000;
	sram_mem[88652] = 16'b0000000000000000;
	sram_mem[88653] = 16'b0000000000000000;
	sram_mem[88654] = 16'b0000000000000000;
	sram_mem[88655] = 16'b0000000000000000;
	sram_mem[88656] = 16'b0000000000000000;
	sram_mem[88657] = 16'b0000000000000000;
	sram_mem[88658] = 16'b0000000000000000;
	sram_mem[88659] = 16'b0000000000000000;
	sram_mem[88660] = 16'b0000000000000000;
	sram_mem[88661] = 16'b0000000000000000;
	sram_mem[88662] = 16'b0000000000000000;
	sram_mem[88663] = 16'b0000000000000000;
	sram_mem[88664] = 16'b0000000000000000;
	sram_mem[88665] = 16'b0000000000000000;
	sram_mem[88666] = 16'b0000000000000000;
	sram_mem[88667] = 16'b0000000000000000;
	sram_mem[88668] = 16'b0000000000000000;
	sram_mem[88669] = 16'b0000000000000000;
	sram_mem[88670] = 16'b0000000000000000;
	sram_mem[88671] = 16'b0000000000000000;
	sram_mem[88672] = 16'b0000000000000000;
	sram_mem[88673] = 16'b0000000000000000;
	sram_mem[88674] = 16'b0000000000000000;
	sram_mem[88675] = 16'b0000000000000000;
	sram_mem[88676] = 16'b0000000000000000;
	sram_mem[88677] = 16'b0000000000000000;
	sram_mem[88678] = 16'b0000000000000000;
	sram_mem[88679] = 16'b0000000000000000;
	sram_mem[88680] = 16'b0000000000000000;
	sram_mem[88681] = 16'b0000000000000000;
	sram_mem[88682] = 16'b0000000000000000;
	sram_mem[88683] = 16'b0000000000000000;
	sram_mem[88684] = 16'b0000000000000000;
	sram_mem[88685] = 16'b0000000000000000;
	sram_mem[88686] = 16'b0000000000000000;
	sram_mem[88687] = 16'b0000000000000000;
	sram_mem[88688] = 16'b0000000000000000;
	sram_mem[88689] = 16'b0000000000000000;
	sram_mem[88690] = 16'b0000000000000000;
	sram_mem[88691] = 16'b0000000000000000;
	sram_mem[88692] = 16'b0000000000000000;
	sram_mem[88693] = 16'b0000000000000000;
	sram_mem[88694] = 16'b0000000000000000;
	sram_mem[88695] = 16'b0000000000000000;
	sram_mem[88696] = 16'b0000000000000000;
	sram_mem[88697] = 16'b0000000000000000;
	sram_mem[88698] = 16'b0000000000000000;
	sram_mem[88699] = 16'b0000000000000000;
	sram_mem[88700] = 16'b0000000000000000;
	sram_mem[88701] = 16'b0000000000000000;
	sram_mem[88702] = 16'b0000000000000000;
	sram_mem[88703] = 16'b0000000000000000;
	sram_mem[88704] = 16'b0000000000000000;
	sram_mem[88705] = 16'b0000000000000000;
	sram_mem[88706] = 16'b0000000000000000;
	sram_mem[88707] = 16'b0000000000000000;
	sram_mem[88708] = 16'b0000000000000000;
	sram_mem[88709] = 16'b0000000000000000;
	sram_mem[88710] = 16'b0000000000000000;
	sram_mem[88711] = 16'b0000000000000000;
	sram_mem[88712] = 16'b0000000000000000;
	sram_mem[88713] = 16'b0000000000000000;
	sram_mem[88714] = 16'b0000000000000000;
	sram_mem[88715] = 16'b0000000000000000;
	sram_mem[88716] = 16'b0000000000000000;
	sram_mem[88717] = 16'b0000000000000000;
	sram_mem[88718] = 16'b0000000000000000;
	sram_mem[88719] = 16'b0000000000000000;
	sram_mem[88720] = 16'b0000000000000000;
	sram_mem[88721] = 16'b0000000000000000;
	sram_mem[88722] = 16'b0000000000000000;
	sram_mem[88723] = 16'b0000000000000000;
	sram_mem[88724] = 16'b0000000000000000;
	sram_mem[88725] = 16'b0000000000000000;
	sram_mem[88726] = 16'b0000000000000000;
	sram_mem[88727] = 16'b0000000000000000;
	sram_mem[88728] = 16'b0000000000000000;
	sram_mem[88729] = 16'b0000000000000000;
	sram_mem[88730] = 16'b0000000000000000;
	sram_mem[88731] = 16'b0000000000000000;
	sram_mem[88732] = 16'b0000000000000000;
	sram_mem[88733] = 16'b0000000000000000;
	sram_mem[88734] = 16'b0000000000000000;
	sram_mem[88735] = 16'b0000000000000000;
	sram_mem[88736] = 16'b0000000000000000;
	sram_mem[88737] = 16'b0000000000000000;
	sram_mem[88738] = 16'b0000000000000000;
	sram_mem[88739] = 16'b0000000000000000;
	sram_mem[88740] = 16'b0000000000000000;
	sram_mem[88741] = 16'b0000000000000000;
	sram_mem[88742] = 16'b0000000000000000;
	sram_mem[88743] = 16'b0000000000000000;
	sram_mem[88744] = 16'b0000000000000000;
	sram_mem[88745] = 16'b0000000000000000;
	sram_mem[88746] = 16'b0000000000000000;
	sram_mem[88747] = 16'b0000000000000000;
	sram_mem[88748] = 16'b0000000000000000;
	sram_mem[88749] = 16'b0000000000000000;
	sram_mem[88750] = 16'b0000000000000000;
	sram_mem[88751] = 16'b0000000000000000;
	sram_mem[88752] = 16'b0000000000000000;
	sram_mem[88753] = 16'b0000000000000000;
	sram_mem[88754] = 16'b0000000000000000;
	sram_mem[88755] = 16'b0000000000000000;
	sram_mem[88756] = 16'b0000000000000000;
	sram_mem[88757] = 16'b0000000000000000;
	sram_mem[88758] = 16'b0000000000000000;
	sram_mem[88759] = 16'b0000000000000000;
	sram_mem[88760] = 16'b0000000000000000;
	sram_mem[88761] = 16'b0000000000000000;
	sram_mem[88762] = 16'b0000000000000000;
	sram_mem[88763] = 16'b0000000000000000;
	sram_mem[88764] = 16'b0000000000000000;
	sram_mem[88765] = 16'b0000000000000000;
	sram_mem[88766] = 16'b0000000000000000;
	sram_mem[88767] = 16'b0000000000000000;
	sram_mem[88768] = 16'b0000000000000000;
	sram_mem[88769] = 16'b0000000000000000;
	sram_mem[88770] = 16'b0000000000000000;
	sram_mem[88771] = 16'b0000000000000000;
	sram_mem[88772] = 16'b0000000000000000;
	sram_mem[88773] = 16'b0000000000000000;
	sram_mem[88774] = 16'b0000000000000000;
	sram_mem[88775] = 16'b0000000000000000;
	sram_mem[88776] = 16'b0000000000000000;
	sram_mem[88777] = 16'b0000000000000000;
	sram_mem[88778] = 16'b0000000000000000;
	sram_mem[88779] = 16'b0000000000000000;
	sram_mem[88780] = 16'b0000000000000000;
	sram_mem[88781] = 16'b0000000000000000;
	sram_mem[88782] = 16'b0000000000000000;
	sram_mem[88783] = 16'b0000000000000000;
	sram_mem[88784] = 16'b0000000000000000;
	sram_mem[88785] = 16'b0000000000000000;
	sram_mem[88786] = 16'b0000000000000000;
	sram_mem[88787] = 16'b0000000000000000;
	sram_mem[88788] = 16'b0000000000000000;
	sram_mem[88789] = 16'b0000000000000000;
	sram_mem[88790] = 16'b0000000000000000;
	sram_mem[88791] = 16'b0000000000000000;
	sram_mem[88792] = 16'b0000000000000000;
	sram_mem[88793] = 16'b0000000000000000;
	sram_mem[88794] = 16'b0000000000000000;
	sram_mem[88795] = 16'b0000000000000000;
	sram_mem[88796] = 16'b0000000000000000;
	sram_mem[88797] = 16'b0000000000000000;
	sram_mem[88798] = 16'b0000000000000000;
	sram_mem[88799] = 16'b0000000000000000;
	sram_mem[88800] = 16'b0000000000000000;
	sram_mem[88801] = 16'b0000000000000000;
	sram_mem[88802] = 16'b0000000000000000;
	sram_mem[88803] = 16'b0000000000000000;
	sram_mem[88804] = 16'b0000000000000000;
	sram_mem[88805] = 16'b0000000000000000;
	sram_mem[88806] = 16'b0000000000000000;
	sram_mem[88807] = 16'b0000000000000000;
	sram_mem[88808] = 16'b0000000000000000;
	sram_mem[88809] = 16'b0000000000000000;
	sram_mem[88810] = 16'b0000000000000000;
	sram_mem[88811] = 16'b0000000000000000;
	sram_mem[88812] = 16'b0000000000000000;
	sram_mem[88813] = 16'b0000000000000000;
	sram_mem[88814] = 16'b0000000000000000;
	sram_mem[88815] = 16'b0000000000000000;
	sram_mem[88816] = 16'b0000000000000000;
	sram_mem[88817] = 16'b0000000000000000;
	sram_mem[88818] = 16'b0000000000000000;
	sram_mem[88819] = 16'b0000000000000000;
	sram_mem[88820] = 16'b0000000000000000;
	sram_mem[88821] = 16'b0000000000000000;
	sram_mem[88822] = 16'b0000000000000000;
	sram_mem[88823] = 16'b0000000000000000;
	sram_mem[88824] = 16'b0000000000000000;
	sram_mem[88825] = 16'b0000000000000000;
	sram_mem[88826] = 16'b0000000000000000;
	sram_mem[88827] = 16'b0000000000000000;
	sram_mem[88828] = 16'b0000000000000000;
	sram_mem[88829] = 16'b0000000000000000;
	sram_mem[88830] = 16'b0000000000000000;
	sram_mem[88831] = 16'b0000000000000000;
	sram_mem[88832] = 16'b0000000000000000;
	sram_mem[88833] = 16'b0000000000000000;
	sram_mem[88834] = 16'b0000000000000000;
	sram_mem[88835] = 16'b0000000000000000;
	sram_mem[88836] = 16'b0000000000000000;
	sram_mem[88837] = 16'b0000000000000000;
	sram_mem[88838] = 16'b0000000000000000;
	sram_mem[88839] = 16'b0000000000000000;
	sram_mem[88840] = 16'b0000000000000000;
	sram_mem[88841] = 16'b0000000000000000;
	sram_mem[88842] = 16'b0000000000000000;
	sram_mem[88843] = 16'b0000000000000000;
	sram_mem[88844] = 16'b0000000000000000;
	sram_mem[88845] = 16'b0000000000000000;
	sram_mem[88846] = 16'b0000000000000000;
	sram_mem[88847] = 16'b0000000000000000;
	sram_mem[88848] = 16'b0000000000000000;
	sram_mem[88849] = 16'b0000000000000000;
	sram_mem[88850] = 16'b0000000000000000;
	sram_mem[88851] = 16'b0000000000000000;
	sram_mem[88852] = 16'b0000000000000000;
	sram_mem[88853] = 16'b0000000000000000;
	sram_mem[88854] = 16'b0000000000000000;
	sram_mem[88855] = 16'b0000000000000000;
	sram_mem[88856] = 16'b0000000000000000;
	sram_mem[88857] = 16'b0000000000000000;
	sram_mem[88858] = 16'b0000000000000000;
	sram_mem[88859] = 16'b0000000000000000;
	sram_mem[88860] = 16'b0000000000000000;
	sram_mem[88861] = 16'b0000000000000000;
	sram_mem[88862] = 16'b0000000000000000;
	sram_mem[88863] = 16'b0000000000000000;
	sram_mem[88864] = 16'b0000000000000000;
	sram_mem[88865] = 16'b0000000000000000;
	sram_mem[88866] = 16'b0000000000000000;
	sram_mem[88867] = 16'b0000000000000000;
	sram_mem[88868] = 16'b0000000000000000;
	sram_mem[88869] = 16'b0000000000000000;
	sram_mem[88870] = 16'b0000000000000000;
	sram_mem[88871] = 16'b0000000000000000;
	sram_mem[88872] = 16'b0000000000000000;
	sram_mem[88873] = 16'b0000000000000000;
	sram_mem[88874] = 16'b0000000000000000;
	sram_mem[88875] = 16'b0000000000000000;
	sram_mem[88876] = 16'b0000000000000000;
	sram_mem[88877] = 16'b0000000000000000;
	sram_mem[88878] = 16'b0000000000000000;
	sram_mem[88879] = 16'b0000000000000000;
	sram_mem[88880] = 16'b0000000000000000;
	sram_mem[88881] = 16'b0000000000000000;
	sram_mem[88882] = 16'b0000000000000000;
	sram_mem[88883] = 16'b0000000000000000;
	sram_mem[88884] = 16'b0000000000000000;
	sram_mem[88885] = 16'b0000000000000000;
	sram_mem[88886] = 16'b0000000000000000;
	sram_mem[88887] = 16'b0000000000000000;
	sram_mem[88888] = 16'b0000000000000000;
	sram_mem[88889] = 16'b0000000000000000;
	sram_mem[88890] = 16'b0000000000000000;
	sram_mem[88891] = 16'b0000000000000000;
	sram_mem[88892] = 16'b0000000000000000;
	sram_mem[88893] = 16'b0000000000000000;
	sram_mem[88894] = 16'b0000000000000000;
	sram_mem[88895] = 16'b0000000000000000;
	sram_mem[88896] = 16'b0000000000000000;
	sram_mem[88897] = 16'b0000000000000000;
	sram_mem[88898] = 16'b0000000000000000;
	sram_mem[88899] = 16'b0000000000000000;
	sram_mem[88900] = 16'b0000000000000000;
	sram_mem[88901] = 16'b0000000000000000;
	sram_mem[88902] = 16'b0000000000000000;
	sram_mem[88903] = 16'b0000000000000000;
	sram_mem[88904] = 16'b0000000000000000;
	sram_mem[88905] = 16'b0000000000000000;
	sram_mem[88906] = 16'b0000000000000000;
	sram_mem[88907] = 16'b0000000000000000;
	sram_mem[88908] = 16'b0000000000000000;
	sram_mem[88909] = 16'b0000000000000000;
	sram_mem[88910] = 16'b0000000000000000;
	sram_mem[88911] = 16'b0000000000000000;
	sram_mem[88912] = 16'b0000000000000000;
	sram_mem[88913] = 16'b0000000000000000;
	sram_mem[88914] = 16'b0000000000000000;
	sram_mem[88915] = 16'b0000000000000000;
	sram_mem[88916] = 16'b0000000000000000;
	sram_mem[88917] = 16'b0000000000000000;
	sram_mem[88918] = 16'b0000000000000000;
	sram_mem[88919] = 16'b0000000000000000;
	sram_mem[88920] = 16'b0000000000000000;
	sram_mem[88921] = 16'b0000000000000000;
	sram_mem[88922] = 16'b0000000000000000;
	sram_mem[88923] = 16'b0000000000000000;
	sram_mem[88924] = 16'b0000000000000000;
	sram_mem[88925] = 16'b0000000000000000;
	sram_mem[88926] = 16'b0000000000000000;
	sram_mem[88927] = 16'b0000000000000000;
	sram_mem[88928] = 16'b0000000000000000;
	sram_mem[88929] = 16'b0000000000000000;
	sram_mem[88930] = 16'b0000000000000000;
	sram_mem[88931] = 16'b0000000000000000;
	sram_mem[88932] = 16'b0000000000000000;
	sram_mem[88933] = 16'b0000000000000000;
	sram_mem[88934] = 16'b0000000000000000;
	sram_mem[88935] = 16'b0000000000000000;
	sram_mem[88936] = 16'b0000000000000000;
	sram_mem[88937] = 16'b0000000000000000;
	sram_mem[88938] = 16'b0000000000000000;
	sram_mem[88939] = 16'b0000000000000000;
	sram_mem[88940] = 16'b0000000000000000;
	sram_mem[88941] = 16'b0000000000000000;
	sram_mem[88942] = 16'b0000000000000000;
	sram_mem[88943] = 16'b0000000000000000;
	sram_mem[88944] = 16'b0000000000000000;
	sram_mem[88945] = 16'b0000000000000000;
	sram_mem[88946] = 16'b0000000000000000;
	sram_mem[88947] = 16'b0000000000000000;
	sram_mem[88948] = 16'b0000000000000000;
	sram_mem[88949] = 16'b0000000000000000;
	sram_mem[88950] = 16'b0000000000000000;
	sram_mem[88951] = 16'b0000000000000000;
	sram_mem[88952] = 16'b0000000000000000;
	sram_mem[88953] = 16'b0000000000000000;
	sram_mem[88954] = 16'b0000000000000000;
	sram_mem[88955] = 16'b0000000000000000;
	sram_mem[88956] = 16'b0000000000000000;
	sram_mem[88957] = 16'b0000000000000000;
	sram_mem[88958] = 16'b0000000000000000;
	sram_mem[88959] = 16'b0000000000000000;
	sram_mem[88960] = 16'b0000000000000000;
	sram_mem[88961] = 16'b0000000000000000;
	sram_mem[88962] = 16'b0000000000000000;
	sram_mem[88963] = 16'b0000000000000000;
	sram_mem[88964] = 16'b0000000000000000;
	sram_mem[88965] = 16'b0000000000000000;
	sram_mem[88966] = 16'b0000000000000000;
	sram_mem[88967] = 16'b0000000000000000;
	sram_mem[88968] = 16'b0000000000000000;
	sram_mem[88969] = 16'b0000000000000000;
	sram_mem[88970] = 16'b0000000000000000;
	sram_mem[88971] = 16'b0000000000000000;
	sram_mem[88972] = 16'b0000000000000000;
	sram_mem[88973] = 16'b0000000000000000;
	sram_mem[88974] = 16'b0000000000000000;
	sram_mem[88975] = 16'b0000000000000000;
	sram_mem[88976] = 16'b0000000000000000;
	sram_mem[88977] = 16'b0000000000000000;
	sram_mem[88978] = 16'b0000000000000000;
	sram_mem[88979] = 16'b0000000000000000;
	sram_mem[88980] = 16'b0000000000000000;
	sram_mem[88981] = 16'b0000000000000000;
	sram_mem[88982] = 16'b0000000000000000;
	sram_mem[88983] = 16'b0000000000000000;
	sram_mem[88984] = 16'b0000000000000000;
	sram_mem[88985] = 16'b0000000000000000;
	sram_mem[88986] = 16'b0000000000000000;
	sram_mem[88987] = 16'b0000000000000000;
	sram_mem[88988] = 16'b0000000000000000;
	sram_mem[88989] = 16'b0000000000000000;
	sram_mem[88990] = 16'b0000000000000000;
	sram_mem[88991] = 16'b0000000000000000;
	sram_mem[88992] = 16'b0000000000000000;
	sram_mem[88993] = 16'b0000000000000000;
	sram_mem[88994] = 16'b0000000000000000;
	sram_mem[88995] = 16'b0000000000000000;
	sram_mem[88996] = 16'b0000000000000000;
	sram_mem[88997] = 16'b0000000000000000;
	sram_mem[88998] = 16'b0000000000000000;
	sram_mem[88999] = 16'b0000000000000000;
	sram_mem[89000] = 16'b0000000000000000;
	sram_mem[89001] = 16'b0000000000000000;
	sram_mem[89002] = 16'b0000000000000000;
	sram_mem[89003] = 16'b0000000000000000;
	sram_mem[89004] = 16'b0000000000000000;
	sram_mem[89005] = 16'b0000000000000000;
	sram_mem[89006] = 16'b0000000000000000;
	sram_mem[89007] = 16'b0000000000000000;
	sram_mem[89008] = 16'b0000000000000000;
	sram_mem[89009] = 16'b0000000000000000;
	sram_mem[89010] = 16'b0000000000000000;
	sram_mem[89011] = 16'b0000000000000000;
	sram_mem[89012] = 16'b0000000000000000;
	sram_mem[89013] = 16'b0000000000000000;
	sram_mem[89014] = 16'b0000000000000000;
	sram_mem[89015] = 16'b0000000000000000;
	sram_mem[89016] = 16'b0000000000000000;
	sram_mem[89017] = 16'b0000000000000000;
	sram_mem[89018] = 16'b0000000000000000;
	sram_mem[89019] = 16'b0000000000000000;
	sram_mem[89020] = 16'b0000000000000000;
	sram_mem[89021] = 16'b0000000000000000;
	sram_mem[89022] = 16'b0000000000000000;
	sram_mem[89023] = 16'b0000000000000000;
	sram_mem[89024] = 16'b0000000000000000;
	sram_mem[89025] = 16'b0000000000000000;
	sram_mem[89026] = 16'b0000000000000000;
	sram_mem[89027] = 16'b0000000000000000;
	sram_mem[89028] = 16'b0000000000000000;
	sram_mem[89029] = 16'b0000000000000000;
	sram_mem[89030] = 16'b0000000000000000;
	sram_mem[89031] = 16'b0000000000000000;
	sram_mem[89032] = 16'b0000000000000000;
	sram_mem[89033] = 16'b0000000000000000;
	sram_mem[89034] = 16'b0000000000000000;
	sram_mem[89035] = 16'b0000000000000000;
	sram_mem[89036] = 16'b0000000000000000;
	sram_mem[89037] = 16'b0000000000000000;
	sram_mem[89038] = 16'b0000000000000000;
	sram_mem[89039] = 16'b0000000000000000;
	sram_mem[89040] = 16'b0000000000000000;
	sram_mem[89041] = 16'b0000000000000000;
	sram_mem[89042] = 16'b0000000000000000;
	sram_mem[89043] = 16'b0000000000000000;
	sram_mem[89044] = 16'b0000000000000000;
	sram_mem[89045] = 16'b0000000000000000;
	sram_mem[89046] = 16'b0000000000000000;
	sram_mem[89047] = 16'b0000000000000000;
	sram_mem[89048] = 16'b0000000000000000;
	sram_mem[89049] = 16'b0000000000000000;
	sram_mem[89050] = 16'b0000000000000000;
	sram_mem[89051] = 16'b0000000000000000;
	sram_mem[89052] = 16'b0000000000000000;
	sram_mem[89053] = 16'b0000000000000000;
	sram_mem[89054] = 16'b0000000000000000;
	sram_mem[89055] = 16'b0000000000000000;
	sram_mem[89056] = 16'b0000000000000000;
	sram_mem[89057] = 16'b0000000000000000;
	sram_mem[89058] = 16'b0000000000000000;
	sram_mem[89059] = 16'b0000000000000000;
	sram_mem[89060] = 16'b0000000000000000;
	sram_mem[89061] = 16'b0000000000000000;
	sram_mem[89062] = 16'b0000000000000000;
	sram_mem[89063] = 16'b0000000000000000;
	sram_mem[89064] = 16'b0000000000000000;
	sram_mem[89065] = 16'b0000000000000000;
	sram_mem[89066] = 16'b0000000000000000;
	sram_mem[89067] = 16'b0000000000000000;
	sram_mem[89068] = 16'b0000000000000000;
	sram_mem[89069] = 16'b0000000000000000;
	sram_mem[89070] = 16'b0000000000000000;
	sram_mem[89071] = 16'b0000000000000000;
	sram_mem[89072] = 16'b0000000000000000;
	sram_mem[89073] = 16'b0000000000000000;
	sram_mem[89074] = 16'b0000000000000000;
	sram_mem[89075] = 16'b0000000000000000;
	sram_mem[89076] = 16'b0000000000000000;
	sram_mem[89077] = 16'b0000000000000000;
	sram_mem[89078] = 16'b0000000000000000;
	sram_mem[89079] = 16'b0000000000000000;
	sram_mem[89080] = 16'b0000000000000000;
	sram_mem[89081] = 16'b0000000000000000;
	sram_mem[89082] = 16'b0000000000000000;
	sram_mem[89083] = 16'b0000000000000000;
	sram_mem[89084] = 16'b0000000000000000;
	sram_mem[89085] = 16'b0000000000000000;
	sram_mem[89086] = 16'b0000000000000000;
	sram_mem[89087] = 16'b0000000000000000;
	sram_mem[89088] = 16'b0000000000000000;
	sram_mem[89089] = 16'b0000000000000000;
	sram_mem[89090] = 16'b0000000000000000;
	sram_mem[89091] = 16'b0000000000000000;
	sram_mem[89092] = 16'b0000000000000000;
	sram_mem[89093] = 16'b0000000000000000;
	sram_mem[89094] = 16'b0000000000000000;
	sram_mem[89095] = 16'b0000000000000000;
	sram_mem[89096] = 16'b0000000000000000;
	sram_mem[89097] = 16'b0000000000000000;
	sram_mem[89098] = 16'b0000000000000000;
	sram_mem[89099] = 16'b0000000000000000;
	sram_mem[89100] = 16'b0000000000000000;
	sram_mem[89101] = 16'b0000000000000000;
	sram_mem[89102] = 16'b0000000000000000;
	sram_mem[89103] = 16'b0000000000000000;
	sram_mem[89104] = 16'b0000000000000000;
	sram_mem[89105] = 16'b0000000000000000;
	sram_mem[89106] = 16'b0000000000000000;
	sram_mem[89107] = 16'b0000000000000000;
	sram_mem[89108] = 16'b0000000000000000;
	sram_mem[89109] = 16'b0000000000000000;
	sram_mem[89110] = 16'b0000000000000000;
	sram_mem[89111] = 16'b0000000000000000;
	sram_mem[89112] = 16'b0000000000000000;
	sram_mem[89113] = 16'b0000000000000000;
	sram_mem[89114] = 16'b0000000000000000;
	sram_mem[89115] = 16'b0000000000000000;
	sram_mem[89116] = 16'b0000000000000000;
	sram_mem[89117] = 16'b0000000000000000;
	sram_mem[89118] = 16'b0000000000000000;
	sram_mem[89119] = 16'b0000000000000000;
	sram_mem[89120] = 16'b0000000000000000;
	sram_mem[89121] = 16'b0000000000000000;
	sram_mem[89122] = 16'b0000000000000000;
	sram_mem[89123] = 16'b0000000000000000;
	sram_mem[89124] = 16'b0000000000000000;
	sram_mem[89125] = 16'b0000000000000000;
	sram_mem[89126] = 16'b0000000000000000;
	sram_mem[89127] = 16'b0000000000000000;
	sram_mem[89128] = 16'b0000000000000000;
	sram_mem[89129] = 16'b0000000000000000;
	sram_mem[89130] = 16'b0000000000000000;
	sram_mem[89131] = 16'b0000000000000000;
	sram_mem[89132] = 16'b0000000000000000;
	sram_mem[89133] = 16'b0000000000000000;
	sram_mem[89134] = 16'b0000000000000000;
	sram_mem[89135] = 16'b0000000000000000;
	sram_mem[89136] = 16'b0000000000000000;
	sram_mem[89137] = 16'b0000000000000000;
	sram_mem[89138] = 16'b0000000000000000;
	sram_mem[89139] = 16'b0000000000000000;
	sram_mem[89140] = 16'b0000000000000000;
	sram_mem[89141] = 16'b0000000000000000;
	sram_mem[89142] = 16'b0000000000000000;
	sram_mem[89143] = 16'b0000000000000000;
	sram_mem[89144] = 16'b0000000000000000;
	sram_mem[89145] = 16'b0000000000000000;
	sram_mem[89146] = 16'b0000000000000000;
	sram_mem[89147] = 16'b0000000000000000;
	sram_mem[89148] = 16'b0000000000000000;
	sram_mem[89149] = 16'b0000000000000000;
	sram_mem[89150] = 16'b0000000000000000;
	sram_mem[89151] = 16'b0000000000000000;
	sram_mem[89152] = 16'b0000000000000000;
	sram_mem[89153] = 16'b0000000000000000;
	sram_mem[89154] = 16'b0000000000000000;
	sram_mem[89155] = 16'b0000000000000000;
	sram_mem[89156] = 16'b0000000000000000;
	sram_mem[89157] = 16'b0000000000000000;
	sram_mem[89158] = 16'b0000000000000000;
	sram_mem[89159] = 16'b0000000000000000;
	sram_mem[89160] = 16'b0000000000000000;
	sram_mem[89161] = 16'b0000000000000000;
	sram_mem[89162] = 16'b0000000000000000;
	sram_mem[89163] = 16'b0000000000000000;
	sram_mem[89164] = 16'b0000000000000000;
	sram_mem[89165] = 16'b0000000000000000;
	sram_mem[89166] = 16'b0000000000000000;
	sram_mem[89167] = 16'b0000000000000000;
	sram_mem[89168] = 16'b0000000000000000;
	sram_mem[89169] = 16'b0000000000000000;
	sram_mem[89170] = 16'b0000000000000000;
	sram_mem[89171] = 16'b0000000000000000;
	sram_mem[89172] = 16'b0000000000000000;
	sram_mem[89173] = 16'b0000000000000000;
	sram_mem[89174] = 16'b0000000000000000;
	sram_mem[89175] = 16'b0000000000000000;
	sram_mem[89176] = 16'b0000000000000000;
	sram_mem[89177] = 16'b0000000000000000;
	sram_mem[89178] = 16'b0000000000000000;
	sram_mem[89179] = 16'b0000000000000000;
	sram_mem[89180] = 16'b0000000000000000;
	sram_mem[89181] = 16'b0000000000000000;
	sram_mem[89182] = 16'b0000000000000000;
	sram_mem[89183] = 16'b0000000000000000;
	sram_mem[89184] = 16'b0000000000000000;
	sram_mem[89185] = 16'b0000000000000000;
	sram_mem[89186] = 16'b0000000000000000;
	sram_mem[89187] = 16'b0000000000000000;
	sram_mem[89188] = 16'b0000000000000000;
	sram_mem[89189] = 16'b0000000000000000;
	sram_mem[89190] = 16'b0000000000000000;
	sram_mem[89191] = 16'b0000000000000000;
	sram_mem[89192] = 16'b0000000000000000;
	sram_mem[89193] = 16'b0000000000000000;
	sram_mem[89194] = 16'b0000000000000000;
	sram_mem[89195] = 16'b0000000000000000;
	sram_mem[89196] = 16'b0000000000000000;
	sram_mem[89197] = 16'b0000000000000000;
	sram_mem[89198] = 16'b0000000000000000;
	sram_mem[89199] = 16'b0000000000000000;
	sram_mem[89200] = 16'b0000000000000000;
	sram_mem[89201] = 16'b0000000000000000;
	sram_mem[89202] = 16'b0000000000000000;
	sram_mem[89203] = 16'b0000000000000000;
	sram_mem[89204] = 16'b0000000000000000;
	sram_mem[89205] = 16'b0000000000000000;
	sram_mem[89206] = 16'b0000000000000000;
	sram_mem[89207] = 16'b0000000000000000;
	sram_mem[89208] = 16'b0000000000000000;
	sram_mem[89209] = 16'b0000000000000000;
	sram_mem[89210] = 16'b0000000000000000;
	sram_mem[89211] = 16'b0000000000000000;
	sram_mem[89212] = 16'b0000000000000000;
	sram_mem[89213] = 16'b0000000000000000;
	sram_mem[89214] = 16'b0000000000000000;
	sram_mem[89215] = 16'b0000000000000000;
	sram_mem[89216] = 16'b0000000000000000;
	sram_mem[89217] = 16'b0000000000000000;
	sram_mem[89218] = 16'b0000000000000000;
	sram_mem[89219] = 16'b0000000000000000;
	sram_mem[89220] = 16'b0000000000000000;
	sram_mem[89221] = 16'b0000000000000000;
	sram_mem[89222] = 16'b0000000000000000;
	sram_mem[89223] = 16'b0000000000000000;
	sram_mem[89224] = 16'b0000000000000000;
	sram_mem[89225] = 16'b0000000000000000;
	sram_mem[89226] = 16'b0000000000000000;
	sram_mem[89227] = 16'b0000000000000000;
	sram_mem[89228] = 16'b0000000000000000;
	sram_mem[89229] = 16'b0000000000000000;
	sram_mem[89230] = 16'b0000000000000000;
	sram_mem[89231] = 16'b0000000000000000;
	sram_mem[89232] = 16'b0000000000000000;
	sram_mem[89233] = 16'b0000000000000000;
	sram_mem[89234] = 16'b0000000000000000;
	sram_mem[89235] = 16'b0000000000000000;
	sram_mem[89236] = 16'b0000000000000000;
	sram_mem[89237] = 16'b0000000000000000;
	sram_mem[89238] = 16'b0000000000000000;
	sram_mem[89239] = 16'b0000000000000000;
	sram_mem[89240] = 16'b0000000000000000;
	sram_mem[89241] = 16'b0000000000000000;
	sram_mem[89242] = 16'b0000000000000000;
	sram_mem[89243] = 16'b0000000000000000;
	sram_mem[89244] = 16'b0000000000000000;
	sram_mem[89245] = 16'b0000000000000000;
	sram_mem[89246] = 16'b0000000000000000;
	sram_mem[89247] = 16'b0000000000000000;
	sram_mem[89248] = 16'b0000000000000000;
	sram_mem[89249] = 16'b0000000000000000;
	sram_mem[89250] = 16'b0000000000000000;
	sram_mem[89251] = 16'b0000000000000000;
	sram_mem[89252] = 16'b0000000000000000;
	sram_mem[89253] = 16'b0000000000000000;
	sram_mem[89254] = 16'b0000000000000000;
	sram_mem[89255] = 16'b0000000000000000;
	sram_mem[89256] = 16'b0000000000000000;
	sram_mem[89257] = 16'b0000000000000000;
	sram_mem[89258] = 16'b0000000000000000;
	sram_mem[89259] = 16'b0000000000000000;
	sram_mem[89260] = 16'b0000000000000000;
	sram_mem[89261] = 16'b0000000000000000;
	sram_mem[89262] = 16'b0000000000000000;
	sram_mem[89263] = 16'b0000000000000000;
	sram_mem[89264] = 16'b0000000000000000;
	sram_mem[89265] = 16'b0000000000000000;
	sram_mem[89266] = 16'b0000000000000000;
	sram_mem[89267] = 16'b0000000000000000;
	sram_mem[89268] = 16'b0000000000000000;
	sram_mem[89269] = 16'b0000000000000000;
	sram_mem[89270] = 16'b0000000000000000;
	sram_mem[89271] = 16'b0000000000000000;
	sram_mem[89272] = 16'b0000000000000000;
	sram_mem[89273] = 16'b0000000000000000;
	sram_mem[89274] = 16'b0000000000000000;
	sram_mem[89275] = 16'b0000000000000000;
	sram_mem[89276] = 16'b0000000000000000;
	sram_mem[89277] = 16'b0000000000000000;
	sram_mem[89278] = 16'b0000000000000000;
	sram_mem[89279] = 16'b0000000000000000;
	sram_mem[89280] = 16'b0000000000000000;
	sram_mem[89281] = 16'b0000000000000000;
	sram_mem[89282] = 16'b0000000000000000;
	sram_mem[89283] = 16'b0000000000000000;
	sram_mem[89284] = 16'b0000000000000000;
	sram_mem[89285] = 16'b0000000000000000;
	sram_mem[89286] = 16'b0000000000000000;
	sram_mem[89287] = 16'b0000000000000000;
	sram_mem[89288] = 16'b0000000000000000;
	sram_mem[89289] = 16'b0000000000000000;
	sram_mem[89290] = 16'b0000000000000000;
	sram_mem[89291] = 16'b0000000000000000;
	sram_mem[89292] = 16'b0000000000000000;
	sram_mem[89293] = 16'b0000000000000000;
	sram_mem[89294] = 16'b0000000000000000;
	sram_mem[89295] = 16'b0000000000000000;
	sram_mem[89296] = 16'b0000000000000000;
	sram_mem[89297] = 16'b0000000000000000;
	sram_mem[89298] = 16'b0000000000000000;
	sram_mem[89299] = 16'b0000000000000000;
	sram_mem[89300] = 16'b0000000000000000;
	sram_mem[89301] = 16'b0000000000000000;
	sram_mem[89302] = 16'b0000000000000000;
	sram_mem[89303] = 16'b0000000000000000;
	sram_mem[89304] = 16'b0000000000000000;
	sram_mem[89305] = 16'b0000000000000000;
	sram_mem[89306] = 16'b0000000000000000;
	sram_mem[89307] = 16'b0000000000000000;
	sram_mem[89308] = 16'b0000000000000000;
	sram_mem[89309] = 16'b0000000000000000;
	sram_mem[89310] = 16'b0000000000000000;
	sram_mem[89311] = 16'b0000000000000000;
	sram_mem[89312] = 16'b0000000000000000;
	sram_mem[89313] = 16'b0000000000000000;
	sram_mem[89314] = 16'b0000000000000000;
	sram_mem[89315] = 16'b0000000000000000;
	sram_mem[89316] = 16'b0000000000000000;
	sram_mem[89317] = 16'b0000000000000000;
	sram_mem[89318] = 16'b0000000000000000;
	sram_mem[89319] = 16'b0000000000000000;
	sram_mem[89320] = 16'b0000000000000000;
	sram_mem[89321] = 16'b0000000000000000;
	sram_mem[89322] = 16'b0000000000000000;
	sram_mem[89323] = 16'b0000000000000000;
	sram_mem[89324] = 16'b0000000000000000;
	sram_mem[89325] = 16'b0000000000000000;
	sram_mem[89326] = 16'b0000000000000000;
	sram_mem[89327] = 16'b0000000000000000;
	sram_mem[89328] = 16'b0000000000000000;
	sram_mem[89329] = 16'b0000000000000000;
	sram_mem[89330] = 16'b0000000000000000;
	sram_mem[89331] = 16'b0000000000000000;
	sram_mem[89332] = 16'b0000000000000000;
	sram_mem[89333] = 16'b0000000000000000;
	sram_mem[89334] = 16'b0000000000000000;
	sram_mem[89335] = 16'b0000000000000000;
	sram_mem[89336] = 16'b0000000000000000;
	sram_mem[89337] = 16'b0000000000000000;
	sram_mem[89338] = 16'b0000000000000000;
	sram_mem[89339] = 16'b0000000000000000;
	sram_mem[89340] = 16'b0000000000000000;
	sram_mem[89341] = 16'b0000000000000000;
	sram_mem[89342] = 16'b0000000000000000;
	sram_mem[89343] = 16'b0000000000000000;
	sram_mem[89344] = 16'b0000000000000000;
	sram_mem[89345] = 16'b0000000000000000;
	sram_mem[89346] = 16'b0000000000000000;
	sram_mem[89347] = 16'b0000000000000000;
	sram_mem[89348] = 16'b0000000000000000;
	sram_mem[89349] = 16'b0000000000000000;
	sram_mem[89350] = 16'b0000000000000000;
	sram_mem[89351] = 16'b0000000000000000;
	sram_mem[89352] = 16'b0000000000000000;
	sram_mem[89353] = 16'b0000000000000000;
	sram_mem[89354] = 16'b0000000000000000;
	sram_mem[89355] = 16'b0000000000000000;
	sram_mem[89356] = 16'b0000000000000000;
	sram_mem[89357] = 16'b0000000000000000;
	sram_mem[89358] = 16'b0000000000000000;
	sram_mem[89359] = 16'b0000000000000000;
	sram_mem[89360] = 16'b0000000000000000;
	sram_mem[89361] = 16'b0000000000000000;
	sram_mem[89362] = 16'b0000000000000000;
	sram_mem[89363] = 16'b0000000000000000;
	sram_mem[89364] = 16'b0000000000000000;
	sram_mem[89365] = 16'b0000000000000000;
	sram_mem[89366] = 16'b0000000000000000;
	sram_mem[89367] = 16'b0000000000000000;
	sram_mem[89368] = 16'b0000000000000000;
	sram_mem[89369] = 16'b0000000000000000;
	sram_mem[89370] = 16'b0000000000000000;
	sram_mem[89371] = 16'b0000000000000000;
	sram_mem[89372] = 16'b0000000000000000;
	sram_mem[89373] = 16'b0000000000000000;
	sram_mem[89374] = 16'b0000000000000000;
	sram_mem[89375] = 16'b0000000000000000;
	sram_mem[89376] = 16'b0000000000000000;
	sram_mem[89377] = 16'b0000000000000000;
	sram_mem[89378] = 16'b0000000000000000;
	sram_mem[89379] = 16'b0000000000000000;
	sram_mem[89380] = 16'b0000000000000000;
	sram_mem[89381] = 16'b0000000000000000;
	sram_mem[89382] = 16'b0000000000000000;
	sram_mem[89383] = 16'b0000000000000000;
	sram_mem[89384] = 16'b0000000000000000;
	sram_mem[89385] = 16'b0000000000000000;
	sram_mem[89386] = 16'b0000000000000000;
	sram_mem[89387] = 16'b0000000000000000;
	sram_mem[89388] = 16'b0000000000000000;
	sram_mem[89389] = 16'b0000000000000000;
	sram_mem[89390] = 16'b0000000000000000;
	sram_mem[89391] = 16'b0000000000000000;
	sram_mem[89392] = 16'b0000000000000000;
	sram_mem[89393] = 16'b0000000000000000;
	sram_mem[89394] = 16'b0000000000000000;
	sram_mem[89395] = 16'b0000000000000000;
	sram_mem[89396] = 16'b0000000000000000;
	sram_mem[89397] = 16'b0000000000000000;
	sram_mem[89398] = 16'b0000000000000000;
	sram_mem[89399] = 16'b0000000000000000;
	sram_mem[89400] = 16'b0000000000000000;
	sram_mem[89401] = 16'b0000000000000000;
	sram_mem[89402] = 16'b0000000000000000;
	sram_mem[89403] = 16'b0000000000000000;
	sram_mem[89404] = 16'b0000000000000000;
	sram_mem[89405] = 16'b0000000000000000;
	sram_mem[89406] = 16'b0000000000000000;
	sram_mem[89407] = 16'b0000000000000000;
	sram_mem[89408] = 16'b0000000000000000;
	sram_mem[89409] = 16'b0000000000000000;
	sram_mem[89410] = 16'b0000000000000000;
	sram_mem[89411] = 16'b0000000000000000;
	sram_mem[89412] = 16'b0000000000000000;
	sram_mem[89413] = 16'b0000000000000000;
	sram_mem[89414] = 16'b0000000000000000;
	sram_mem[89415] = 16'b0000000000000000;
	sram_mem[89416] = 16'b0000000000000000;
	sram_mem[89417] = 16'b0000000000000000;
	sram_mem[89418] = 16'b0000000000000000;
	sram_mem[89419] = 16'b0000000000000000;
	sram_mem[89420] = 16'b0000000000000000;
	sram_mem[89421] = 16'b0000000000000000;
	sram_mem[89422] = 16'b0000000000000000;
	sram_mem[89423] = 16'b0000000000000000;
	sram_mem[89424] = 16'b0000000000000000;
	sram_mem[89425] = 16'b0000000000000000;
	sram_mem[89426] = 16'b0000000000000000;
	sram_mem[89427] = 16'b0000000000000000;
	sram_mem[89428] = 16'b0000000000000000;
	sram_mem[89429] = 16'b0000000000000000;
	sram_mem[89430] = 16'b0000000000000000;
	sram_mem[89431] = 16'b0000000000000000;
	sram_mem[89432] = 16'b0000000000000000;
	sram_mem[89433] = 16'b0000000000000000;
	sram_mem[89434] = 16'b0000000000000000;
	sram_mem[89435] = 16'b0000000000000000;
	sram_mem[89436] = 16'b0000000000000000;
	sram_mem[89437] = 16'b0000000000000000;
	sram_mem[89438] = 16'b0000000000000000;
	sram_mem[89439] = 16'b0000000000000000;
	sram_mem[89440] = 16'b0000000000000000;
	sram_mem[89441] = 16'b0000000000000000;
	sram_mem[89442] = 16'b0000000000000000;
	sram_mem[89443] = 16'b0000000000000000;
	sram_mem[89444] = 16'b0000000000000000;
	sram_mem[89445] = 16'b0000000000000000;
	sram_mem[89446] = 16'b0000000000000000;
	sram_mem[89447] = 16'b0000000000000000;
	sram_mem[89448] = 16'b0000000000000000;
	sram_mem[89449] = 16'b0000000000000000;
	sram_mem[89450] = 16'b0000000000000000;
	sram_mem[89451] = 16'b0000000000000000;
	sram_mem[89452] = 16'b0000000000000000;
	sram_mem[89453] = 16'b0000000000000000;
	sram_mem[89454] = 16'b0000000000000000;
	sram_mem[89455] = 16'b0000000000000000;
	sram_mem[89456] = 16'b0000000000000000;
	sram_mem[89457] = 16'b0000000000000000;
	sram_mem[89458] = 16'b0000000000000000;
	sram_mem[89459] = 16'b0000000000000000;
	sram_mem[89460] = 16'b0000000000000000;
	sram_mem[89461] = 16'b0000000000000000;
	sram_mem[89462] = 16'b0000000000000000;
	sram_mem[89463] = 16'b0000000000000000;
	sram_mem[89464] = 16'b0000000000000000;
	sram_mem[89465] = 16'b0000000000000000;
	sram_mem[89466] = 16'b0000000000000000;
	sram_mem[89467] = 16'b0000000000000000;
	sram_mem[89468] = 16'b0000000000000000;
	sram_mem[89469] = 16'b0000000000000000;
	sram_mem[89470] = 16'b0000000000000000;
	sram_mem[89471] = 16'b0000000000000000;
	sram_mem[89472] = 16'b0000000000000000;
	sram_mem[89473] = 16'b0000000000000000;
	sram_mem[89474] = 16'b0000000000000000;
	sram_mem[89475] = 16'b0000000000000000;
	sram_mem[89476] = 16'b0000000000000000;
	sram_mem[89477] = 16'b0000000000000000;
	sram_mem[89478] = 16'b0000000000000000;
	sram_mem[89479] = 16'b0000000000000000;
	sram_mem[89480] = 16'b0000000000000000;
	sram_mem[89481] = 16'b0000000000000000;
	sram_mem[89482] = 16'b0000000000000000;
	sram_mem[89483] = 16'b0000000000000000;
	sram_mem[89484] = 16'b0000000000000000;
	sram_mem[89485] = 16'b0000000000000000;
	sram_mem[89486] = 16'b0000000000000000;
	sram_mem[89487] = 16'b0000000000000000;
	sram_mem[89488] = 16'b0000000000000000;
	sram_mem[89489] = 16'b0000000000000000;
	sram_mem[89490] = 16'b0000000000000000;
	sram_mem[89491] = 16'b0000000000000000;
	sram_mem[89492] = 16'b0000000000000000;
	sram_mem[89493] = 16'b0000000000000000;
	sram_mem[89494] = 16'b0000000000000000;
	sram_mem[89495] = 16'b0000000000000000;
	sram_mem[89496] = 16'b0000000000000000;
	sram_mem[89497] = 16'b0000000000000000;
	sram_mem[89498] = 16'b0000000000000000;
	sram_mem[89499] = 16'b0000000000000000;
	sram_mem[89500] = 16'b0000000000000000;
	sram_mem[89501] = 16'b0000000000000000;
	sram_mem[89502] = 16'b0000000000000000;
	sram_mem[89503] = 16'b0000000000000000;
	sram_mem[89504] = 16'b0000000000000000;
	sram_mem[89505] = 16'b0000000000000000;
	sram_mem[89506] = 16'b0000000000000000;
	sram_mem[89507] = 16'b0000000000000000;
	sram_mem[89508] = 16'b0000000000000000;
	sram_mem[89509] = 16'b0000000000000000;
	sram_mem[89510] = 16'b0000000000000000;
	sram_mem[89511] = 16'b0000000000000000;
	sram_mem[89512] = 16'b0000000000000000;
	sram_mem[89513] = 16'b0000000000000000;
	sram_mem[89514] = 16'b0000000000000000;
	sram_mem[89515] = 16'b0000000000000000;
	sram_mem[89516] = 16'b0000000000000000;
	sram_mem[89517] = 16'b0000000000000000;
	sram_mem[89518] = 16'b0000000000000000;
	sram_mem[89519] = 16'b0000000000000000;
	sram_mem[89520] = 16'b0000000000000000;
	sram_mem[89521] = 16'b0000000000000000;
	sram_mem[89522] = 16'b0000000000000000;
	sram_mem[89523] = 16'b0000000000000000;
	sram_mem[89524] = 16'b0000000000000000;
	sram_mem[89525] = 16'b0000000000000000;
	sram_mem[89526] = 16'b0000000000000000;
	sram_mem[89527] = 16'b0000000000000000;
	sram_mem[89528] = 16'b0000000000000000;
	sram_mem[89529] = 16'b0000000000000000;
	sram_mem[89530] = 16'b0000000000000000;
	sram_mem[89531] = 16'b0000000000000000;
	sram_mem[89532] = 16'b0000000000000000;
	sram_mem[89533] = 16'b0000000000000000;
	sram_mem[89534] = 16'b0000000000000000;
	sram_mem[89535] = 16'b0000000000000000;
	sram_mem[89536] = 16'b0000000000000000;
	sram_mem[89537] = 16'b0000000000000000;
	sram_mem[89538] = 16'b0000000000000000;
	sram_mem[89539] = 16'b0000000000000000;
	sram_mem[89540] = 16'b0000000000000000;
	sram_mem[89541] = 16'b0000000000000000;
	sram_mem[89542] = 16'b0000000000000000;
	sram_mem[89543] = 16'b0000000000000000;
	sram_mem[89544] = 16'b0000000000000000;
	sram_mem[89545] = 16'b0000000000000000;
	sram_mem[89546] = 16'b0000000000000000;
	sram_mem[89547] = 16'b0000000000000000;
	sram_mem[89548] = 16'b0000000000000000;
	sram_mem[89549] = 16'b0000000000000000;
	sram_mem[89550] = 16'b0000000000000000;
	sram_mem[89551] = 16'b0000000000000000;
	sram_mem[89552] = 16'b0000000000000000;
	sram_mem[89553] = 16'b0000000000000000;
	sram_mem[89554] = 16'b0000000000000000;
	sram_mem[89555] = 16'b0000000000000000;
	sram_mem[89556] = 16'b0000000000000000;
	sram_mem[89557] = 16'b0000000000000000;
	sram_mem[89558] = 16'b0000000000000000;
	sram_mem[89559] = 16'b0000000000000000;
	sram_mem[89560] = 16'b0000000000000000;
	sram_mem[89561] = 16'b0000000000000000;
	sram_mem[89562] = 16'b0000000000000000;
	sram_mem[89563] = 16'b0000000000000000;
	sram_mem[89564] = 16'b0000000000000000;
	sram_mem[89565] = 16'b0000000000000000;
	sram_mem[89566] = 16'b0000000000000000;
	sram_mem[89567] = 16'b0000000000000000;
	sram_mem[89568] = 16'b0000000000000000;
	sram_mem[89569] = 16'b0000000000000000;
	sram_mem[89570] = 16'b0000000000000000;
	sram_mem[89571] = 16'b0000000000000000;
	sram_mem[89572] = 16'b0000000000000000;
	sram_mem[89573] = 16'b0000000000000000;
	sram_mem[89574] = 16'b0000000000000000;
	sram_mem[89575] = 16'b0000000000000000;
	sram_mem[89576] = 16'b0000000000000000;
	sram_mem[89577] = 16'b0000000000000000;
	sram_mem[89578] = 16'b0000000000000000;
	sram_mem[89579] = 16'b0000000000000000;
	sram_mem[89580] = 16'b0000000000000000;
	sram_mem[89581] = 16'b0000000000000000;
	sram_mem[89582] = 16'b0000000000000000;
	sram_mem[89583] = 16'b0000000000000000;
	sram_mem[89584] = 16'b0000000000000000;
	sram_mem[89585] = 16'b0000000000000000;
	sram_mem[89586] = 16'b0000000000000000;
	sram_mem[89587] = 16'b0000000000000000;
	sram_mem[89588] = 16'b0000000000000000;
	sram_mem[89589] = 16'b0000000000000000;
	sram_mem[89590] = 16'b0000000000000000;
	sram_mem[89591] = 16'b0000000000000000;
	sram_mem[89592] = 16'b0000000000000000;
	sram_mem[89593] = 16'b0000000000000000;
	sram_mem[89594] = 16'b0000000000000000;
	sram_mem[89595] = 16'b0000000000000000;
	sram_mem[89596] = 16'b0000000000000000;
	sram_mem[89597] = 16'b0000000000000000;
	sram_mem[89598] = 16'b0000000000000000;
	sram_mem[89599] = 16'b0000000000000000;
	sram_mem[89600] = 16'b0000000000000000;
	sram_mem[89601] = 16'b0000000000000000;
	sram_mem[89602] = 16'b0000000000000000;
	sram_mem[89603] = 16'b0000000000000000;
	sram_mem[89604] = 16'b0000000000000000;
	sram_mem[89605] = 16'b0000000000000000;
	sram_mem[89606] = 16'b0000000000000000;
	sram_mem[89607] = 16'b0000000000000000;
	sram_mem[89608] = 16'b0000000000000000;
	sram_mem[89609] = 16'b0000000000000000;
	sram_mem[89610] = 16'b0000000000000000;
	sram_mem[89611] = 16'b0000000000000000;
	sram_mem[89612] = 16'b0000000000000000;
	sram_mem[89613] = 16'b0000000000000000;
	sram_mem[89614] = 16'b0000000000000000;
	sram_mem[89615] = 16'b0000000000000000;
	sram_mem[89616] = 16'b0000000000000000;
	sram_mem[89617] = 16'b0000000000000000;
	sram_mem[89618] = 16'b0000000000000000;
	sram_mem[89619] = 16'b0000000000000000;
	sram_mem[89620] = 16'b0000000000000000;
	sram_mem[89621] = 16'b0000000000000000;
	sram_mem[89622] = 16'b0000000000000000;
	sram_mem[89623] = 16'b0000000000000000;
	sram_mem[89624] = 16'b0000000000000000;
	sram_mem[89625] = 16'b0000000000000000;
	sram_mem[89626] = 16'b0000000000000000;
	sram_mem[89627] = 16'b0000000000000000;
	sram_mem[89628] = 16'b0000000000000000;
	sram_mem[89629] = 16'b0000000000000000;
	sram_mem[89630] = 16'b0000000000000000;
	sram_mem[89631] = 16'b0000000000000000;
	sram_mem[89632] = 16'b0000000000000000;
	sram_mem[89633] = 16'b0000000000000000;
	sram_mem[89634] = 16'b0000000000000000;
	sram_mem[89635] = 16'b0000000000000000;
	sram_mem[89636] = 16'b0000000000000000;
	sram_mem[89637] = 16'b0000000000000000;
	sram_mem[89638] = 16'b0000000000000000;
	sram_mem[89639] = 16'b0000000000000000;
	sram_mem[89640] = 16'b0000000000000000;
	sram_mem[89641] = 16'b0000000000000000;
	sram_mem[89642] = 16'b0000000000000000;
	sram_mem[89643] = 16'b0000000000000000;
	sram_mem[89644] = 16'b0000000000000000;
	sram_mem[89645] = 16'b0000000000000000;
	sram_mem[89646] = 16'b0000000000000000;
	sram_mem[89647] = 16'b0000000000000000;
	sram_mem[89648] = 16'b0000000000000000;
	sram_mem[89649] = 16'b0000000000000000;
	sram_mem[89650] = 16'b0000000000000000;
	sram_mem[89651] = 16'b0000000000000000;
	sram_mem[89652] = 16'b0000000000000000;
	sram_mem[89653] = 16'b0000000000000000;
	sram_mem[89654] = 16'b0000000000000000;
	sram_mem[89655] = 16'b0000000000000000;
	sram_mem[89656] = 16'b0000000000000000;
	sram_mem[89657] = 16'b0000000000000000;
	sram_mem[89658] = 16'b0000000000000000;
	sram_mem[89659] = 16'b0000000000000000;
	sram_mem[89660] = 16'b0000000000000000;
	sram_mem[89661] = 16'b0000000000000000;
	sram_mem[89662] = 16'b0000000000000000;
	sram_mem[89663] = 16'b0000000000000000;
	sram_mem[89664] = 16'b0000000000000000;
	sram_mem[89665] = 16'b0000000000000000;
	sram_mem[89666] = 16'b0000000000000000;
	sram_mem[89667] = 16'b0000000000000000;
	sram_mem[89668] = 16'b0000000000000000;
	sram_mem[89669] = 16'b0000000000000000;
	sram_mem[89670] = 16'b0000000000000000;
	sram_mem[89671] = 16'b0000000000000000;
	sram_mem[89672] = 16'b0000000000000000;
	sram_mem[89673] = 16'b0000000000000000;
	sram_mem[89674] = 16'b0000000000000000;
	sram_mem[89675] = 16'b0000000000000000;
	sram_mem[89676] = 16'b0000000000000000;
	sram_mem[89677] = 16'b0000000000000000;
	sram_mem[89678] = 16'b0000000000000000;
	sram_mem[89679] = 16'b0000000000000000;
	sram_mem[89680] = 16'b0000000000000000;
	sram_mem[89681] = 16'b0000000000000000;
	sram_mem[89682] = 16'b0000000000000000;
	sram_mem[89683] = 16'b0000000000000000;
	sram_mem[89684] = 16'b0000000000000000;
	sram_mem[89685] = 16'b0000000000000000;
	sram_mem[89686] = 16'b0000000000000000;
	sram_mem[89687] = 16'b0000000000000000;
	sram_mem[89688] = 16'b0000000000000000;
	sram_mem[89689] = 16'b0000000000000000;
	sram_mem[89690] = 16'b0000000000000000;
	sram_mem[89691] = 16'b0000000000000000;
	sram_mem[89692] = 16'b0000000000000000;
	sram_mem[89693] = 16'b0000000000000000;
	sram_mem[89694] = 16'b0000000000000000;
	sram_mem[89695] = 16'b0000000000000000;
	sram_mem[89696] = 16'b0000000000000000;
	sram_mem[89697] = 16'b0000000000000000;
	sram_mem[89698] = 16'b0000000000000000;
	sram_mem[89699] = 16'b0000000000000000;
	sram_mem[89700] = 16'b0000000000000000;
	sram_mem[89701] = 16'b0000000000000000;
	sram_mem[89702] = 16'b0000000000000000;
	sram_mem[89703] = 16'b0000000000000000;
	sram_mem[89704] = 16'b0000000000000000;
	sram_mem[89705] = 16'b0000000000000000;
	sram_mem[89706] = 16'b0000000000000000;
	sram_mem[89707] = 16'b0000000000000000;
	sram_mem[89708] = 16'b0000000000000000;
	sram_mem[89709] = 16'b0000000000000000;
	sram_mem[89710] = 16'b0000000000000000;
	sram_mem[89711] = 16'b0000000000000000;
	sram_mem[89712] = 16'b0000000000000000;
	sram_mem[89713] = 16'b0000000000000000;
	sram_mem[89714] = 16'b0000000000000000;
	sram_mem[89715] = 16'b0000000000000000;
	sram_mem[89716] = 16'b0000000000000000;
	sram_mem[89717] = 16'b0000000000000000;
	sram_mem[89718] = 16'b0000000000000000;
	sram_mem[89719] = 16'b0000000000000000;
	sram_mem[89720] = 16'b0000000000000000;
	sram_mem[89721] = 16'b0000000000000000;
	sram_mem[89722] = 16'b0000000000000000;
	sram_mem[89723] = 16'b0000000000000000;
	sram_mem[89724] = 16'b0000000000000000;
	sram_mem[89725] = 16'b0000000000000000;
	sram_mem[89726] = 16'b0000000000000000;
	sram_mem[89727] = 16'b0000000000000000;
	sram_mem[89728] = 16'b0000000000000000;
	sram_mem[89729] = 16'b0000000000000000;
	sram_mem[89730] = 16'b0000000000000000;
	sram_mem[89731] = 16'b0000000000000000;
	sram_mem[89732] = 16'b0000000000000000;
	sram_mem[89733] = 16'b0000000000000000;
	sram_mem[89734] = 16'b0000000000000000;
	sram_mem[89735] = 16'b0000000000000000;
	sram_mem[89736] = 16'b0000000000000000;
	sram_mem[89737] = 16'b0000000000000000;
	sram_mem[89738] = 16'b0000000000000000;
	sram_mem[89739] = 16'b0000000000000000;
	sram_mem[89740] = 16'b0000000000000000;
	sram_mem[89741] = 16'b0000000000000000;
	sram_mem[89742] = 16'b0000000000000000;
	sram_mem[89743] = 16'b0000000000000000;
	sram_mem[89744] = 16'b0000000000000000;
	sram_mem[89745] = 16'b0000000000000000;
	sram_mem[89746] = 16'b0000000000000000;
	sram_mem[89747] = 16'b0000000000000000;
	sram_mem[89748] = 16'b0000000000000000;
	sram_mem[89749] = 16'b0000000000000000;
	sram_mem[89750] = 16'b0000000000000000;
	sram_mem[89751] = 16'b0000000000000000;
	sram_mem[89752] = 16'b0000000000000000;
	sram_mem[89753] = 16'b0000000000000000;
	sram_mem[89754] = 16'b0000000000000000;
	sram_mem[89755] = 16'b0000000000000000;
	sram_mem[89756] = 16'b0000000000000000;
	sram_mem[89757] = 16'b0000000000000000;
	sram_mem[89758] = 16'b0000000000000000;
	sram_mem[89759] = 16'b0000000000000000;
	sram_mem[89760] = 16'b0000000000000000;
	sram_mem[89761] = 16'b0000000000000000;
	sram_mem[89762] = 16'b0000000000000000;
	sram_mem[89763] = 16'b0000000000000000;
	sram_mem[89764] = 16'b0000000000000000;
	sram_mem[89765] = 16'b0000000000000000;
	sram_mem[89766] = 16'b0000000000000000;
	sram_mem[89767] = 16'b0000000000000000;
	sram_mem[89768] = 16'b0000000000000000;
	sram_mem[89769] = 16'b0000000000000000;
	sram_mem[89770] = 16'b0000000000000000;
	sram_mem[89771] = 16'b0000000000000000;
	sram_mem[89772] = 16'b0000000000000000;
	sram_mem[89773] = 16'b0000000000000000;
	sram_mem[89774] = 16'b0000000000000000;
	sram_mem[89775] = 16'b0000000000000000;
	sram_mem[89776] = 16'b0000000000000000;
	sram_mem[89777] = 16'b0000000000000000;
	sram_mem[89778] = 16'b0000000000000000;
	sram_mem[89779] = 16'b0000000000000000;
	sram_mem[89780] = 16'b0000000000000000;
	sram_mem[89781] = 16'b0000000000000000;
	sram_mem[89782] = 16'b0000000000000000;
	sram_mem[89783] = 16'b0000000000000000;
	sram_mem[89784] = 16'b0000000000000000;
	sram_mem[89785] = 16'b0000000000000000;
	sram_mem[89786] = 16'b0000000000000000;
	sram_mem[89787] = 16'b0000000000000000;
	sram_mem[89788] = 16'b0000000000000000;
	sram_mem[89789] = 16'b0000000000000000;
	sram_mem[89790] = 16'b0000000000000000;
	sram_mem[89791] = 16'b0000000000000000;
	sram_mem[89792] = 16'b0000000000000000;
	sram_mem[89793] = 16'b0000000000000000;
	sram_mem[89794] = 16'b0000000000000000;
	sram_mem[89795] = 16'b0000000000000000;
	sram_mem[89796] = 16'b0000000000000000;
	sram_mem[89797] = 16'b0000000000000000;
	sram_mem[89798] = 16'b0000000000000000;
	sram_mem[89799] = 16'b0000000000000000;
	sram_mem[89800] = 16'b0000000000000000;
	sram_mem[89801] = 16'b0000000000000000;
	sram_mem[89802] = 16'b0000000000000000;
	sram_mem[89803] = 16'b0000000000000000;
	sram_mem[89804] = 16'b0000000000000000;
	sram_mem[89805] = 16'b0000000000000000;
	sram_mem[89806] = 16'b0000000000000000;
	sram_mem[89807] = 16'b0000000000000000;
	sram_mem[89808] = 16'b0000000000000000;
	sram_mem[89809] = 16'b0000000000000000;
	sram_mem[89810] = 16'b0000000000000000;
	sram_mem[89811] = 16'b0000000000000000;
	sram_mem[89812] = 16'b0000000000000000;
	sram_mem[89813] = 16'b0000000000000000;
	sram_mem[89814] = 16'b0000000000000000;
	sram_mem[89815] = 16'b0000000000000000;
	sram_mem[89816] = 16'b0000000000000000;
	sram_mem[89817] = 16'b0000000000000000;
	sram_mem[89818] = 16'b0000000000000000;
	sram_mem[89819] = 16'b0000000000000000;
	sram_mem[89820] = 16'b0000000000000000;
	sram_mem[89821] = 16'b0000000000000000;
	sram_mem[89822] = 16'b0000000000000000;
	sram_mem[89823] = 16'b0000000000000000;
	sram_mem[89824] = 16'b0000000000000000;
	sram_mem[89825] = 16'b0000000000000000;
	sram_mem[89826] = 16'b0000000000000000;
	sram_mem[89827] = 16'b0000000000000000;
	sram_mem[89828] = 16'b0000000000000000;
	sram_mem[89829] = 16'b0000000000000000;
	sram_mem[89830] = 16'b0000000000000000;
	sram_mem[89831] = 16'b0000000000000000;
	sram_mem[89832] = 16'b0000000000000000;
	sram_mem[89833] = 16'b0000000000000000;
	sram_mem[89834] = 16'b0000000000000000;
	sram_mem[89835] = 16'b0000000000000000;
	sram_mem[89836] = 16'b0000000000000000;
	sram_mem[89837] = 16'b0000000000000000;
	sram_mem[89838] = 16'b0000000000000000;
	sram_mem[89839] = 16'b0000000000000000;
	sram_mem[89840] = 16'b0000000000000000;
	sram_mem[89841] = 16'b0000000000000000;
	sram_mem[89842] = 16'b0000000000000000;
	sram_mem[89843] = 16'b0000000000000000;
	sram_mem[89844] = 16'b0000000000000000;
	sram_mem[89845] = 16'b0000000000000000;
	sram_mem[89846] = 16'b0000000000000000;
	sram_mem[89847] = 16'b0000000000000000;
	sram_mem[89848] = 16'b0000000000000000;
	sram_mem[89849] = 16'b0000000000000000;
	sram_mem[89850] = 16'b0000000000000000;
	sram_mem[89851] = 16'b0000000000000000;
	sram_mem[89852] = 16'b0000000000000000;
	sram_mem[89853] = 16'b0000000000000000;
	sram_mem[89854] = 16'b0000000000000000;
	sram_mem[89855] = 16'b0000000000000000;
	sram_mem[89856] = 16'b0000000000000000;
	sram_mem[89857] = 16'b0000000000000000;
	sram_mem[89858] = 16'b0000000000000000;
	sram_mem[89859] = 16'b0000000000000000;
	sram_mem[89860] = 16'b0000000000000000;
	sram_mem[89861] = 16'b0000000000000000;
	sram_mem[89862] = 16'b0000000000000000;
	sram_mem[89863] = 16'b0000000000000000;
	sram_mem[89864] = 16'b0000000000000000;
	sram_mem[89865] = 16'b0000000000000000;
	sram_mem[89866] = 16'b0000000000000000;
	sram_mem[89867] = 16'b0000000000000000;
	sram_mem[89868] = 16'b0000000000000000;
	sram_mem[89869] = 16'b0000000000000000;
	sram_mem[89870] = 16'b0000000000000000;
	sram_mem[89871] = 16'b0000000000000000;
	sram_mem[89872] = 16'b0000000000000000;
	sram_mem[89873] = 16'b0000000000000000;
	sram_mem[89874] = 16'b0000000000000000;
	sram_mem[89875] = 16'b0000000000000000;
	sram_mem[89876] = 16'b0000000000000000;
	sram_mem[89877] = 16'b0000000000000000;
	sram_mem[89878] = 16'b0000000000000000;
	sram_mem[89879] = 16'b0000000000000000;
	sram_mem[89880] = 16'b0000000000000000;
	sram_mem[89881] = 16'b0000000000000000;
	sram_mem[89882] = 16'b0000000000000000;
	sram_mem[89883] = 16'b0000000000000000;
	sram_mem[89884] = 16'b0000000000000000;
	sram_mem[89885] = 16'b0000000000000000;
	sram_mem[89886] = 16'b0000000000000000;
	sram_mem[89887] = 16'b0000000000000000;
	sram_mem[89888] = 16'b0000000000000000;
	sram_mem[89889] = 16'b0000000000000000;
	sram_mem[89890] = 16'b0000000000000000;
	sram_mem[89891] = 16'b0000000000000000;
	sram_mem[89892] = 16'b0000000000000000;
	sram_mem[89893] = 16'b0000000000000000;
	sram_mem[89894] = 16'b0000000000000000;
	sram_mem[89895] = 16'b0000000000000000;
	sram_mem[89896] = 16'b0000000000000000;
	sram_mem[89897] = 16'b0000000000000000;
	sram_mem[89898] = 16'b0000000000000000;
	sram_mem[89899] = 16'b0000000000000000;
	sram_mem[89900] = 16'b0000000000000000;
	sram_mem[89901] = 16'b0000000000000000;
	sram_mem[89902] = 16'b0000000000000000;
	sram_mem[89903] = 16'b0000000000000000;
	sram_mem[89904] = 16'b0000000000000000;
	sram_mem[89905] = 16'b0000000000000000;
	sram_mem[89906] = 16'b0000000000000000;
	sram_mem[89907] = 16'b0000000000000000;
	sram_mem[89908] = 16'b0000000000000000;
	sram_mem[89909] = 16'b0000000000000000;
	sram_mem[89910] = 16'b0000000000000000;
	sram_mem[89911] = 16'b0000000000000000;
	sram_mem[89912] = 16'b0000000000000000;
	sram_mem[89913] = 16'b0000000000000000;
	sram_mem[89914] = 16'b0000000000000000;
	sram_mem[89915] = 16'b0000000000000000;
	sram_mem[89916] = 16'b0000000000000000;
	sram_mem[89917] = 16'b0000000000000000;
	sram_mem[89918] = 16'b0000000000000000;
	sram_mem[89919] = 16'b0000000000000000;
	sram_mem[89920] = 16'b0000000000000000;
	sram_mem[89921] = 16'b0000000000000000;
	sram_mem[89922] = 16'b0000000000000000;
	sram_mem[89923] = 16'b0000000000000000;
	sram_mem[89924] = 16'b0000000000000000;
	sram_mem[89925] = 16'b0000000000000000;
	sram_mem[89926] = 16'b0000000000000000;
	sram_mem[89927] = 16'b0000000000000000;
	sram_mem[89928] = 16'b0000000000000000;
	sram_mem[89929] = 16'b0000000000000000;
	sram_mem[89930] = 16'b0000000000000000;
	sram_mem[89931] = 16'b0000000000000000;
	sram_mem[89932] = 16'b0000000000000000;
	sram_mem[89933] = 16'b0000000000000000;
	sram_mem[89934] = 16'b0000000000000000;
	sram_mem[89935] = 16'b0000000000000000;
	sram_mem[89936] = 16'b0000000000000000;
	sram_mem[89937] = 16'b0000000000000000;
	sram_mem[89938] = 16'b0000000000000000;
	sram_mem[89939] = 16'b0000000000000000;
	sram_mem[89940] = 16'b0000000000000000;
	sram_mem[89941] = 16'b0000000000000000;
	sram_mem[89942] = 16'b0000000000000000;
	sram_mem[89943] = 16'b0000000000000000;
	sram_mem[89944] = 16'b0000000000000000;
	sram_mem[89945] = 16'b0000000000000000;
	sram_mem[89946] = 16'b0000000000000000;
	sram_mem[89947] = 16'b0000000000000000;
	sram_mem[89948] = 16'b0000000000000000;
	sram_mem[89949] = 16'b0000000000000000;
	sram_mem[89950] = 16'b0000000000000000;
	sram_mem[89951] = 16'b0000000000000000;
	sram_mem[89952] = 16'b0000000000000000;
	sram_mem[89953] = 16'b0000000000000000;
	sram_mem[89954] = 16'b0000000000000000;
	sram_mem[89955] = 16'b0000000000000000;
	sram_mem[89956] = 16'b0000000000000000;
	sram_mem[89957] = 16'b0000000000000000;
	sram_mem[89958] = 16'b0000000000000000;
	sram_mem[89959] = 16'b0000000000000000;
	sram_mem[89960] = 16'b0000000000000000;
	sram_mem[89961] = 16'b0000000000000000;
	sram_mem[89962] = 16'b0000000000000000;
	sram_mem[89963] = 16'b0000000000000000;
	sram_mem[89964] = 16'b0000000000000000;
	sram_mem[89965] = 16'b0000000000000000;
	sram_mem[89966] = 16'b0000000000000000;
	sram_mem[89967] = 16'b0000000000000000;
	sram_mem[89968] = 16'b0000000000000000;
	sram_mem[89969] = 16'b0000000000000000;
	sram_mem[89970] = 16'b0000000000000000;
	sram_mem[89971] = 16'b0000000000000000;
	sram_mem[89972] = 16'b0000000000000000;
	sram_mem[89973] = 16'b0000000000000000;
	sram_mem[89974] = 16'b0000000000000000;
	sram_mem[89975] = 16'b0000000000000000;
	sram_mem[89976] = 16'b0000000000000000;
	sram_mem[89977] = 16'b0000000000000000;
	sram_mem[89978] = 16'b0000000000000000;
	sram_mem[89979] = 16'b0000000000000000;
	sram_mem[89980] = 16'b0000000000000000;
	sram_mem[89981] = 16'b0000000000000000;
	sram_mem[89982] = 16'b0000000000000000;
	sram_mem[89983] = 16'b0000000000000000;
	sram_mem[89984] = 16'b0000000000000000;
	sram_mem[89985] = 16'b0000000000000000;
	sram_mem[89986] = 16'b0000000000000000;
	sram_mem[89987] = 16'b0000000000000000;
	sram_mem[89988] = 16'b0000000000000000;
	sram_mem[89989] = 16'b0000000000000000;
	sram_mem[89990] = 16'b0000000000000000;
	sram_mem[89991] = 16'b0000000000000000;
	sram_mem[89992] = 16'b0000000000000000;
	sram_mem[89993] = 16'b0000000000000000;
	sram_mem[89994] = 16'b0000000000000000;
	sram_mem[89995] = 16'b0000000000000000;
	sram_mem[89996] = 16'b0000000000000000;
	sram_mem[89997] = 16'b0000000000000000;
	sram_mem[89998] = 16'b0000000000000000;
	sram_mem[89999] = 16'b0000000000000000;
	sram_mem[90000] = 16'b0000000000000000;
	sram_mem[90001] = 16'b0000000000000000;
	sram_mem[90002] = 16'b0000000000000000;
	sram_mem[90003] = 16'b0000000000000000;
	sram_mem[90004] = 16'b0000000000000000;
	sram_mem[90005] = 16'b0000000000000000;
	sram_mem[90006] = 16'b0000000000000000;
	sram_mem[90007] = 16'b0000000000000000;
	sram_mem[90008] = 16'b0000000000000000;
	sram_mem[90009] = 16'b0000000000000000;
	sram_mem[90010] = 16'b0000000000000000;
	sram_mem[90011] = 16'b0000000000000000;
	sram_mem[90012] = 16'b0000000000000000;
	sram_mem[90013] = 16'b0000000000000000;
	sram_mem[90014] = 16'b0000000000000000;
	sram_mem[90015] = 16'b0000000000000000;
	sram_mem[90016] = 16'b0000000000000000;
	sram_mem[90017] = 16'b0000000000000000;
	sram_mem[90018] = 16'b0000000000000000;
	sram_mem[90019] = 16'b0000000000000000;
	sram_mem[90020] = 16'b0000000000000000;
	sram_mem[90021] = 16'b0000000000000000;
	sram_mem[90022] = 16'b0000000000000000;
	sram_mem[90023] = 16'b0000000000000000;
	sram_mem[90024] = 16'b0000000000000000;
	sram_mem[90025] = 16'b0000000000000000;
	sram_mem[90026] = 16'b0000000000000000;
	sram_mem[90027] = 16'b0000000000000000;
	sram_mem[90028] = 16'b0000000000000000;
	sram_mem[90029] = 16'b0000000000000000;
	sram_mem[90030] = 16'b0000000000000000;
	sram_mem[90031] = 16'b0000000000000000;
	sram_mem[90032] = 16'b0000000000000000;
	sram_mem[90033] = 16'b0000000000000000;
	sram_mem[90034] = 16'b0000000000000000;
	sram_mem[90035] = 16'b0000000000000000;
	sram_mem[90036] = 16'b0000000000000000;
	sram_mem[90037] = 16'b0000000000000000;
	sram_mem[90038] = 16'b0000000000000000;
	sram_mem[90039] = 16'b0000000000000000;
	sram_mem[90040] = 16'b0000000000000000;
	sram_mem[90041] = 16'b0000000000000000;
	sram_mem[90042] = 16'b0000000000000000;
	sram_mem[90043] = 16'b0000000000000000;
	sram_mem[90044] = 16'b0000000000000000;
	sram_mem[90045] = 16'b0000000000000000;
	sram_mem[90046] = 16'b0000000000000000;
	sram_mem[90047] = 16'b0000000000000000;
	sram_mem[90048] = 16'b0000000000000000;
	sram_mem[90049] = 16'b0000000000000000;
	sram_mem[90050] = 16'b0000000000000000;
	sram_mem[90051] = 16'b0000000000000000;
	sram_mem[90052] = 16'b0000000000000000;
	sram_mem[90053] = 16'b0000000000000000;
	sram_mem[90054] = 16'b0000000000000000;
	sram_mem[90055] = 16'b0000000000000000;
	sram_mem[90056] = 16'b0000000000000000;
	sram_mem[90057] = 16'b0000000000000000;
	sram_mem[90058] = 16'b0000000000000000;
	sram_mem[90059] = 16'b0000000000000000;
	sram_mem[90060] = 16'b0000000000000000;
	sram_mem[90061] = 16'b0000000000000000;
	sram_mem[90062] = 16'b0000000000000000;
	sram_mem[90063] = 16'b0000000000000000;
	sram_mem[90064] = 16'b0000000000000000;
	sram_mem[90065] = 16'b0000000000000000;
	sram_mem[90066] = 16'b0000000000000000;
	sram_mem[90067] = 16'b0000000000000000;
	sram_mem[90068] = 16'b0000000000000000;
	sram_mem[90069] = 16'b0000000000000000;
	sram_mem[90070] = 16'b0000000000000000;
	sram_mem[90071] = 16'b0000000000000000;
	sram_mem[90072] = 16'b0000000000000000;
	sram_mem[90073] = 16'b0000000000000000;
	sram_mem[90074] = 16'b0000000000000000;
	sram_mem[90075] = 16'b0000000000000000;
	sram_mem[90076] = 16'b0000000000000000;
	sram_mem[90077] = 16'b0000000000000000;
	sram_mem[90078] = 16'b0000000000000000;
	sram_mem[90079] = 16'b0000000000000000;
	sram_mem[90080] = 16'b0000000000000000;
	sram_mem[90081] = 16'b0000000000000000;
	sram_mem[90082] = 16'b0000000000000000;
	sram_mem[90083] = 16'b0000000000000000;
	sram_mem[90084] = 16'b0000000000000000;
	sram_mem[90085] = 16'b0000000000000000;
	sram_mem[90086] = 16'b0000000000000000;
	sram_mem[90087] = 16'b0000000000000000;
	sram_mem[90088] = 16'b0000000000000000;
	sram_mem[90089] = 16'b0000000000000000;
	sram_mem[90090] = 16'b0000000000000000;
	sram_mem[90091] = 16'b0000000000000000;
	sram_mem[90092] = 16'b0000000000000000;
	sram_mem[90093] = 16'b0000000000000000;
	sram_mem[90094] = 16'b0000000000000000;
	sram_mem[90095] = 16'b0000000000000000;
	sram_mem[90096] = 16'b0000000000000000;
	sram_mem[90097] = 16'b0000000000000000;
	sram_mem[90098] = 16'b0000000000000000;
	sram_mem[90099] = 16'b0000000000000000;
	sram_mem[90100] = 16'b0000000000000000;
	sram_mem[90101] = 16'b0000000000000000;
	sram_mem[90102] = 16'b0000000000000000;
	sram_mem[90103] = 16'b0000000000000000;
	sram_mem[90104] = 16'b0000000000000000;
	sram_mem[90105] = 16'b0000000000000000;
	sram_mem[90106] = 16'b0000000000000000;
	sram_mem[90107] = 16'b0000000000000000;
	sram_mem[90108] = 16'b0000000000000000;
	sram_mem[90109] = 16'b0000000000000000;
	sram_mem[90110] = 16'b0000000000000000;
	sram_mem[90111] = 16'b0000000000000000;
	sram_mem[90112] = 16'b0000000000000000;
	sram_mem[90113] = 16'b0000000000000000;
	sram_mem[90114] = 16'b0000000000000000;
	sram_mem[90115] = 16'b0000000000000000;
	sram_mem[90116] = 16'b0000000000000000;
	sram_mem[90117] = 16'b0000000000000000;
	sram_mem[90118] = 16'b0000000000000000;
	sram_mem[90119] = 16'b0000000000000000;
	sram_mem[90120] = 16'b0000000000000000;
	sram_mem[90121] = 16'b0000000000000000;
	sram_mem[90122] = 16'b0000000000000000;
	sram_mem[90123] = 16'b0000000000000000;
	sram_mem[90124] = 16'b0000000000000000;
	sram_mem[90125] = 16'b0000000000000000;
	sram_mem[90126] = 16'b0000000000000000;
	sram_mem[90127] = 16'b0000000000000000;
	sram_mem[90128] = 16'b0000000000000000;
	sram_mem[90129] = 16'b0000000000000000;
	sram_mem[90130] = 16'b0000000000000000;
	sram_mem[90131] = 16'b0000000000000000;
	sram_mem[90132] = 16'b0000000000000000;
	sram_mem[90133] = 16'b0000000000000000;
	sram_mem[90134] = 16'b0000000000000000;
	sram_mem[90135] = 16'b0000000000000000;
	sram_mem[90136] = 16'b0000000000000000;
	sram_mem[90137] = 16'b0000000000000000;
	sram_mem[90138] = 16'b0000000000000000;
	sram_mem[90139] = 16'b0000000000000000;
	sram_mem[90140] = 16'b0000000000000000;
	sram_mem[90141] = 16'b0000000000000000;
	sram_mem[90142] = 16'b0000000000000000;
	sram_mem[90143] = 16'b0000000000000000;
	sram_mem[90144] = 16'b0000000000000000;
	sram_mem[90145] = 16'b0000000000000000;
	sram_mem[90146] = 16'b0000000000000000;
	sram_mem[90147] = 16'b0000000000000000;
	sram_mem[90148] = 16'b0000000000000000;
	sram_mem[90149] = 16'b0000000000000000;
	sram_mem[90150] = 16'b0000000000000000;
	sram_mem[90151] = 16'b0000000000000000;
	sram_mem[90152] = 16'b0000000000000000;
	sram_mem[90153] = 16'b0000000000000000;
	sram_mem[90154] = 16'b0000000000000000;
	sram_mem[90155] = 16'b0000000000000000;
	sram_mem[90156] = 16'b0000000000000000;
	sram_mem[90157] = 16'b0000000000000000;
	sram_mem[90158] = 16'b0000000000000000;
	sram_mem[90159] = 16'b0000000000000000;
	sram_mem[90160] = 16'b0000000000000000;
	sram_mem[90161] = 16'b0000000000000000;
	sram_mem[90162] = 16'b0000000000000000;
	sram_mem[90163] = 16'b0000000000000000;
	sram_mem[90164] = 16'b0000000000000000;
	sram_mem[90165] = 16'b0000000000000000;
	sram_mem[90166] = 16'b0000000000000000;
	sram_mem[90167] = 16'b0000000000000000;
	sram_mem[90168] = 16'b0000000000000000;
	sram_mem[90169] = 16'b0000000000000000;
	sram_mem[90170] = 16'b0000000000000000;
	sram_mem[90171] = 16'b0000000000000000;
	sram_mem[90172] = 16'b0000000000000000;
	sram_mem[90173] = 16'b0000000000000000;
	sram_mem[90174] = 16'b0000000000000000;
	sram_mem[90175] = 16'b0000000000000000;
	sram_mem[90176] = 16'b0000000000000000;
	sram_mem[90177] = 16'b0000000000000000;
	sram_mem[90178] = 16'b0000000000000000;
	sram_mem[90179] = 16'b0000000000000000;
	sram_mem[90180] = 16'b0000000000000000;
	sram_mem[90181] = 16'b0000000000000000;
	sram_mem[90182] = 16'b0000000000000000;
	sram_mem[90183] = 16'b0000000000000000;
	sram_mem[90184] = 16'b0000000000000000;
	sram_mem[90185] = 16'b0000000000000000;
	sram_mem[90186] = 16'b0000000000000000;
	sram_mem[90187] = 16'b0000000000000000;
	sram_mem[90188] = 16'b0000000000000000;
	sram_mem[90189] = 16'b0000000000000000;
	sram_mem[90190] = 16'b0000000000000000;
	sram_mem[90191] = 16'b0000000000000000;
	sram_mem[90192] = 16'b0000000000000000;
	sram_mem[90193] = 16'b0000000000000000;
	sram_mem[90194] = 16'b0000000000000000;
	sram_mem[90195] = 16'b0000000000000000;
	sram_mem[90196] = 16'b0000000000000000;
	sram_mem[90197] = 16'b0000000000000000;
	sram_mem[90198] = 16'b0000000000000000;
	sram_mem[90199] = 16'b0000000000000000;
	sram_mem[90200] = 16'b0000000000000000;
	sram_mem[90201] = 16'b0000000000000000;
	sram_mem[90202] = 16'b0000000000000000;
	sram_mem[90203] = 16'b0000000000000000;
	sram_mem[90204] = 16'b0000000000000000;
	sram_mem[90205] = 16'b0000000000000000;
	sram_mem[90206] = 16'b0000000000000000;
	sram_mem[90207] = 16'b0000000000000000;
	sram_mem[90208] = 16'b0000000000000000;
	sram_mem[90209] = 16'b0000000000000000;
	sram_mem[90210] = 16'b0000000000000000;
	sram_mem[90211] = 16'b0000000000000000;
	sram_mem[90212] = 16'b0000000000000000;
	sram_mem[90213] = 16'b0000000000000000;
	sram_mem[90214] = 16'b0000000000000000;
	sram_mem[90215] = 16'b0000000000000000;
	sram_mem[90216] = 16'b0000000000000000;
	sram_mem[90217] = 16'b0000000000000000;
	sram_mem[90218] = 16'b0000000000000000;
	sram_mem[90219] = 16'b0000000000000000;
	sram_mem[90220] = 16'b0000000000000000;
	sram_mem[90221] = 16'b0000000000000000;
	sram_mem[90222] = 16'b0000000000000000;
	sram_mem[90223] = 16'b0000000000000000;
	sram_mem[90224] = 16'b0000000000000000;
	sram_mem[90225] = 16'b0000000000000000;
	sram_mem[90226] = 16'b0000000000000000;
	sram_mem[90227] = 16'b0000000000000000;
	sram_mem[90228] = 16'b0000000000000000;
	sram_mem[90229] = 16'b0000000000000000;
	sram_mem[90230] = 16'b0000000000000000;
	sram_mem[90231] = 16'b0000000000000000;
	sram_mem[90232] = 16'b0000000000000000;
	sram_mem[90233] = 16'b0000000000000000;
	sram_mem[90234] = 16'b0000000000000000;
	sram_mem[90235] = 16'b0000000000000000;
	sram_mem[90236] = 16'b0000000000000000;
	sram_mem[90237] = 16'b0000000000000000;
	sram_mem[90238] = 16'b0000000000000000;
	sram_mem[90239] = 16'b0000000000000000;
	sram_mem[90240] = 16'b0000000000000000;
	sram_mem[90241] = 16'b0000000000000000;
	sram_mem[90242] = 16'b0000000000000000;
	sram_mem[90243] = 16'b0000000000000000;
	sram_mem[90244] = 16'b0000000000000000;
	sram_mem[90245] = 16'b0000000000000000;
	sram_mem[90246] = 16'b0000000000000000;
	sram_mem[90247] = 16'b0000000000000000;
	sram_mem[90248] = 16'b0000000000000000;
	sram_mem[90249] = 16'b0000000000000000;
	sram_mem[90250] = 16'b0000000000000000;
	sram_mem[90251] = 16'b0000000000000000;
	sram_mem[90252] = 16'b0000000000000000;
	sram_mem[90253] = 16'b0000000000000000;
	sram_mem[90254] = 16'b0000000000000000;
	sram_mem[90255] = 16'b0000000000000000;
	sram_mem[90256] = 16'b0000000000000000;
	sram_mem[90257] = 16'b0000000000000000;
	sram_mem[90258] = 16'b0000000000000000;
	sram_mem[90259] = 16'b0000000000000000;
	sram_mem[90260] = 16'b0000000000000000;
	sram_mem[90261] = 16'b0000000000000000;
	sram_mem[90262] = 16'b0000000000000000;
	sram_mem[90263] = 16'b0000000000000000;
	sram_mem[90264] = 16'b0000000000000000;
	sram_mem[90265] = 16'b0000000000000000;
	sram_mem[90266] = 16'b0000000000000000;
	sram_mem[90267] = 16'b0000000000000000;
	sram_mem[90268] = 16'b0000000000000000;
	sram_mem[90269] = 16'b0000000000000000;
	sram_mem[90270] = 16'b0000000000000000;
	sram_mem[90271] = 16'b0000000000000000;
	sram_mem[90272] = 16'b0000000000000000;
	sram_mem[90273] = 16'b0000000000000000;
	sram_mem[90274] = 16'b0000000000000000;
	sram_mem[90275] = 16'b0000000000000000;
	sram_mem[90276] = 16'b0000000000000000;
	sram_mem[90277] = 16'b0000000000000000;
	sram_mem[90278] = 16'b0000000000000000;
	sram_mem[90279] = 16'b0000000000000000;
	sram_mem[90280] = 16'b0000000000000000;
	sram_mem[90281] = 16'b0000000000000000;
	sram_mem[90282] = 16'b0000000000000000;
	sram_mem[90283] = 16'b0000000000000000;
	sram_mem[90284] = 16'b0000000000000000;
	sram_mem[90285] = 16'b0000000000000000;
	sram_mem[90286] = 16'b0000000000000000;
	sram_mem[90287] = 16'b0000000000000000;
	sram_mem[90288] = 16'b0000000000000000;
	sram_mem[90289] = 16'b0000000000000000;
	sram_mem[90290] = 16'b0000000000000000;
	sram_mem[90291] = 16'b0000000000000000;
	sram_mem[90292] = 16'b0000000000000000;
	sram_mem[90293] = 16'b0000000000000000;
	sram_mem[90294] = 16'b0000000000000000;
	sram_mem[90295] = 16'b0000000000000000;
	sram_mem[90296] = 16'b0000000000000000;
	sram_mem[90297] = 16'b0000000000000000;
	sram_mem[90298] = 16'b0000000000000000;
	sram_mem[90299] = 16'b0000000000000000;
	sram_mem[90300] = 16'b0000000000000000;
	sram_mem[90301] = 16'b0000000000000000;
	sram_mem[90302] = 16'b0000000000000000;
	sram_mem[90303] = 16'b0000000000000000;
	sram_mem[90304] = 16'b0000000000000000;
	sram_mem[90305] = 16'b0000000000000000;
	sram_mem[90306] = 16'b0000000000000000;
	sram_mem[90307] = 16'b0000000000000000;
	sram_mem[90308] = 16'b0000000000000000;
	sram_mem[90309] = 16'b0000000000000000;
	sram_mem[90310] = 16'b0000000000000000;
	sram_mem[90311] = 16'b0000000000000000;
	sram_mem[90312] = 16'b0000000000000000;
	sram_mem[90313] = 16'b0000000000000000;
	sram_mem[90314] = 16'b0000000000000000;
	sram_mem[90315] = 16'b0000000000000000;
	sram_mem[90316] = 16'b0000000000000000;
	sram_mem[90317] = 16'b0000000000000000;
	sram_mem[90318] = 16'b0000000000000000;
	sram_mem[90319] = 16'b0000000000000000;
	sram_mem[90320] = 16'b0000000000000000;
	sram_mem[90321] = 16'b0000000000000000;
	sram_mem[90322] = 16'b0000000000000000;
	sram_mem[90323] = 16'b0000000000000000;
	sram_mem[90324] = 16'b0000000000000000;
	sram_mem[90325] = 16'b0000000000000000;
	sram_mem[90326] = 16'b0000000000000000;
	sram_mem[90327] = 16'b0000000000000000;
	sram_mem[90328] = 16'b0000000000000000;
	sram_mem[90329] = 16'b0000000000000000;
	sram_mem[90330] = 16'b0000000000000000;
	sram_mem[90331] = 16'b0000000000000000;
	sram_mem[90332] = 16'b0000000000000000;
	sram_mem[90333] = 16'b0000000000000000;
	sram_mem[90334] = 16'b0000000000000000;
	sram_mem[90335] = 16'b0000000000000000;
	sram_mem[90336] = 16'b0000000000000000;
	sram_mem[90337] = 16'b0000000000000000;
	sram_mem[90338] = 16'b0000000000000000;
	sram_mem[90339] = 16'b0000000000000000;
	sram_mem[90340] = 16'b0000000000000000;
	sram_mem[90341] = 16'b0000000000000000;
	sram_mem[90342] = 16'b0000000000000000;
	sram_mem[90343] = 16'b0000000000000000;
	sram_mem[90344] = 16'b0000000000000000;
	sram_mem[90345] = 16'b0000000000000000;
	sram_mem[90346] = 16'b0000000000000000;
	sram_mem[90347] = 16'b0000000000000000;
	sram_mem[90348] = 16'b0000000000000000;
	sram_mem[90349] = 16'b0000000000000000;
	sram_mem[90350] = 16'b0000000000000000;
	sram_mem[90351] = 16'b0000000000000000;
	sram_mem[90352] = 16'b0000000000000000;
	sram_mem[90353] = 16'b0000000000000000;
	sram_mem[90354] = 16'b0000000000000000;
	sram_mem[90355] = 16'b0000000000000000;
	sram_mem[90356] = 16'b0000000000000000;
	sram_mem[90357] = 16'b0000000000000000;
	sram_mem[90358] = 16'b0000000000000000;
	sram_mem[90359] = 16'b0000000000000000;
	sram_mem[90360] = 16'b0000000000000000;
	sram_mem[90361] = 16'b0000000000000000;
	sram_mem[90362] = 16'b0000000000000000;
	sram_mem[90363] = 16'b0000000000000000;
	sram_mem[90364] = 16'b0000000000000000;
	sram_mem[90365] = 16'b0000000000000000;
	sram_mem[90366] = 16'b0000000000000000;
	sram_mem[90367] = 16'b0000000000000000;
	sram_mem[90368] = 16'b0000000000000000;
	sram_mem[90369] = 16'b0000000000000000;
	sram_mem[90370] = 16'b0000000000000000;
	sram_mem[90371] = 16'b0000000000000000;
	sram_mem[90372] = 16'b0000000000000000;
	sram_mem[90373] = 16'b0000000000000000;
	sram_mem[90374] = 16'b0000000000000000;
	sram_mem[90375] = 16'b0000000000000000;
	sram_mem[90376] = 16'b0000000000000000;
	sram_mem[90377] = 16'b0000000000000000;
	sram_mem[90378] = 16'b0000000000000000;
	sram_mem[90379] = 16'b0000000000000000;
	sram_mem[90380] = 16'b0000000000000000;
	sram_mem[90381] = 16'b0000000000000000;
	sram_mem[90382] = 16'b0000000000000000;
	sram_mem[90383] = 16'b0000000000000000;
	sram_mem[90384] = 16'b0000000000000000;
	sram_mem[90385] = 16'b0000000000000000;
	sram_mem[90386] = 16'b0000000000000000;
	sram_mem[90387] = 16'b0000000000000000;
	sram_mem[90388] = 16'b0000000000000000;
	sram_mem[90389] = 16'b0000000000000000;
	sram_mem[90390] = 16'b0000000000000000;
	sram_mem[90391] = 16'b0000000000000000;
	sram_mem[90392] = 16'b0000000000000000;
	sram_mem[90393] = 16'b0000000000000000;
	sram_mem[90394] = 16'b0000000000000000;
	sram_mem[90395] = 16'b0000000000000000;
	sram_mem[90396] = 16'b0000000000000000;
	sram_mem[90397] = 16'b0000000000000000;
	sram_mem[90398] = 16'b0000000000000000;
	sram_mem[90399] = 16'b0000000000000000;
	sram_mem[90400] = 16'b0000000000000000;
	sram_mem[90401] = 16'b0000000000000000;
	sram_mem[90402] = 16'b0000000000000000;
	sram_mem[90403] = 16'b0000000000000000;
	sram_mem[90404] = 16'b0000000000000000;
	sram_mem[90405] = 16'b0000000000000000;
	sram_mem[90406] = 16'b0000000000000000;
	sram_mem[90407] = 16'b0000000000000000;
	sram_mem[90408] = 16'b0000000000000000;
	sram_mem[90409] = 16'b0000000000000000;
	sram_mem[90410] = 16'b0000000000000000;
	sram_mem[90411] = 16'b0000000000000000;
	sram_mem[90412] = 16'b0000000000000000;
	sram_mem[90413] = 16'b0000000000000000;
	sram_mem[90414] = 16'b0000000000000000;
	sram_mem[90415] = 16'b0000000000000000;
	sram_mem[90416] = 16'b0000000000000000;
	sram_mem[90417] = 16'b0000000000000000;
	sram_mem[90418] = 16'b0000000000000000;
	sram_mem[90419] = 16'b0000000000000000;
	sram_mem[90420] = 16'b0000000000000000;
	sram_mem[90421] = 16'b0000000000000000;
	sram_mem[90422] = 16'b0000000000000000;
	sram_mem[90423] = 16'b0000000000000000;
	sram_mem[90424] = 16'b0000000000000000;
	sram_mem[90425] = 16'b0000000000000000;
	sram_mem[90426] = 16'b0000000000000000;
	sram_mem[90427] = 16'b0000000000000000;
	sram_mem[90428] = 16'b0000000000000000;
	sram_mem[90429] = 16'b0000000000000000;
	sram_mem[90430] = 16'b0000000000000000;
	sram_mem[90431] = 16'b0000000000000000;
	sram_mem[90432] = 16'b0000000000000000;
	sram_mem[90433] = 16'b0000000000000000;
	sram_mem[90434] = 16'b0000000000000000;
	sram_mem[90435] = 16'b0000000000000000;
	sram_mem[90436] = 16'b0000000000000000;
	sram_mem[90437] = 16'b0000000000000000;
	sram_mem[90438] = 16'b0000000000000000;
	sram_mem[90439] = 16'b0000000000000000;
	sram_mem[90440] = 16'b0000000000000000;
	sram_mem[90441] = 16'b0000000000000000;
	sram_mem[90442] = 16'b0000000000000000;
	sram_mem[90443] = 16'b0000000000000000;
	sram_mem[90444] = 16'b0000000000000000;
	sram_mem[90445] = 16'b0000000000000000;
	sram_mem[90446] = 16'b0000000000000000;
	sram_mem[90447] = 16'b0000000000000000;
	sram_mem[90448] = 16'b0000000000000000;
	sram_mem[90449] = 16'b0000000000000000;
	sram_mem[90450] = 16'b0000000000000000;
	sram_mem[90451] = 16'b0000000000000000;
	sram_mem[90452] = 16'b0000000000000000;
	sram_mem[90453] = 16'b0000000000000000;
	sram_mem[90454] = 16'b0000000000000000;
	sram_mem[90455] = 16'b0000000000000000;
	sram_mem[90456] = 16'b0000000000000000;
	sram_mem[90457] = 16'b0000000000000000;
	sram_mem[90458] = 16'b0000000000000000;
	sram_mem[90459] = 16'b0000000000000000;
	sram_mem[90460] = 16'b0000000000000000;
	sram_mem[90461] = 16'b0000000000000000;
	sram_mem[90462] = 16'b0000000000000000;
	sram_mem[90463] = 16'b0000000000000000;
	sram_mem[90464] = 16'b0000000000000000;
	sram_mem[90465] = 16'b0000000000000000;
	sram_mem[90466] = 16'b0000000000000000;
	sram_mem[90467] = 16'b0000000000000000;
	sram_mem[90468] = 16'b0000000000000000;
	sram_mem[90469] = 16'b0000000000000000;
	sram_mem[90470] = 16'b0000000000000000;
	sram_mem[90471] = 16'b0000000000000000;
	sram_mem[90472] = 16'b0000000000000000;
	sram_mem[90473] = 16'b0000000000000000;
	sram_mem[90474] = 16'b0000000000000000;
	sram_mem[90475] = 16'b0000000000000000;
	sram_mem[90476] = 16'b0000000000000000;
	sram_mem[90477] = 16'b0000000000000000;
	sram_mem[90478] = 16'b0000000000000000;
	sram_mem[90479] = 16'b0000000000000000;
	sram_mem[90480] = 16'b0000000000000000;
	sram_mem[90481] = 16'b0000000000000000;
	sram_mem[90482] = 16'b0000000000000000;
	sram_mem[90483] = 16'b0000000000000000;
	sram_mem[90484] = 16'b0000000000000000;
	sram_mem[90485] = 16'b0000000000000000;
	sram_mem[90486] = 16'b0000000000000000;
	sram_mem[90487] = 16'b0000000000000000;
	sram_mem[90488] = 16'b0000000000000000;
	sram_mem[90489] = 16'b0000000000000000;
	sram_mem[90490] = 16'b0000000000000000;
	sram_mem[90491] = 16'b0000000000000000;
	sram_mem[90492] = 16'b0000000000000000;
	sram_mem[90493] = 16'b0000000000000000;
	sram_mem[90494] = 16'b0000000000000000;
	sram_mem[90495] = 16'b0000000000000000;
	sram_mem[90496] = 16'b0000000000000000;
	sram_mem[90497] = 16'b0000000000000000;
	sram_mem[90498] = 16'b0000000000000000;
	sram_mem[90499] = 16'b0000000000000000;
	sram_mem[90500] = 16'b0000000000000000;
	sram_mem[90501] = 16'b0000000000000000;
	sram_mem[90502] = 16'b0000000000000000;
	sram_mem[90503] = 16'b0000000000000000;
	sram_mem[90504] = 16'b0000000000000000;
	sram_mem[90505] = 16'b0000000000000000;
	sram_mem[90506] = 16'b0000000000000000;
	sram_mem[90507] = 16'b0000000000000000;
	sram_mem[90508] = 16'b0000000000000000;
	sram_mem[90509] = 16'b0000000000000000;
	sram_mem[90510] = 16'b0000000000000000;
	sram_mem[90511] = 16'b0000000000000000;
	sram_mem[90512] = 16'b0000000000000000;
	sram_mem[90513] = 16'b0000000000000000;
	sram_mem[90514] = 16'b0000000000000000;
	sram_mem[90515] = 16'b0000000000000000;
	sram_mem[90516] = 16'b0000000000000000;
	sram_mem[90517] = 16'b0000000000000000;
	sram_mem[90518] = 16'b0000000000000000;
	sram_mem[90519] = 16'b0000000000000000;
	sram_mem[90520] = 16'b0000000000000000;
	sram_mem[90521] = 16'b0000000000000000;
	sram_mem[90522] = 16'b0000000000000000;
	sram_mem[90523] = 16'b0000000000000000;
	sram_mem[90524] = 16'b0000000000000000;
	sram_mem[90525] = 16'b0000000000000000;
	sram_mem[90526] = 16'b0000000000000000;
	sram_mem[90527] = 16'b0000000000000000;
	sram_mem[90528] = 16'b0000000000000000;
	sram_mem[90529] = 16'b0000000000000000;
	sram_mem[90530] = 16'b0000000000000000;
	sram_mem[90531] = 16'b0000000000000000;
	sram_mem[90532] = 16'b0000000000000000;
	sram_mem[90533] = 16'b0000000000000000;
	sram_mem[90534] = 16'b0000000000000000;
	sram_mem[90535] = 16'b0000000000000000;
	sram_mem[90536] = 16'b0000000000000000;
	sram_mem[90537] = 16'b0000000000000000;
	sram_mem[90538] = 16'b0000000000000000;
	sram_mem[90539] = 16'b0000000000000000;
	sram_mem[90540] = 16'b0000000000000000;
	sram_mem[90541] = 16'b0000000000000000;
	sram_mem[90542] = 16'b0000000000000000;
	sram_mem[90543] = 16'b0000000000000000;
	sram_mem[90544] = 16'b0000000000000000;
	sram_mem[90545] = 16'b0000000000000000;
	sram_mem[90546] = 16'b0000000000000000;
	sram_mem[90547] = 16'b0000000000000000;
	sram_mem[90548] = 16'b0000000000000000;
	sram_mem[90549] = 16'b0000000000000000;
	sram_mem[90550] = 16'b0000000000000000;
	sram_mem[90551] = 16'b0000000000000000;
	sram_mem[90552] = 16'b0000000000000000;
	sram_mem[90553] = 16'b0000000000000000;
	sram_mem[90554] = 16'b0000000000000000;
	sram_mem[90555] = 16'b0000000000000000;
	sram_mem[90556] = 16'b0000000000000000;
	sram_mem[90557] = 16'b0000000000000000;
	sram_mem[90558] = 16'b0000000000000000;
	sram_mem[90559] = 16'b0000000000000000;
	sram_mem[90560] = 16'b0000000000000000;
	sram_mem[90561] = 16'b0000000000000000;
	sram_mem[90562] = 16'b0000000000000000;
	sram_mem[90563] = 16'b0000000000000000;
	sram_mem[90564] = 16'b0000000000000000;
	sram_mem[90565] = 16'b0000000000000000;
	sram_mem[90566] = 16'b0000000000000000;
	sram_mem[90567] = 16'b0000000000000000;
	sram_mem[90568] = 16'b0000000000000000;
	sram_mem[90569] = 16'b0000000000000000;
	sram_mem[90570] = 16'b0000000000000000;
	sram_mem[90571] = 16'b0000000000000000;
	sram_mem[90572] = 16'b0000000000000000;
	sram_mem[90573] = 16'b0000000000000000;
	sram_mem[90574] = 16'b0000000000000000;
	sram_mem[90575] = 16'b0000000000000000;
	sram_mem[90576] = 16'b0000000000000000;
	sram_mem[90577] = 16'b0000000000000000;
	sram_mem[90578] = 16'b0000000000000000;
	sram_mem[90579] = 16'b0000000000000000;
	sram_mem[90580] = 16'b0000000000000000;
	sram_mem[90581] = 16'b0000000000000000;
	sram_mem[90582] = 16'b0000000000000000;
	sram_mem[90583] = 16'b0000000000000000;
	sram_mem[90584] = 16'b0000000000000000;
	sram_mem[90585] = 16'b0000000000000000;
	sram_mem[90586] = 16'b0000000000000000;
	sram_mem[90587] = 16'b0000000000000000;
	sram_mem[90588] = 16'b0000000000000000;
	sram_mem[90589] = 16'b0000000000000000;
	sram_mem[90590] = 16'b0000000000000000;
	sram_mem[90591] = 16'b0000000000000000;
	sram_mem[90592] = 16'b0000000000000000;
	sram_mem[90593] = 16'b0000000000000000;
	sram_mem[90594] = 16'b0000000000000000;
	sram_mem[90595] = 16'b0000000000000000;
	sram_mem[90596] = 16'b0000000000000000;
	sram_mem[90597] = 16'b0000000000000000;
	sram_mem[90598] = 16'b0000000000000000;
	sram_mem[90599] = 16'b0000000000000000;
	sram_mem[90600] = 16'b0000000000000000;
	sram_mem[90601] = 16'b0000000000000000;
	sram_mem[90602] = 16'b0000000000000000;
	sram_mem[90603] = 16'b0000000000000000;
	sram_mem[90604] = 16'b0000000000000000;
	sram_mem[90605] = 16'b0000000000000000;
	sram_mem[90606] = 16'b0000000000000000;
	sram_mem[90607] = 16'b0000000000000000;
	sram_mem[90608] = 16'b0000000000000000;
	sram_mem[90609] = 16'b0000000000000000;
	sram_mem[90610] = 16'b0000000000000000;
	sram_mem[90611] = 16'b0000000000000000;
	sram_mem[90612] = 16'b0000000000000000;
	sram_mem[90613] = 16'b0000000000000000;
	sram_mem[90614] = 16'b0000000000000000;
	sram_mem[90615] = 16'b0000000000000000;
	sram_mem[90616] = 16'b0000000000000000;
	sram_mem[90617] = 16'b0000000000000000;
	sram_mem[90618] = 16'b0000000000000000;
	sram_mem[90619] = 16'b0000000000000000;
	sram_mem[90620] = 16'b0000000000000000;
	sram_mem[90621] = 16'b0000000000000000;
	sram_mem[90622] = 16'b0000000000000000;
	sram_mem[90623] = 16'b0000000000000000;
	sram_mem[90624] = 16'b0000000000000000;
	sram_mem[90625] = 16'b0000000000000000;
	sram_mem[90626] = 16'b0000000000000000;
	sram_mem[90627] = 16'b0000000000000000;
	sram_mem[90628] = 16'b0000000000000000;
	sram_mem[90629] = 16'b0000000000000000;
	sram_mem[90630] = 16'b0000000000000000;
	sram_mem[90631] = 16'b0000000000000000;
	sram_mem[90632] = 16'b0000000000000000;
	sram_mem[90633] = 16'b0000000000000000;
	sram_mem[90634] = 16'b0000000000000000;
	sram_mem[90635] = 16'b0000000000000000;
	sram_mem[90636] = 16'b0000000000000000;
	sram_mem[90637] = 16'b0000000000000000;
	sram_mem[90638] = 16'b0000000000000000;
	sram_mem[90639] = 16'b0000000000000000;
	sram_mem[90640] = 16'b0000000000000000;
	sram_mem[90641] = 16'b0000000000000000;
	sram_mem[90642] = 16'b0000000000000000;
	sram_mem[90643] = 16'b0000000000000000;
	sram_mem[90644] = 16'b0000000000000000;
	sram_mem[90645] = 16'b0000000000000000;
	sram_mem[90646] = 16'b0000000000000000;
	sram_mem[90647] = 16'b0000000000000000;
	sram_mem[90648] = 16'b0000000000000000;
	sram_mem[90649] = 16'b0000000000000000;
	sram_mem[90650] = 16'b0000000000000000;
	sram_mem[90651] = 16'b0000000000000000;
	sram_mem[90652] = 16'b0000000000000000;
	sram_mem[90653] = 16'b0000000000000000;
	sram_mem[90654] = 16'b0000000000000000;
	sram_mem[90655] = 16'b0000000000000000;
	sram_mem[90656] = 16'b0000000000000000;
	sram_mem[90657] = 16'b0000000000000000;
	sram_mem[90658] = 16'b0000000000000000;
	sram_mem[90659] = 16'b0000000000000000;
	sram_mem[90660] = 16'b0000000000000000;
	sram_mem[90661] = 16'b0000000000000000;
	sram_mem[90662] = 16'b0000000000000000;
	sram_mem[90663] = 16'b0000000000000000;
	sram_mem[90664] = 16'b0000000000000000;
	sram_mem[90665] = 16'b0000000000000000;
	sram_mem[90666] = 16'b0000000000000000;
	sram_mem[90667] = 16'b0000000000000000;
	sram_mem[90668] = 16'b0000000000000000;
	sram_mem[90669] = 16'b0000000000000000;
	sram_mem[90670] = 16'b0000000000000000;
	sram_mem[90671] = 16'b0000000000000000;
	sram_mem[90672] = 16'b0000000000000000;
	sram_mem[90673] = 16'b0000000000000000;
	sram_mem[90674] = 16'b0000000000000000;
	sram_mem[90675] = 16'b0000000000000000;
	sram_mem[90676] = 16'b0000000000000000;
	sram_mem[90677] = 16'b0000000000000000;
	sram_mem[90678] = 16'b0000000000000000;
	sram_mem[90679] = 16'b0000000000000000;
	sram_mem[90680] = 16'b0000000000000000;
	sram_mem[90681] = 16'b0000000000000000;
	sram_mem[90682] = 16'b0000000000000000;
	sram_mem[90683] = 16'b0000000000000000;
	sram_mem[90684] = 16'b0000000000000000;
	sram_mem[90685] = 16'b0000000000000000;
	sram_mem[90686] = 16'b0000000000000000;
	sram_mem[90687] = 16'b0000000000000000;
	sram_mem[90688] = 16'b0000000000000000;
	sram_mem[90689] = 16'b0000000000000000;
	sram_mem[90690] = 16'b0000000000000000;
	sram_mem[90691] = 16'b0000000000000000;
	sram_mem[90692] = 16'b0000000000000000;
	sram_mem[90693] = 16'b0000000000000000;
	sram_mem[90694] = 16'b0000000000000000;
	sram_mem[90695] = 16'b0000000000000000;
	sram_mem[90696] = 16'b0000000000000000;
	sram_mem[90697] = 16'b0000000000000000;
	sram_mem[90698] = 16'b0000000000000000;
	sram_mem[90699] = 16'b0000000000000000;
	sram_mem[90700] = 16'b0000000000000000;
	sram_mem[90701] = 16'b0000000000000000;
	sram_mem[90702] = 16'b0000000000000000;
	sram_mem[90703] = 16'b0000000000000000;
	sram_mem[90704] = 16'b0000000000000000;
	sram_mem[90705] = 16'b0000000000000000;
	sram_mem[90706] = 16'b0000000000000000;
	sram_mem[90707] = 16'b0000000000000000;
	sram_mem[90708] = 16'b0000000000000000;
	sram_mem[90709] = 16'b0000000000000000;
	sram_mem[90710] = 16'b0000000000000000;
	sram_mem[90711] = 16'b0000000000000000;
	sram_mem[90712] = 16'b0000000000000000;
	sram_mem[90713] = 16'b0000000000000000;
	sram_mem[90714] = 16'b0000000000000000;
	sram_mem[90715] = 16'b0000000000000000;
	sram_mem[90716] = 16'b0000000000000000;
	sram_mem[90717] = 16'b0000000000000000;
	sram_mem[90718] = 16'b0000000000000000;
	sram_mem[90719] = 16'b0000000000000000;
	sram_mem[90720] = 16'b0000000000000000;
	sram_mem[90721] = 16'b0000000000000000;
	sram_mem[90722] = 16'b0000000000000000;
	sram_mem[90723] = 16'b0000000000000000;
	sram_mem[90724] = 16'b0000000000000000;
	sram_mem[90725] = 16'b0000000000000000;
	sram_mem[90726] = 16'b0000000000000000;
	sram_mem[90727] = 16'b0000000000000000;
	sram_mem[90728] = 16'b0000000000000000;
	sram_mem[90729] = 16'b0000000000000000;
	sram_mem[90730] = 16'b0000000000000000;
	sram_mem[90731] = 16'b0000000000000000;
	sram_mem[90732] = 16'b0000000000000000;
	sram_mem[90733] = 16'b0000000000000000;
	sram_mem[90734] = 16'b0000000000000000;
	sram_mem[90735] = 16'b0000000000000000;
	sram_mem[90736] = 16'b0000000000000000;
	sram_mem[90737] = 16'b0000000000000000;
	sram_mem[90738] = 16'b0000000000000000;
	sram_mem[90739] = 16'b0000000000000000;
	sram_mem[90740] = 16'b0000000000000000;
	sram_mem[90741] = 16'b0000000000000000;
	sram_mem[90742] = 16'b0000000000000000;
	sram_mem[90743] = 16'b0000000000000000;
	sram_mem[90744] = 16'b0000000000000000;
	sram_mem[90745] = 16'b0000000000000000;
	sram_mem[90746] = 16'b0000000000000000;
	sram_mem[90747] = 16'b0000000000000000;
	sram_mem[90748] = 16'b0000000000000000;
	sram_mem[90749] = 16'b0000000000000000;
	sram_mem[90750] = 16'b0000000000000000;
	sram_mem[90751] = 16'b0000000000000000;
	sram_mem[90752] = 16'b0000000000000000;
	sram_mem[90753] = 16'b0000000000000000;
	sram_mem[90754] = 16'b0000000000000000;
	sram_mem[90755] = 16'b0000000000000000;
	sram_mem[90756] = 16'b0000000000000000;
	sram_mem[90757] = 16'b0000000000000000;
	sram_mem[90758] = 16'b0000000000000000;
	sram_mem[90759] = 16'b0000000000000000;
	sram_mem[90760] = 16'b0000000000000000;
	sram_mem[90761] = 16'b0000000000000000;
	sram_mem[90762] = 16'b0000000000000000;
	sram_mem[90763] = 16'b0000000000000000;
	sram_mem[90764] = 16'b0000000000000000;
	sram_mem[90765] = 16'b0000000000000000;
	sram_mem[90766] = 16'b0000000000000000;
	sram_mem[90767] = 16'b0000000000000000;
	sram_mem[90768] = 16'b0000000000000000;
	sram_mem[90769] = 16'b0000000000000000;
	sram_mem[90770] = 16'b0000000000000000;
	sram_mem[90771] = 16'b0000000000000000;
	sram_mem[90772] = 16'b0000000000000000;
	sram_mem[90773] = 16'b0000000000000000;
	sram_mem[90774] = 16'b0000000000000000;
	sram_mem[90775] = 16'b0000000000000000;
	sram_mem[90776] = 16'b0000000000000000;
	sram_mem[90777] = 16'b0000000000000000;
	sram_mem[90778] = 16'b0000000000000000;
	sram_mem[90779] = 16'b0000000000000000;
	sram_mem[90780] = 16'b0000000000000000;
	sram_mem[90781] = 16'b0000000000000000;
	sram_mem[90782] = 16'b0000000000000000;
	sram_mem[90783] = 16'b0000000000000000;
	sram_mem[90784] = 16'b0000000000000000;
	sram_mem[90785] = 16'b0000000000000000;
	sram_mem[90786] = 16'b0000000000000000;
	sram_mem[90787] = 16'b0000000000000000;
	sram_mem[90788] = 16'b0000000000000000;
	sram_mem[90789] = 16'b0000000000000000;
	sram_mem[90790] = 16'b0000000000000000;
	sram_mem[90791] = 16'b0000000000000000;
	sram_mem[90792] = 16'b0000000000000000;
	sram_mem[90793] = 16'b0000000000000000;
	sram_mem[90794] = 16'b0000000000000000;
	sram_mem[90795] = 16'b0000000000000000;
	sram_mem[90796] = 16'b0000000000000000;
	sram_mem[90797] = 16'b0000000000000000;
	sram_mem[90798] = 16'b0000000000000000;
	sram_mem[90799] = 16'b0000000000000000;
	sram_mem[90800] = 16'b0000000000000000;
	sram_mem[90801] = 16'b0000000000000000;
	sram_mem[90802] = 16'b0000000000000000;
	sram_mem[90803] = 16'b0000000000000000;
	sram_mem[90804] = 16'b0000000000000000;
	sram_mem[90805] = 16'b0000000000000000;
	sram_mem[90806] = 16'b0000000000000000;
	sram_mem[90807] = 16'b0000000000000000;
	sram_mem[90808] = 16'b0000000000000000;
	sram_mem[90809] = 16'b0000000000000000;
	sram_mem[90810] = 16'b0000000000000000;
	sram_mem[90811] = 16'b0000000000000000;
	sram_mem[90812] = 16'b0000000000000000;
	sram_mem[90813] = 16'b0000000000000000;
	sram_mem[90814] = 16'b0000000000000000;
	sram_mem[90815] = 16'b0000000000000000;
	sram_mem[90816] = 16'b0000000000000000;
	sram_mem[90817] = 16'b0000000000000000;
	sram_mem[90818] = 16'b0000000000000000;
	sram_mem[90819] = 16'b0000000000000000;
	sram_mem[90820] = 16'b0000000000000000;
	sram_mem[90821] = 16'b0000000000000000;
	sram_mem[90822] = 16'b0000000000000000;
	sram_mem[90823] = 16'b0000000000000000;
	sram_mem[90824] = 16'b0000000000000000;
	sram_mem[90825] = 16'b0000000000000000;
	sram_mem[90826] = 16'b0000000000000000;
	sram_mem[90827] = 16'b0000000000000000;
	sram_mem[90828] = 16'b0000000000000000;
	sram_mem[90829] = 16'b0000000000000000;
	sram_mem[90830] = 16'b0000000000000000;
	sram_mem[90831] = 16'b0000000000000000;
	sram_mem[90832] = 16'b0000000000000000;
	sram_mem[90833] = 16'b0000000000000000;
	sram_mem[90834] = 16'b0000000000000000;
	sram_mem[90835] = 16'b0000000000000000;
	sram_mem[90836] = 16'b0000000000000000;
	sram_mem[90837] = 16'b0000000000000000;
	sram_mem[90838] = 16'b0000000000000000;
	sram_mem[90839] = 16'b0000000000000000;
	sram_mem[90840] = 16'b0000000000000000;
	sram_mem[90841] = 16'b0000000000000000;
	sram_mem[90842] = 16'b0000000000000000;
	sram_mem[90843] = 16'b0000000000000000;
	sram_mem[90844] = 16'b0000000000000000;
	sram_mem[90845] = 16'b0000000000000000;
	sram_mem[90846] = 16'b0000000000000000;
	sram_mem[90847] = 16'b0000000000000000;
	sram_mem[90848] = 16'b0000000000000000;
	sram_mem[90849] = 16'b0000000000000000;
	sram_mem[90850] = 16'b0000000000000000;
	sram_mem[90851] = 16'b0000000000000000;
	sram_mem[90852] = 16'b0000000000000000;
	sram_mem[90853] = 16'b0000000000000000;
	sram_mem[90854] = 16'b0000000000000000;
	sram_mem[90855] = 16'b0000000000000000;
	sram_mem[90856] = 16'b0000000000000000;
	sram_mem[90857] = 16'b0000000000000000;
	sram_mem[90858] = 16'b0000000000000000;
	sram_mem[90859] = 16'b0000000000000000;
	sram_mem[90860] = 16'b0000000000000000;
	sram_mem[90861] = 16'b0000000000000000;
	sram_mem[90862] = 16'b0000000000000000;
	sram_mem[90863] = 16'b0000000000000000;
	sram_mem[90864] = 16'b0000000000000000;
	sram_mem[90865] = 16'b0000000000000000;
	sram_mem[90866] = 16'b0000000000000000;
	sram_mem[90867] = 16'b0000000000000000;
	sram_mem[90868] = 16'b0000000000000000;
	sram_mem[90869] = 16'b0000000000000000;
	sram_mem[90870] = 16'b0000000000000000;
	sram_mem[90871] = 16'b0000000000000000;
	sram_mem[90872] = 16'b0000000000000000;
	sram_mem[90873] = 16'b0000000000000000;
	sram_mem[90874] = 16'b0000000000000000;
	sram_mem[90875] = 16'b0000000000000000;
	sram_mem[90876] = 16'b0000000000000000;
	sram_mem[90877] = 16'b0000000000000000;
	sram_mem[90878] = 16'b0000000000000000;
	sram_mem[90879] = 16'b0000000000000000;
	sram_mem[90880] = 16'b0000000000000000;
	sram_mem[90881] = 16'b0000000000000000;
	sram_mem[90882] = 16'b0000000000000000;
	sram_mem[90883] = 16'b0000000000000000;
	sram_mem[90884] = 16'b0000000000000000;
	sram_mem[90885] = 16'b0000000000000000;
	sram_mem[90886] = 16'b0000000000000000;
	sram_mem[90887] = 16'b0000000000000000;
	sram_mem[90888] = 16'b0000000000000000;
	sram_mem[90889] = 16'b0000000000000000;
	sram_mem[90890] = 16'b0000000000000000;
	sram_mem[90891] = 16'b0000000000000000;
	sram_mem[90892] = 16'b0000000000000000;
	sram_mem[90893] = 16'b0000000000000000;
	sram_mem[90894] = 16'b0000000000000000;
	sram_mem[90895] = 16'b0000000000000000;
	sram_mem[90896] = 16'b0000000000000000;
	sram_mem[90897] = 16'b0000000000000000;
	sram_mem[90898] = 16'b0000000000000000;
	sram_mem[90899] = 16'b0000000000000000;
	sram_mem[90900] = 16'b0000000000000000;
	sram_mem[90901] = 16'b0000000000000000;
	sram_mem[90902] = 16'b0000000000000000;
	sram_mem[90903] = 16'b0000000000000000;
	sram_mem[90904] = 16'b0000000000000000;
	sram_mem[90905] = 16'b0000000000000000;
	sram_mem[90906] = 16'b0000000000000000;
	sram_mem[90907] = 16'b0000000000000000;
	sram_mem[90908] = 16'b0000000000000000;
	sram_mem[90909] = 16'b0000000000000000;
	sram_mem[90910] = 16'b0000000000000000;
	sram_mem[90911] = 16'b0000000000000000;
	sram_mem[90912] = 16'b0000000000000000;
	sram_mem[90913] = 16'b0000000000000000;
	sram_mem[90914] = 16'b0000000000000000;
	sram_mem[90915] = 16'b0000000000000000;
	sram_mem[90916] = 16'b0000000000000000;
	sram_mem[90917] = 16'b0000000000000000;
	sram_mem[90918] = 16'b0000000000000000;
	sram_mem[90919] = 16'b0000000000000000;
	sram_mem[90920] = 16'b0000000000000000;
	sram_mem[90921] = 16'b0000000000000000;
	sram_mem[90922] = 16'b0000000000000000;
	sram_mem[90923] = 16'b0000000000000000;
	sram_mem[90924] = 16'b0000000000000000;
	sram_mem[90925] = 16'b0000000000000000;
	sram_mem[90926] = 16'b0000000000000000;
	sram_mem[90927] = 16'b0000000000000000;
	sram_mem[90928] = 16'b0000000000000000;
	sram_mem[90929] = 16'b0000000000000000;
	sram_mem[90930] = 16'b0000000000000000;
	sram_mem[90931] = 16'b0000000000000000;
	sram_mem[90932] = 16'b0000000000000000;
	sram_mem[90933] = 16'b0000000000000000;
	sram_mem[90934] = 16'b0000000000000000;
	sram_mem[90935] = 16'b0000000000000000;
	sram_mem[90936] = 16'b0000000000000000;
	sram_mem[90937] = 16'b0000000000000000;
	sram_mem[90938] = 16'b0000000000000000;
	sram_mem[90939] = 16'b0000000000000000;
	sram_mem[90940] = 16'b0000000000000000;
	sram_mem[90941] = 16'b0000000000000000;
	sram_mem[90942] = 16'b0000000000000000;
	sram_mem[90943] = 16'b0000000000000000;
	sram_mem[90944] = 16'b0000000000000000;
	sram_mem[90945] = 16'b0000000000000000;
	sram_mem[90946] = 16'b0000000000000000;
	sram_mem[90947] = 16'b0000000000000000;
	sram_mem[90948] = 16'b0000000000000000;
	sram_mem[90949] = 16'b0000000000000000;
	sram_mem[90950] = 16'b0000000000000000;
	sram_mem[90951] = 16'b0000000000000000;
	sram_mem[90952] = 16'b0000000000000000;
	sram_mem[90953] = 16'b0000000000000000;
	sram_mem[90954] = 16'b0000000000000000;
	sram_mem[90955] = 16'b0000000000000000;
	sram_mem[90956] = 16'b0000000000000000;
	sram_mem[90957] = 16'b0000000000000000;
	sram_mem[90958] = 16'b0000000000000000;
	sram_mem[90959] = 16'b0000000000000000;
	sram_mem[90960] = 16'b0000000000000000;
	sram_mem[90961] = 16'b0000000000000000;
	sram_mem[90962] = 16'b0000000000000000;
	sram_mem[90963] = 16'b0000000000000000;
	sram_mem[90964] = 16'b0000000000000000;
	sram_mem[90965] = 16'b0000000000000000;
	sram_mem[90966] = 16'b0000000000000000;
	sram_mem[90967] = 16'b0000000000000000;
	sram_mem[90968] = 16'b0000000000000000;
	sram_mem[90969] = 16'b0000000000000000;
	sram_mem[90970] = 16'b0000000000000000;
	sram_mem[90971] = 16'b0000000000000000;
	sram_mem[90972] = 16'b0000000000000000;
	sram_mem[90973] = 16'b0000000000000000;
	sram_mem[90974] = 16'b0000000000000000;
	sram_mem[90975] = 16'b0000000000000000;
	sram_mem[90976] = 16'b0000000000000000;
	sram_mem[90977] = 16'b0000000000000000;
	sram_mem[90978] = 16'b0000000000000000;
	sram_mem[90979] = 16'b0000000000000000;
	sram_mem[90980] = 16'b0000000000000000;
	sram_mem[90981] = 16'b0000000000000000;
	sram_mem[90982] = 16'b0000000000000000;
	sram_mem[90983] = 16'b0000000000000000;
	sram_mem[90984] = 16'b0000000000000000;
	sram_mem[90985] = 16'b0000000000000000;
	sram_mem[90986] = 16'b0000000000000000;
	sram_mem[90987] = 16'b0000000000000000;
	sram_mem[90988] = 16'b0000000000000000;
	sram_mem[90989] = 16'b0000000000000000;
	sram_mem[90990] = 16'b0000000000000000;
	sram_mem[90991] = 16'b0000000000000000;
	sram_mem[90992] = 16'b0000000000000000;
	sram_mem[90993] = 16'b0000000000000000;
	sram_mem[90994] = 16'b0000000000000000;
	sram_mem[90995] = 16'b0000000000000000;
	sram_mem[90996] = 16'b0000000000000000;
	sram_mem[90997] = 16'b0000000000000000;
	sram_mem[90998] = 16'b0000000000000000;
	sram_mem[90999] = 16'b0000000000000000;
	sram_mem[91000] = 16'b0000000000000000;
	sram_mem[91001] = 16'b0000000000000000;
	sram_mem[91002] = 16'b0000000000000000;
	sram_mem[91003] = 16'b0000000000000000;
	sram_mem[91004] = 16'b0000000000000000;
	sram_mem[91005] = 16'b0000000000000000;
	sram_mem[91006] = 16'b0000000000000000;
	sram_mem[91007] = 16'b0000000000000000;
	sram_mem[91008] = 16'b0000000000000000;
	sram_mem[91009] = 16'b0000000000000000;
	sram_mem[91010] = 16'b0000000000000000;
	sram_mem[91011] = 16'b0000000000000000;
	sram_mem[91012] = 16'b0000000000000000;
	sram_mem[91013] = 16'b0000000000000000;
	sram_mem[91014] = 16'b0000000000000000;
	sram_mem[91015] = 16'b0000000000000000;
	sram_mem[91016] = 16'b0000000000000000;
	sram_mem[91017] = 16'b0000000000000000;
	sram_mem[91018] = 16'b0000000000000000;
	sram_mem[91019] = 16'b0000000000000000;
	sram_mem[91020] = 16'b0000000000000000;
	sram_mem[91021] = 16'b0000000000000000;
	sram_mem[91022] = 16'b0000000000000000;
	sram_mem[91023] = 16'b0000000000000000;
	sram_mem[91024] = 16'b0000000000000000;
	sram_mem[91025] = 16'b0000000000000000;
	sram_mem[91026] = 16'b0000000000000000;
	sram_mem[91027] = 16'b0000000000000000;
	sram_mem[91028] = 16'b0000000000000000;
	sram_mem[91029] = 16'b0000000000000000;
	sram_mem[91030] = 16'b0000000000000000;
	sram_mem[91031] = 16'b0000000000000000;
	sram_mem[91032] = 16'b0000000000000000;
	sram_mem[91033] = 16'b0000000000000000;
	sram_mem[91034] = 16'b0000000000000000;
	sram_mem[91035] = 16'b0000000000000000;
	sram_mem[91036] = 16'b0000000000000000;
	sram_mem[91037] = 16'b0000000000000000;
	sram_mem[91038] = 16'b0000000000000000;
	sram_mem[91039] = 16'b0000000000000000;
	sram_mem[91040] = 16'b0000000000000000;
	sram_mem[91041] = 16'b0000000000000000;
	sram_mem[91042] = 16'b0000000000000000;
	sram_mem[91043] = 16'b0000000000000000;
	sram_mem[91044] = 16'b0000000000000000;
	sram_mem[91045] = 16'b0000000000000000;
	sram_mem[91046] = 16'b0000000000000000;
	sram_mem[91047] = 16'b0000000000000000;
	sram_mem[91048] = 16'b0000000000000000;
	sram_mem[91049] = 16'b0000000000000000;
	sram_mem[91050] = 16'b0000000000000000;
	sram_mem[91051] = 16'b0000000000000000;
	sram_mem[91052] = 16'b0000000000000000;
	sram_mem[91053] = 16'b0000000000000000;
	sram_mem[91054] = 16'b0000000000000000;
	sram_mem[91055] = 16'b0000000000000000;
	sram_mem[91056] = 16'b0000000000000000;
	sram_mem[91057] = 16'b0000000000000000;
	sram_mem[91058] = 16'b0000000000000000;
	sram_mem[91059] = 16'b0000000000000000;
	sram_mem[91060] = 16'b0000000000000000;
	sram_mem[91061] = 16'b0000000000000000;
	sram_mem[91062] = 16'b0000000000000000;
	sram_mem[91063] = 16'b0000000000000000;
	sram_mem[91064] = 16'b0000000000000000;
	sram_mem[91065] = 16'b0000000000000000;
	sram_mem[91066] = 16'b0000000000000000;
	sram_mem[91067] = 16'b0000000000000000;
	sram_mem[91068] = 16'b0000000000000000;
	sram_mem[91069] = 16'b0000000000000000;
	sram_mem[91070] = 16'b0000000000000000;
	sram_mem[91071] = 16'b0000000000000000;
	sram_mem[91072] = 16'b0000000000000000;
	sram_mem[91073] = 16'b0000000000000000;
	sram_mem[91074] = 16'b0000000000000000;
	sram_mem[91075] = 16'b0000000000000000;
	sram_mem[91076] = 16'b0000000000000000;
	sram_mem[91077] = 16'b0000000000000000;
	sram_mem[91078] = 16'b0000000000000000;
	sram_mem[91079] = 16'b0000000000000000;
	sram_mem[91080] = 16'b0000000000000000;
	sram_mem[91081] = 16'b0000000000000000;
	sram_mem[91082] = 16'b0000000000000000;
	sram_mem[91083] = 16'b0000000000000000;
	sram_mem[91084] = 16'b0000000000000000;
	sram_mem[91085] = 16'b0000000000000000;
	sram_mem[91086] = 16'b0000000000000000;
	sram_mem[91087] = 16'b0000000000000000;
	sram_mem[91088] = 16'b0000000000000000;
	sram_mem[91089] = 16'b0000000000000000;
	sram_mem[91090] = 16'b0000000000000000;
	sram_mem[91091] = 16'b0000000000000000;
	sram_mem[91092] = 16'b0000000000000000;
	sram_mem[91093] = 16'b0000000000000000;
	sram_mem[91094] = 16'b0000000000000000;
	sram_mem[91095] = 16'b0000000000000000;
	sram_mem[91096] = 16'b0000000000000000;
	sram_mem[91097] = 16'b0000000000000000;
	sram_mem[91098] = 16'b0000000000000000;
	sram_mem[91099] = 16'b0000000000000000;
	sram_mem[91100] = 16'b0000000000000000;
	sram_mem[91101] = 16'b0000000000000000;
	sram_mem[91102] = 16'b0000000000000000;
	sram_mem[91103] = 16'b0000000000000000;
	sram_mem[91104] = 16'b0000000000000000;
	sram_mem[91105] = 16'b0000000000000000;
	sram_mem[91106] = 16'b0000000000000000;
	sram_mem[91107] = 16'b0000000000000000;
	sram_mem[91108] = 16'b0000000000000000;
	sram_mem[91109] = 16'b0000000000000000;
	sram_mem[91110] = 16'b0000000000000000;
	sram_mem[91111] = 16'b0000000000000000;
	sram_mem[91112] = 16'b0000000000000000;
	sram_mem[91113] = 16'b0000000000000000;
	sram_mem[91114] = 16'b0000000000000000;
	sram_mem[91115] = 16'b0000000000000000;
	sram_mem[91116] = 16'b0000000000000000;
	sram_mem[91117] = 16'b0000000000000000;
	sram_mem[91118] = 16'b0000000000000000;
	sram_mem[91119] = 16'b0000000000000000;
	sram_mem[91120] = 16'b0000000000000000;
	sram_mem[91121] = 16'b0000000000000000;
	sram_mem[91122] = 16'b0000000000000000;
	sram_mem[91123] = 16'b0000000000000000;
	sram_mem[91124] = 16'b0000000000000000;
	sram_mem[91125] = 16'b0000000000000000;
	sram_mem[91126] = 16'b0000000000000000;
	sram_mem[91127] = 16'b0000000000000000;
	sram_mem[91128] = 16'b0000000000000000;
	sram_mem[91129] = 16'b0000000000000000;
	sram_mem[91130] = 16'b0000000000000000;
	sram_mem[91131] = 16'b0000000000000000;
	sram_mem[91132] = 16'b0000000000000000;
	sram_mem[91133] = 16'b0000000000000000;
	sram_mem[91134] = 16'b0000000000000000;
	sram_mem[91135] = 16'b0000000000000000;
	sram_mem[91136] = 16'b0000000000000000;
	sram_mem[91137] = 16'b0000000000000000;
	sram_mem[91138] = 16'b0000000000000000;
	sram_mem[91139] = 16'b0000000000000000;
	sram_mem[91140] = 16'b0000000000000000;
	sram_mem[91141] = 16'b0000000000000000;
	sram_mem[91142] = 16'b0000000000000000;
	sram_mem[91143] = 16'b0000000000000000;
	sram_mem[91144] = 16'b0000000000000000;
	sram_mem[91145] = 16'b0000000000000000;
	sram_mem[91146] = 16'b0000000000000000;
	sram_mem[91147] = 16'b0000000000000000;
	sram_mem[91148] = 16'b0000000000000000;
	sram_mem[91149] = 16'b0000000000000000;
	sram_mem[91150] = 16'b0000000000000000;
	sram_mem[91151] = 16'b0000000000000000;
	sram_mem[91152] = 16'b0000000000000000;
	sram_mem[91153] = 16'b0000000000000000;
	sram_mem[91154] = 16'b0000000000000000;
	sram_mem[91155] = 16'b0000000000000000;
	sram_mem[91156] = 16'b0000000000000000;
	sram_mem[91157] = 16'b0000000000000000;
	sram_mem[91158] = 16'b0000000000000000;
	sram_mem[91159] = 16'b0000000000000000;
	sram_mem[91160] = 16'b0000000000000000;
	sram_mem[91161] = 16'b0000000000000000;
	sram_mem[91162] = 16'b0000000000000000;
	sram_mem[91163] = 16'b0000000000000000;
	sram_mem[91164] = 16'b0000000000000000;
	sram_mem[91165] = 16'b0000000000000000;
	sram_mem[91166] = 16'b0000000000000000;
	sram_mem[91167] = 16'b0000000000000000;
	sram_mem[91168] = 16'b0000000000000000;
	sram_mem[91169] = 16'b0000000000000000;
	sram_mem[91170] = 16'b0000000000000000;
	sram_mem[91171] = 16'b0000000000000000;
	sram_mem[91172] = 16'b0000000000000000;
	sram_mem[91173] = 16'b0000000000000000;
	sram_mem[91174] = 16'b0000000000000000;
	sram_mem[91175] = 16'b0000000000000000;
	sram_mem[91176] = 16'b0000000000000000;
	sram_mem[91177] = 16'b0000000000000000;
	sram_mem[91178] = 16'b0000000000000000;
	sram_mem[91179] = 16'b0000000000000000;
	sram_mem[91180] = 16'b0000000000000000;
	sram_mem[91181] = 16'b0000000000000000;
	sram_mem[91182] = 16'b0000000000000000;
	sram_mem[91183] = 16'b0000000000000000;
	sram_mem[91184] = 16'b0000000000000000;
	sram_mem[91185] = 16'b0000000000000000;
	sram_mem[91186] = 16'b0000000000000000;
	sram_mem[91187] = 16'b0000000000000000;
	sram_mem[91188] = 16'b0000000000000000;
	sram_mem[91189] = 16'b0000000000000000;
	sram_mem[91190] = 16'b0000000000000000;
	sram_mem[91191] = 16'b0000000000000000;
	sram_mem[91192] = 16'b0000000000000000;
	sram_mem[91193] = 16'b0000000000000000;
	sram_mem[91194] = 16'b0000000000000000;
	sram_mem[91195] = 16'b0000000000000000;
	sram_mem[91196] = 16'b0000000000000000;
	sram_mem[91197] = 16'b0000000000000000;
	sram_mem[91198] = 16'b0000000000000000;
	sram_mem[91199] = 16'b0000000000000000;
	sram_mem[91200] = 16'b0000000000000000;
	sram_mem[91201] = 16'b0000000000000000;
	sram_mem[91202] = 16'b0000000000000000;
	sram_mem[91203] = 16'b0000000000000000;
	sram_mem[91204] = 16'b0000000000000000;
	sram_mem[91205] = 16'b0000000000000000;
	sram_mem[91206] = 16'b0000000000000000;
	sram_mem[91207] = 16'b0000000000000000;
	sram_mem[91208] = 16'b0000000000000000;
	sram_mem[91209] = 16'b0000000000000000;
	sram_mem[91210] = 16'b0000000000000000;
	sram_mem[91211] = 16'b0000000000000000;
	sram_mem[91212] = 16'b0000000000000000;
	sram_mem[91213] = 16'b0000000000000000;
	sram_mem[91214] = 16'b0000000000000000;
	sram_mem[91215] = 16'b0000000000000000;
	sram_mem[91216] = 16'b0000000000000000;
	sram_mem[91217] = 16'b0000000000000000;
	sram_mem[91218] = 16'b0000000000000000;
	sram_mem[91219] = 16'b0000000000000000;
	sram_mem[91220] = 16'b0000000000000000;
	sram_mem[91221] = 16'b0000000000000000;
	sram_mem[91222] = 16'b0000000000000000;
	sram_mem[91223] = 16'b0000000000000000;
	sram_mem[91224] = 16'b0000000000000000;
	sram_mem[91225] = 16'b0000000000000000;
	sram_mem[91226] = 16'b0000000000000000;
	sram_mem[91227] = 16'b0000000000000000;
	sram_mem[91228] = 16'b0000000000000000;
	sram_mem[91229] = 16'b0000000000000000;
	sram_mem[91230] = 16'b0000000000000000;
	sram_mem[91231] = 16'b0000000000000000;
	sram_mem[91232] = 16'b0000000000000000;
	sram_mem[91233] = 16'b0000000000000000;
	sram_mem[91234] = 16'b0000000000000000;
	sram_mem[91235] = 16'b0000000000000000;
	sram_mem[91236] = 16'b0000000000000000;
	sram_mem[91237] = 16'b0000000000000000;
	sram_mem[91238] = 16'b0000000000000000;
	sram_mem[91239] = 16'b0000000000000000;
	sram_mem[91240] = 16'b0000000000000000;
	sram_mem[91241] = 16'b0000000000000000;
	sram_mem[91242] = 16'b0000000000000000;
	sram_mem[91243] = 16'b0000000000000000;
	sram_mem[91244] = 16'b0000000000000000;
	sram_mem[91245] = 16'b0000000000000000;
	sram_mem[91246] = 16'b0000000000000000;
	sram_mem[91247] = 16'b0000000000000000;
	sram_mem[91248] = 16'b0000000000000000;
	sram_mem[91249] = 16'b0000000000000000;
	sram_mem[91250] = 16'b0000000000000000;
	sram_mem[91251] = 16'b0000000000000000;
	sram_mem[91252] = 16'b0000000000000000;
	sram_mem[91253] = 16'b0000000000000000;
	sram_mem[91254] = 16'b0000000000000000;
	sram_mem[91255] = 16'b0000000000000000;
	sram_mem[91256] = 16'b0000000000000000;
	sram_mem[91257] = 16'b0000000000000000;
	sram_mem[91258] = 16'b0000000000000000;
	sram_mem[91259] = 16'b0000000000000000;
	sram_mem[91260] = 16'b0000000000000000;
	sram_mem[91261] = 16'b0000000000000000;
	sram_mem[91262] = 16'b0000000000000000;
	sram_mem[91263] = 16'b0000000000000000;
	sram_mem[91264] = 16'b0000000000000000;
	sram_mem[91265] = 16'b0000000000000000;
	sram_mem[91266] = 16'b0000000000000000;
	sram_mem[91267] = 16'b0000000000000000;
	sram_mem[91268] = 16'b0000000000000000;
	sram_mem[91269] = 16'b0000000000000000;
	sram_mem[91270] = 16'b0000000000000000;
	sram_mem[91271] = 16'b0000000000000000;
	sram_mem[91272] = 16'b0000000000000000;
	sram_mem[91273] = 16'b0000000000000000;
	sram_mem[91274] = 16'b0000000000000000;
	sram_mem[91275] = 16'b0000000000000000;
	sram_mem[91276] = 16'b0000000000000000;
	sram_mem[91277] = 16'b0000000000000000;
	sram_mem[91278] = 16'b0000000000000000;
	sram_mem[91279] = 16'b0000000000000000;
	sram_mem[91280] = 16'b0000000000000000;
	sram_mem[91281] = 16'b0000000000000000;
	sram_mem[91282] = 16'b0000000000000000;
	sram_mem[91283] = 16'b0000000000000000;
	sram_mem[91284] = 16'b0000000000000000;
	sram_mem[91285] = 16'b0000000000000000;
	sram_mem[91286] = 16'b0000000000000000;
	sram_mem[91287] = 16'b0000000000000000;
	sram_mem[91288] = 16'b0000000000000000;
	sram_mem[91289] = 16'b0000000000000000;
	sram_mem[91290] = 16'b0000000000000000;
	sram_mem[91291] = 16'b0000000000000000;
	sram_mem[91292] = 16'b0000000000000000;
	sram_mem[91293] = 16'b0000000000000000;
	sram_mem[91294] = 16'b0000000000000000;
	sram_mem[91295] = 16'b0000000000000000;
	sram_mem[91296] = 16'b0000000000000000;
	sram_mem[91297] = 16'b0000000000000000;
	sram_mem[91298] = 16'b0000000000000000;
	sram_mem[91299] = 16'b0000000000000000;
	sram_mem[91300] = 16'b0000000000000000;
	sram_mem[91301] = 16'b0000000000000000;
	sram_mem[91302] = 16'b0000000000000000;
	sram_mem[91303] = 16'b0000000000000000;
	sram_mem[91304] = 16'b0000000000000000;
	sram_mem[91305] = 16'b0000000000000000;
	sram_mem[91306] = 16'b0000000000000000;
	sram_mem[91307] = 16'b0000000000000000;
	sram_mem[91308] = 16'b0000000000000000;
	sram_mem[91309] = 16'b0000000000000000;
	sram_mem[91310] = 16'b0000000000000000;
	sram_mem[91311] = 16'b0000000000000000;
	sram_mem[91312] = 16'b0000000000000000;
	sram_mem[91313] = 16'b0000000000000000;
	sram_mem[91314] = 16'b0000000000000000;
	sram_mem[91315] = 16'b0000000000000000;
	sram_mem[91316] = 16'b0000000000000000;
	sram_mem[91317] = 16'b0000000000000000;
	sram_mem[91318] = 16'b0000000000000000;
	sram_mem[91319] = 16'b0000000000000000;
	sram_mem[91320] = 16'b0000000000000000;
	sram_mem[91321] = 16'b0000000000000000;
	sram_mem[91322] = 16'b0000000000000000;
	sram_mem[91323] = 16'b0000000000000000;
	sram_mem[91324] = 16'b0000000000000000;
	sram_mem[91325] = 16'b0000000000000000;
	sram_mem[91326] = 16'b0000000000000000;
	sram_mem[91327] = 16'b0000000000000000;
	sram_mem[91328] = 16'b0000000000000000;
	sram_mem[91329] = 16'b0000000000000000;
	sram_mem[91330] = 16'b0000000000000000;
	sram_mem[91331] = 16'b0000000000000000;
	sram_mem[91332] = 16'b0000000000000000;
	sram_mem[91333] = 16'b0000000000000000;
	sram_mem[91334] = 16'b0000000000000000;
	sram_mem[91335] = 16'b0000000000000000;
	sram_mem[91336] = 16'b0000000000000000;
	sram_mem[91337] = 16'b0000000000000000;
	sram_mem[91338] = 16'b0000000000000000;
	sram_mem[91339] = 16'b0000000000000000;
	sram_mem[91340] = 16'b0000000000000000;
	sram_mem[91341] = 16'b0000000000000000;
	sram_mem[91342] = 16'b0000000000000000;
	sram_mem[91343] = 16'b0000000000000000;
	sram_mem[91344] = 16'b0000000000000000;
	sram_mem[91345] = 16'b0000000000000000;
	sram_mem[91346] = 16'b0000000000000000;
	sram_mem[91347] = 16'b0000000000000000;
	sram_mem[91348] = 16'b0000000000000000;
	sram_mem[91349] = 16'b0000000000000000;
	sram_mem[91350] = 16'b0000000000000000;
	sram_mem[91351] = 16'b0000000000000000;
	sram_mem[91352] = 16'b0000000000000000;
	sram_mem[91353] = 16'b0000000000000000;
	sram_mem[91354] = 16'b0000000000000000;
	sram_mem[91355] = 16'b0000000000000000;
	sram_mem[91356] = 16'b0000000000000000;
	sram_mem[91357] = 16'b0000000000000000;
	sram_mem[91358] = 16'b0000000000000000;
	sram_mem[91359] = 16'b0000000000000000;
	sram_mem[91360] = 16'b0000000000000000;
	sram_mem[91361] = 16'b0000000000000000;
	sram_mem[91362] = 16'b0000000000000000;
	sram_mem[91363] = 16'b0000000000000000;
	sram_mem[91364] = 16'b0000000000000000;
	sram_mem[91365] = 16'b0000000000000000;
	sram_mem[91366] = 16'b0000000000000000;
	sram_mem[91367] = 16'b0000000000000000;
	sram_mem[91368] = 16'b0000000000000000;
	sram_mem[91369] = 16'b0000000000000000;
	sram_mem[91370] = 16'b0000000000000000;
	sram_mem[91371] = 16'b0000000000000000;
	sram_mem[91372] = 16'b0000000000000000;
	sram_mem[91373] = 16'b0000000000000000;
	sram_mem[91374] = 16'b0000000000000000;
	sram_mem[91375] = 16'b0000000000000000;
	sram_mem[91376] = 16'b0000000000000000;
	sram_mem[91377] = 16'b0000000000000000;
	sram_mem[91378] = 16'b0000000000000000;
	sram_mem[91379] = 16'b0000000000000000;
	sram_mem[91380] = 16'b0000000000000000;
	sram_mem[91381] = 16'b0000000000000000;
	sram_mem[91382] = 16'b0000000000000000;
	sram_mem[91383] = 16'b0000000000000000;
	sram_mem[91384] = 16'b0000000000000000;
	sram_mem[91385] = 16'b0000000000000000;
	sram_mem[91386] = 16'b0000000000000000;
	sram_mem[91387] = 16'b0000000000000000;
	sram_mem[91388] = 16'b0000000000000000;
	sram_mem[91389] = 16'b0000000000000000;
	sram_mem[91390] = 16'b0000000000000000;
	sram_mem[91391] = 16'b0000000000000000;
	sram_mem[91392] = 16'b0000000000000000;
	sram_mem[91393] = 16'b0000000000000000;
	sram_mem[91394] = 16'b0000000000000000;
	sram_mem[91395] = 16'b0000000000000000;
	sram_mem[91396] = 16'b0000000000000000;
	sram_mem[91397] = 16'b0000000000000000;
	sram_mem[91398] = 16'b0000000000000000;
	sram_mem[91399] = 16'b0000000000000000;
	sram_mem[91400] = 16'b0000000000000000;
	sram_mem[91401] = 16'b0000000000000000;
	sram_mem[91402] = 16'b0000000000000000;
	sram_mem[91403] = 16'b0000000000000000;
	sram_mem[91404] = 16'b0000000000000000;
	sram_mem[91405] = 16'b0000000000000000;
	sram_mem[91406] = 16'b0000000000000000;
	sram_mem[91407] = 16'b0000000000000000;
	sram_mem[91408] = 16'b0000000000000000;
	sram_mem[91409] = 16'b0000000000000000;
	sram_mem[91410] = 16'b0000000000000000;
	sram_mem[91411] = 16'b0000000000000000;
	sram_mem[91412] = 16'b0000000000000000;
	sram_mem[91413] = 16'b0000000000000000;
	sram_mem[91414] = 16'b0000000000000000;
	sram_mem[91415] = 16'b0000000000000000;
	sram_mem[91416] = 16'b0000000000000000;
	sram_mem[91417] = 16'b0000000000000000;
	sram_mem[91418] = 16'b0000000000000000;
	sram_mem[91419] = 16'b0000000000000000;
	sram_mem[91420] = 16'b0000000000000000;
	sram_mem[91421] = 16'b0000000000000000;
	sram_mem[91422] = 16'b0000000000000000;
	sram_mem[91423] = 16'b0000000000000000;
	sram_mem[91424] = 16'b0000000000000000;
	sram_mem[91425] = 16'b0000000000000000;
	sram_mem[91426] = 16'b0000000000000000;
	sram_mem[91427] = 16'b0000000000000000;
	sram_mem[91428] = 16'b0000000000000000;
	sram_mem[91429] = 16'b0000000000000000;
	sram_mem[91430] = 16'b0000000000000000;
	sram_mem[91431] = 16'b0000000000000000;
	sram_mem[91432] = 16'b0000000000000000;
	sram_mem[91433] = 16'b0000000000000000;
	sram_mem[91434] = 16'b0000000000000000;
	sram_mem[91435] = 16'b0000000000000000;
	sram_mem[91436] = 16'b0000000000000000;
	sram_mem[91437] = 16'b0000000000000000;
	sram_mem[91438] = 16'b0000000000000000;
	sram_mem[91439] = 16'b0000000000000000;
	sram_mem[91440] = 16'b0000000000000000;
	sram_mem[91441] = 16'b0000000000000000;
	sram_mem[91442] = 16'b0000000000000000;
	sram_mem[91443] = 16'b0000000000000000;
	sram_mem[91444] = 16'b0000000000000000;
	sram_mem[91445] = 16'b0000000000000000;
	sram_mem[91446] = 16'b0000000000000000;
	sram_mem[91447] = 16'b0000000000000000;
	sram_mem[91448] = 16'b0000000000000000;
	sram_mem[91449] = 16'b0000000000000000;
	sram_mem[91450] = 16'b0000000000000000;
	sram_mem[91451] = 16'b0000000000000000;
	sram_mem[91452] = 16'b0000000000000000;
	sram_mem[91453] = 16'b0000000000000000;
	sram_mem[91454] = 16'b0000000000000000;
	sram_mem[91455] = 16'b0000000000000000;
	sram_mem[91456] = 16'b0000000000000000;
	sram_mem[91457] = 16'b0000000000000000;
	sram_mem[91458] = 16'b0000000000000000;
	sram_mem[91459] = 16'b0000000000000000;
	sram_mem[91460] = 16'b0000000000000000;
	sram_mem[91461] = 16'b0000000000000000;
	sram_mem[91462] = 16'b0000000000000000;
	sram_mem[91463] = 16'b0000000000000000;
	sram_mem[91464] = 16'b0000000000000000;
	sram_mem[91465] = 16'b0000000000000000;
	sram_mem[91466] = 16'b0000000000000000;
	sram_mem[91467] = 16'b0000000000000000;
	sram_mem[91468] = 16'b0000000000000000;
	sram_mem[91469] = 16'b0000000000000000;
	sram_mem[91470] = 16'b0000000000000000;
	sram_mem[91471] = 16'b0000000000000000;
	sram_mem[91472] = 16'b0000000000000000;
	sram_mem[91473] = 16'b0000000000000000;
	sram_mem[91474] = 16'b0000000000000000;
	sram_mem[91475] = 16'b0000000000000000;
	sram_mem[91476] = 16'b0000000000000000;
	sram_mem[91477] = 16'b0000000000000000;
	sram_mem[91478] = 16'b0000000000000000;
	sram_mem[91479] = 16'b0000000000000000;
	sram_mem[91480] = 16'b0000000000000000;
	sram_mem[91481] = 16'b0000000000000000;
	sram_mem[91482] = 16'b0000000000000000;
	sram_mem[91483] = 16'b0000000000000000;
	sram_mem[91484] = 16'b0000000000000000;
	sram_mem[91485] = 16'b0000000000000000;
	sram_mem[91486] = 16'b0000000000000000;
	sram_mem[91487] = 16'b0000000000000000;
	sram_mem[91488] = 16'b0000000000000000;
	sram_mem[91489] = 16'b0000000000000000;
	sram_mem[91490] = 16'b0000000000000000;
	sram_mem[91491] = 16'b0000000000000000;
	sram_mem[91492] = 16'b0000000000000000;
	sram_mem[91493] = 16'b0000000000000000;
	sram_mem[91494] = 16'b0000000000000000;
	sram_mem[91495] = 16'b0000000000000000;
	sram_mem[91496] = 16'b0000000000000000;
	sram_mem[91497] = 16'b0000000000000000;
	sram_mem[91498] = 16'b0000000000000000;
	sram_mem[91499] = 16'b0000000000000000;
	sram_mem[91500] = 16'b0000000000000000;
	sram_mem[91501] = 16'b0000000000000000;
	sram_mem[91502] = 16'b0000000000000000;
	sram_mem[91503] = 16'b0000000000000000;
	sram_mem[91504] = 16'b0000000000000000;
	sram_mem[91505] = 16'b0000000000000000;
	sram_mem[91506] = 16'b0000000000000000;
	sram_mem[91507] = 16'b0000000000000000;
	sram_mem[91508] = 16'b0000000000000000;
	sram_mem[91509] = 16'b0000000000000000;
	sram_mem[91510] = 16'b0000000000000000;
	sram_mem[91511] = 16'b0000000000000000;
	sram_mem[91512] = 16'b0000000000000000;
	sram_mem[91513] = 16'b0000000000000000;
	sram_mem[91514] = 16'b0000000000000000;
	sram_mem[91515] = 16'b0000000000000000;
	sram_mem[91516] = 16'b0000000000000000;
	sram_mem[91517] = 16'b0000000000000000;
	sram_mem[91518] = 16'b0000000000000000;
	sram_mem[91519] = 16'b0000000000000000;
	sram_mem[91520] = 16'b0000000000000000;
	sram_mem[91521] = 16'b0000000000000000;
	sram_mem[91522] = 16'b0000000000000000;
	sram_mem[91523] = 16'b0000000000000000;
	sram_mem[91524] = 16'b0000000000000000;
	sram_mem[91525] = 16'b0000000000000000;
	sram_mem[91526] = 16'b0000000000000000;
	sram_mem[91527] = 16'b0000000000000000;
	sram_mem[91528] = 16'b0000000000000000;
	sram_mem[91529] = 16'b0000000000000000;
	sram_mem[91530] = 16'b0000000000000000;
	sram_mem[91531] = 16'b0000000000000000;
	sram_mem[91532] = 16'b0000000000000000;
	sram_mem[91533] = 16'b0000000000000000;
	sram_mem[91534] = 16'b0000000000000000;
	sram_mem[91535] = 16'b0000000000000000;
	sram_mem[91536] = 16'b0000000000000000;
	sram_mem[91537] = 16'b0000000000000000;
	sram_mem[91538] = 16'b0000000000000000;
	sram_mem[91539] = 16'b0000000000000000;
	sram_mem[91540] = 16'b0000000000000000;
	sram_mem[91541] = 16'b0000000000000000;
	sram_mem[91542] = 16'b0000000000000000;
	sram_mem[91543] = 16'b0000000000000000;
	sram_mem[91544] = 16'b0000000000000000;
	sram_mem[91545] = 16'b0000000000000000;
	sram_mem[91546] = 16'b0000000000000000;
	sram_mem[91547] = 16'b0000000000000000;
	sram_mem[91548] = 16'b0000000000000000;
	sram_mem[91549] = 16'b0000000000000000;
	sram_mem[91550] = 16'b0000000000000000;
	sram_mem[91551] = 16'b0000000000000000;
	sram_mem[91552] = 16'b0000000000000000;
	sram_mem[91553] = 16'b0000000000000000;
	sram_mem[91554] = 16'b0000000000000000;
	sram_mem[91555] = 16'b0000000000000000;
	sram_mem[91556] = 16'b0000000000000000;
	sram_mem[91557] = 16'b0000000000000000;
	sram_mem[91558] = 16'b0000000000000000;
	sram_mem[91559] = 16'b0000000000000000;
	sram_mem[91560] = 16'b0000000000000000;
	sram_mem[91561] = 16'b0000000000000000;
	sram_mem[91562] = 16'b0000000000000000;
	sram_mem[91563] = 16'b0000000000000000;
	sram_mem[91564] = 16'b0000000000000000;
	sram_mem[91565] = 16'b0000000000000000;
	sram_mem[91566] = 16'b0000000000000000;
	sram_mem[91567] = 16'b0000000000000000;
	sram_mem[91568] = 16'b0000000000000000;
	sram_mem[91569] = 16'b0000000000000000;
	sram_mem[91570] = 16'b0000000000000000;
	sram_mem[91571] = 16'b0000000000000000;
	sram_mem[91572] = 16'b0000000000000000;
	sram_mem[91573] = 16'b0000000000000000;
	sram_mem[91574] = 16'b0000000000000000;
	sram_mem[91575] = 16'b0000000000000000;
	sram_mem[91576] = 16'b0000000000000000;
	sram_mem[91577] = 16'b0000000000000000;
	sram_mem[91578] = 16'b0000000000000000;
	sram_mem[91579] = 16'b0000000000000000;
	sram_mem[91580] = 16'b0000000000000000;
	sram_mem[91581] = 16'b0000000000000000;
	sram_mem[91582] = 16'b0000000000000000;
	sram_mem[91583] = 16'b0000000000000000;
	sram_mem[91584] = 16'b0000000000000000;
	sram_mem[91585] = 16'b0000000000000000;
	sram_mem[91586] = 16'b0000000000000000;
	sram_mem[91587] = 16'b0000000000000000;
	sram_mem[91588] = 16'b0000000000000000;
	sram_mem[91589] = 16'b0000000000000000;
	sram_mem[91590] = 16'b0000000000000000;
	sram_mem[91591] = 16'b0000000000000000;
	sram_mem[91592] = 16'b0000000000000000;
	sram_mem[91593] = 16'b0000000000000000;
	sram_mem[91594] = 16'b0000000000000000;
	sram_mem[91595] = 16'b0000000000000000;
	sram_mem[91596] = 16'b0000000000000000;
	sram_mem[91597] = 16'b0000000000000000;
	sram_mem[91598] = 16'b0000000000000000;
	sram_mem[91599] = 16'b0000000000000000;
	sram_mem[91600] = 16'b0000000000000000;
	sram_mem[91601] = 16'b0000000000000000;
	sram_mem[91602] = 16'b0000000000000000;
	sram_mem[91603] = 16'b0000000000000000;
	sram_mem[91604] = 16'b0000000000000000;
	sram_mem[91605] = 16'b0000000000000000;
	sram_mem[91606] = 16'b0000000000000000;
	sram_mem[91607] = 16'b0000000000000000;
	sram_mem[91608] = 16'b0000000000000000;
	sram_mem[91609] = 16'b0000000000000000;
	sram_mem[91610] = 16'b0000000000000000;
	sram_mem[91611] = 16'b0000000000000000;
	sram_mem[91612] = 16'b0000000000000000;
	sram_mem[91613] = 16'b0000000000000000;
	sram_mem[91614] = 16'b0000000000000000;
	sram_mem[91615] = 16'b0000000000000000;
	sram_mem[91616] = 16'b0000000000000000;
	sram_mem[91617] = 16'b0000000000000000;
	sram_mem[91618] = 16'b0000000000000000;
	sram_mem[91619] = 16'b0000000000000000;
	sram_mem[91620] = 16'b0000000000000000;
	sram_mem[91621] = 16'b0000000000000000;
	sram_mem[91622] = 16'b0000000000000000;
	sram_mem[91623] = 16'b0000000000000000;
	sram_mem[91624] = 16'b0000000000000000;
	sram_mem[91625] = 16'b0000000000000000;
	sram_mem[91626] = 16'b0000000000000000;
	sram_mem[91627] = 16'b0000000000000000;
	sram_mem[91628] = 16'b0000000000000000;
	sram_mem[91629] = 16'b0000000000000000;
	sram_mem[91630] = 16'b0000000000000000;
	sram_mem[91631] = 16'b0000000000000000;
	sram_mem[91632] = 16'b0000000000000000;
	sram_mem[91633] = 16'b0000000000000000;
	sram_mem[91634] = 16'b0000000000000000;
	sram_mem[91635] = 16'b0000000000000000;
	sram_mem[91636] = 16'b0000000000000000;
	sram_mem[91637] = 16'b0000000000000000;
	sram_mem[91638] = 16'b0000000000000000;
	sram_mem[91639] = 16'b0000000000000000;
	sram_mem[91640] = 16'b0000000000000000;
	sram_mem[91641] = 16'b0000000000000000;
	sram_mem[91642] = 16'b0000000000000000;
	sram_mem[91643] = 16'b0000000000000000;
	sram_mem[91644] = 16'b0000000000000000;
	sram_mem[91645] = 16'b0000000000000000;
	sram_mem[91646] = 16'b0000000000000000;
	sram_mem[91647] = 16'b0000000000000000;
	sram_mem[91648] = 16'b0000000000000000;
	sram_mem[91649] = 16'b0000000000000000;
	sram_mem[91650] = 16'b0000000000000000;
	sram_mem[91651] = 16'b0000000000000000;
	sram_mem[91652] = 16'b0000000000000000;
	sram_mem[91653] = 16'b0000000000000000;
	sram_mem[91654] = 16'b0000000000000000;
	sram_mem[91655] = 16'b0000000000000000;
	sram_mem[91656] = 16'b0000000000000000;
	sram_mem[91657] = 16'b0000000000000000;
	sram_mem[91658] = 16'b0000000000000000;
	sram_mem[91659] = 16'b0000000000000000;
	sram_mem[91660] = 16'b0000000000000000;
	sram_mem[91661] = 16'b0000000000000000;
	sram_mem[91662] = 16'b0000000000000000;
	sram_mem[91663] = 16'b0000000000000000;
	sram_mem[91664] = 16'b0000000000000000;
	sram_mem[91665] = 16'b0000000000000000;
	sram_mem[91666] = 16'b0000000000000000;
	sram_mem[91667] = 16'b0000000000000000;
	sram_mem[91668] = 16'b0000000000000000;
	sram_mem[91669] = 16'b0000000000000000;
	sram_mem[91670] = 16'b0000000000000000;
	sram_mem[91671] = 16'b0000000000000000;
	sram_mem[91672] = 16'b0000000000000000;
	sram_mem[91673] = 16'b0000000000000000;
	sram_mem[91674] = 16'b0000000000000000;
	sram_mem[91675] = 16'b0000000000000000;
	sram_mem[91676] = 16'b0000000000000000;
	sram_mem[91677] = 16'b0000000000000000;
	sram_mem[91678] = 16'b0000000000000000;
	sram_mem[91679] = 16'b0000000000000000;
	sram_mem[91680] = 16'b0000000000000000;
	sram_mem[91681] = 16'b0000000000000000;
	sram_mem[91682] = 16'b0000000000000000;
	sram_mem[91683] = 16'b0000000000000000;
	sram_mem[91684] = 16'b0000000000000000;
	sram_mem[91685] = 16'b0000000000000000;
	sram_mem[91686] = 16'b0000000000000000;
	sram_mem[91687] = 16'b0000000000000000;
	sram_mem[91688] = 16'b0000000000000000;
	sram_mem[91689] = 16'b0000000000000000;
	sram_mem[91690] = 16'b0000000000000000;
	sram_mem[91691] = 16'b0000000000000000;
	sram_mem[91692] = 16'b0000000000000000;
	sram_mem[91693] = 16'b0000000000000000;
	sram_mem[91694] = 16'b0000000000000000;
	sram_mem[91695] = 16'b0000000000000000;
	sram_mem[91696] = 16'b0000000000000000;
	sram_mem[91697] = 16'b0000000000000000;
	sram_mem[91698] = 16'b0000000000000000;
	sram_mem[91699] = 16'b0000000000000000;
	sram_mem[91700] = 16'b0000000000000000;
	sram_mem[91701] = 16'b0000000000000000;
	sram_mem[91702] = 16'b0000000000000000;
	sram_mem[91703] = 16'b0000000000000000;
	sram_mem[91704] = 16'b0000000000000000;
	sram_mem[91705] = 16'b0000000000000000;
	sram_mem[91706] = 16'b0000000000000000;
	sram_mem[91707] = 16'b0000000000000000;
	sram_mem[91708] = 16'b0000000000000000;
	sram_mem[91709] = 16'b0000000000000000;
	sram_mem[91710] = 16'b0000000000000000;
	sram_mem[91711] = 16'b0000000000000000;
	sram_mem[91712] = 16'b0000000000000000;
	sram_mem[91713] = 16'b0000000000000000;
	sram_mem[91714] = 16'b0000000000000000;
	sram_mem[91715] = 16'b0000000000000000;
	sram_mem[91716] = 16'b0000000000000000;
	sram_mem[91717] = 16'b0000000000000000;
	sram_mem[91718] = 16'b0000000000000000;
	sram_mem[91719] = 16'b0000000000000000;
	sram_mem[91720] = 16'b0000000000000000;
	sram_mem[91721] = 16'b0000000000000000;
	sram_mem[91722] = 16'b0000000000000000;
	sram_mem[91723] = 16'b0000000000000000;
	sram_mem[91724] = 16'b0000000000000000;
	sram_mem[91725] = 16'b0000000000000000;
	sram_mem[91726] = 16'b0000000000000000;
	sram_mem[91727] = 16'b0000000000000000;
	sram_mem[91728] = 16'b0000000000000000;
	sram_mem[91729] = 16'b0000000000000000;
	sram_mem[91730] = 16'b0000000000000000;
	sram_mem[91731] = 16'b0000000000000000;
	sram_mem[91732] = 16'b0000000000000000;
	sram_mem[91733] = 16'b0000000000000000;
	sram_mem[91734] = 16'b0000000000000000;
	sram_mem[91735] = 16'b0000000000000000;
	sram_mem[91736] = 16'b0000000000000000;
	sram_mem[91737] = 16'b0000000000000000;
	sram_mem[91738] = 16'b0000000000000000;
	sram_mem[91739] = 16'b0000000000000000;
	sram_mem[91740] = 16'b0000000000000000;
	sram_mem[91741] = 16'b0000000000000000;
	sram_mem[91742] = 16'b0000000000000000;
	sram_mem[91743] = 16'b0000000000000000;
	sram_mem[91744] = 16'b0000000000000000;
	sram_mem[91745] = 16'b0000000000000000;
	sram_mem[91746] = 16'b0000000000000000;
	sram_mem[91747] = 16'b0000000000000000;
	sram_mem[91748] = 16'b0000000000000000;
	sram_mem[91749] = 16'b0000000000000000;
	sram_mem[91750] = 16'b0000000000000000;
	sram_mem[91751] = 16'b0000000000000000;
	sram_mem[91752] = 16'b0000000000000000;
	sram_mem[91753] = 16'b0000000000000000;
	sram_mem[91754] = 16'b0000000000000000;
	sram_mem[91755] = 16'b0000000000000000;
	sram_mem[91756] = 16'b0000000000000000;
	sram_mem[91757] = 16'b0000000000000000;
	sram_mem[91758] = 16'b0000000000000000;
	sram_mem[91759] = 16'b0000000000000000;
	sram_mem[91760] = 16'b0000000000000000;
	sram_mem[91761] = 16'b0000000000000000;
	sram_mem[91762] = 16'b0000000000000000;
	sram_mem[91763] = 16'b0000000000000000;
	sram_mem[91764] = 16'b0000000000000000;
	sram_mem[91765] = 16'b0000000000000000;
	sram_mem[91766] = 16'b0000000000000000;
	sram_mem[91767] = 16'b0000000000000000;
	sram_mem[91768] = 16'b0000000000000000;
	sram_mem[91769] = 16'b0000000000000000;
	sram_mem[91770] = 16'b0000000000000000;
	sram_mem[91771] = 16'b0000000000000000;
	sram_mem[91772] = 16'b0000000000000000;
	sram_mem[91773] = 16'b0000000000000000;
	sram_mem[91774] = 16'b0000000000000000;
	sram_mem[91775] = 16'b0000000000000000;
	sram_mem[91776] = 16'b0000000000000000;
	sram_mem[91777] = 16'b0000000000000000;
	sram_mem[91778] = 16'b0000000000000000;
	sram_mem[91779] = 16'b0000000000000000;
	sram_mem[91780] = 16'b0000000000000000;
	sram_mem[91781] = 16'b0000000000000000;
	sram_mem[91782] = 16'b0000000000000000;
	sram_mem[91783] = 16'b0000000000000000;
	sram_mem[91784] = 16'b0000000000000000;
	sram_mem[91785] = 16'b0000000000000000;
	sram_mem[91786] = 16'b0000000000000000;
	sram_mem[91787] = 16'b0000000000000000;
	sram_mem[91788] = 16'b0000000000000000;
	sram_mem[91789] = 16'b0000000000000000;
	sram_mem[91790] = 16'b0000000000000000;
	sram_mem[91791] = 16'b0000000000000000;
	sram_mem[91792] = 16'b0000000000000000;
	sram_mem[91793] = 16'b0000000000000000;
	sram_mem[91794] = 16'b0000000000000000;
	sram_mem[91795] = 16'b0000000000000000;
	sram_mem[91796] = 16'b0000000000000000;
	sram_mem[91797] = 16'b0000000000000000;
	sram_mem[91798] = 16'b0000000000000000;
	sram_mem[91799] = 16'b0000000000000000;
	sram_mem[91800] = 16'b0000000000000000;
	sram_mem[91801] = 16'b0000000000000000;
	sram_mem[91802] = 16'b0000000000000000;
	sram_mem[91803] = 16'b0000000000000000;
	sram_mem[91804] = 16'b0000000000000000;
	sram_mem[91805] = 16'b0000000000000000;
	sram_mem[91806] = 16'b0000000000000000;
	sram_mem[91807] = 16'b0000000000000000;
	sram_mem[91808] = 16'b0000000000000000;
	sram_mem[91809] = 16'b0000000000000000;
	sram_mem[91810] = 16'b0000000000000000;
	sram_mem[91811] = 16'b0000000000000000;
	sram_mem[91812] = 16'b0000000000000000;
	sram_mem[91813] = 16'b0000000000000000;
	sram_mem[91814] = 16'b0000000000000000;
	sram_mem[91815] = 16'b0000000000000000;
	sram_mem[91816] = 16'b0000000000000000;
	sram_mem[91817] = 16'b0000000000000000;
	sram_mem[91818] = 16'b0000000000000000;
	sram_mem[91819] = 16'b0000000000000000;
	sram_mem[91820] = 16'b0000000000000000;
	sram_mem[91821] = 16'b0000000000000000;
	sram_mem[91822] = 16'b0000000000000000;
	sram_mem[91823] = 16'b0000000000000000;
	sram_mem[91824] = 16'b0000000000000000;
	sram_mem[91825] = 16'b0000000000000000;
	sram_mem[91826] = 16'b0000000000000000;
	sram_mem[91827] = 16'b0000000000000000;
	sram_mem[91828] = 16'b0000000000000000;
	sram_mem[91829] = 16'b0000000000000000;
	sram_mem[91830] = 16'b0000000000000000;
	sram_mem[91831] = 16'b0000000000000000;
	sram_mem[91832] = 16'b0000000000000000;
	sram_mem[91833] = 16'b0000000000000000;
	sram_mem[91834] = 16'b0000000000000000;
	sram_mem[91835] = 16'b0000000000000000;
	sram_mem[91836] = 16'b0000000000000000;
	sram_mem[91837] = 16'b0000000000000000;
	sram_mem[91838] = 16'b0000000000000000;
	sram_mem[91839] = 16'b0000000000000000;
	sram_mem[91840] = 16'b0000000000000000;
	sram_mem[91841] = 16'b0000000000000000;
	sram_mem[91842] = 16'b0000000000000000;
	sram_mem[91843] = 16'b0000000000000000;
	sram_mem[91844] = 16'b0000000000000000;
	sram_mem[91845] = 16'b0000000000000000;
	sram_mem[91846] = 16'b0000000000000000;
	sram_mem[91847] = 16'b0000000000000000;
	sram_mem[91848] = 16'b0000000000000000;
	sram_mem[91849] = 16'b0000000000000000;
	sram_mem[91850] = 16'b0000000000000000;
	sram_mem[91851] = 16'b0000000000000000;
	sram_mem[91852] = 16'b0000000000000000;
	sram_mem[91853] = 16'b0000000000000000;
	sram_mem[91854] = 16'b0000000000000000;
	sram_mem[91855] = 16'b0000000000000000;
	sram_mem[91856] = 16'b0000000000000000;
	sram_mem[91857] = 16'b0000000000000000;
	sram_mem[91858] = 16'b0000000000000000;
	sram_mem[91859] = 16'b0000000000000000;
	sram_mem[91860] = 16'b0000000000000000;
	sram_mem[91861] = 16'b0000000000000000;
	sram_mem[91862] = 16'b0000000000000000;
	sram_mem[91863] = 16'b0000000000000000;
	sram_mem[91864] = 16'b0000000000000000;
	sram_mem[91865] = 16'b0000000000000000;
	sram_mem[91866] = 16'b0000000000000000;
	sram_mem[91867] = 16'b0000000000000000;
	sram_mem[91868] = 16'b0000000000000000;
	sram_mem[91869] = 16'b0000000000000000;
	sram_mem[91870] = 16'b0000000000000000;
	sram_mem[91871] = 16'b0000000000000000;
	sram_mem[91872] = 16'b0000000000000000;
	sram_mem[91873] = 16'b0000000000000000;
	sram_mem[91874] = 16'b0000000000000000;
	sram_mem[91875] = 16'b0000000000000000;
	sram_mem[91876] = 16'b0000000000000000;
	sram_mem[91877] = 16'b0000000000000000;
	sram_mem[91878] = 16'b0000000000000000;
	sram_mem[91879] = 16'b0000000000000000;
	sram_mem[91880] = 16'b0000000000000000;
	sram_mem[91881] = 16'b0000000000000000;
	sram_mem[91882] = 16'b0000000000000000;
	sram_mem[91883] = 16'b0000000000000000;
	sram_mem[91884] = 16'b0000000000000000;
	sram_mem[91885] = 16'b0000000000000000;
	sram_mem[91886] = 16'b0000000000000000;
	sram_mem[91887] = 16'b0000000000000000;
	sram_mem[91888] = 16'b0000000000000000;
	sram_mem[91889] = 16'b0000000000000000;
	sram_mem[91890] = 16'b0000000000000000;
	sram_mem[91891] = 16'b0000000000000000;
	sram_mem[91892] = 16'b0000000000000000;
	sram_mem[91893] = 16'b0000000000000000;
	sram_mem[91894] = 16'b0000000000000000;
	sram_mem[91895] = 16'b0000000000000000;
	sram_mem[91896] = 16'b0000000000000000;
	sram_mem[91897] = 16'b0000000000000000;
	sram_mem[91898] = 16'b0000000000000000;
	sram_mem[91899] = 16'b0000000000000000;
	sram_mem[91900] = 16'b0000000000000000;
	sram_mem[91901] = 16'b0000000000000000;
	sram_mem[91902] = 16'b0000000000000000;
	sram_mem[91903] = 16'b0000000000000000;
	sram_mem[91904] = 16'b0000000000000000;
	sram_mem[91905] = 16'b0000000000000000;
	sram_mem[91906] = 16'b0000000000000000;
	sram_mem[91907] = 16'b0000000000000000;
	sram_mem[91908] = 16'b0000000000000000;
	sram_mem[91909] = 16'b0000000000000000;
	sram_mem[91910] = 16'b0000000000000000;
	sram_mem[91911] = 16'b0000000000000000;
	sram_mem[91912] = 16'b0000000000000000;
	sram_mem[91913] = 16'b0000000000000000;
	sram_mem[91914] = 16'b0000000000000000;
	sram_mem[91915] = 16'b0000000000000000;
	sram_mem[91916] = 16'b0000000000000000;
	sram_mem[91917] = 16'b0000000000000000;
	sram_mem[91918] = 16'b0000000000000000;
	sram_mem[91919] = 16'b0000000000000000;
	sram_mem[91920] = 16'b0000000000000000;
	sram_mem[91921] = 16'b0000000000000000;
	sram_mem[91922] = 16'b0000000000000000;
	sram_mem[91923] = 16'b0000000000000000;
	sram_mem[91924] = 16'b0000000000000000;
	sram_mem[91925] = 16'b0000000000000000;
	sram_mem[91926] = 16'b0000000000000000;
	sram_mem[91927] = 16'b0000000000000000;
	sram_mem[91928] = 16'b0000000000000000;
	sram_mem[91929] = 16'b0000000000000000;
	sram_mem[91930] = 16'b0000000000000000;
	sram_mem[91931] = 16'b0000000000000000;
	sram_mem[91932] = 16'b0000000000000000;
	sram_mem[91933] = 16'b0000000000000000;
	sram_mem[91934] = 16'b0000000000000000;
	sram_mem[91935] = 16'b0000000000000000;
	sram_mem[91936] = 16'b0000000000000000;
	sram_mem[91937] = 16'b0000000000000000;
	sram_mem[91938] = 16'b0000000000000000;
	sram_mem[91939] = 16'b0000000000000000;
	sram_mem[91940] = 16'b0000000000000000;
	sram_mem[91941] = 16'b0000000000000000;
	sram_mem[91942] = 16'b0000000000000000;
	sram_mem[91943] = 16'b0000000000000000;
	sram_mem[91944] = 16'b0000000000000000;
	sram_mem[91945] = 16'b0000000000000000;
	sram_mem[91946] = 16'b0000000000000000;
	sram_mem[91947] = 16'b0000000000000000;
	sram_mem[91948] = 16'b0000000000000000;
	sram_mem[91949] = 16'b0000000000000000;
	sram_mem[91950] = 16'b0000000000000000;
	sram_mem[91951] = 16'b0000000000000000;
	sram_mem[91952] = 16'b0000000000000000;
	sram_mem[91953] = 16'b0000000000000000;
	sram_mem[91954] = 16'b0000000000000000;
	sram_mem[91955] = 16'b0000000000000000;
	sram_mem[91956] = 16'b0000000000000000;
	sram_mem[91957] = 16'b0000000000000000;
	sram_mem[91958] = 16'b0000000000000000;
	sram_mem[91959] = 16'b0000000000000000;
	sram_mem[91960] = 16'b0000000000000000;
	sram_mem[91961] = 16'b0000000000000000;
	sram_mem[91962] = 16'b0000000000000000;
	sram_mem[91963] = 16'b0000000000000000;
	sram_mem[91964] = 16'b0000000000000000;
	sram_mem[91965] = 16'b0000000000000000;
	sram_mem[91966] = 16'b0000000000000000;
	sram_mem[91967] = 16'b0000000000000000;
	sram_mem[91968] = 16'b0000000000000000;
	sram_mem[91969] = 16'b0000000000000000;
	sram_mem[91970] = 16'b0000000000000000;
	sram_mem[91971] = 16'b0000000000000000;
	sram_mem[91972] = 16'b0000000000000000;
	sram_mem[91973] = 16'b0000000000000000;
	sram_mem[91974] = 16'b0000000000000000;
	sram_mem[91975] = 16'b0000000000000000;
	sram_mem[91976] = 16'b0000000000000000;
	sram_mem[91977] = 16'b0000000000000000;
	sram_mem[91978] = 16'b0000000000000000;
	sram_mem[91979] = 16'b0000000000000000;
	sram_mem[91980] = 16'b0000000000000000;
	sram_mem[91981] = 16'b0000000000000000;
	sram_mem[91982] = 16'b0000000000000000;
	sram_mem[91983] = 16'b0000000000000000;
	sram_mem[91984] = 16'b0000000000000000;
	sram_mem[91985] = 16'b0000000000000000;
	sram_mem[91986] = 16'b0000000000000000;
	sram_mem[91987] = 16'b0000000000000000;
	sram_mem[91988] = 16'b0000000000000000;
	sram_mem[91989] = 16'b0000000000000000;
	sram_mem[91990] = 16'b0000000000000000;
	sram_mem[91991] = 16'b0000000000000000;
	sram_mem[91992] = 16'b0000000000000000;
	sram_mem[91993] = 16'b0000000000000000;
	sram_mem[91994] = 16'b0000000000000000;
	sram_mem[91995] = 16'b0000000000000000;
	sram_mem[91996] = 16'b0000000000000000;
	sram_mem[91997] = 16'b0000000000000000;
	sram_mem[91998] = 16'b0000000000000000;
	sram_mem[91999] = 16'b0000000000000000;
	sram_mem[92000] = 16'b0000000000000000;
	sram_mem[92001] = 16'b0000000000000000;
	sram_mem[92002] = 16'b0000000000000000;
	sram_mem[92003] = 16'b0000000000000000;
	sram_mem[92004] = 16'b0000000000000000;
	sram_mem[92005] = 16'b0000000000000000;
	sram_mem[92006] = 16'b0000000000000000;
	sram_mem[92007] = 16'b0000000000000000;
	sram_mem[92008] = 16'b0000000000000000;
	sram_mem[92009] = 16'b0000000000000000;
	sram_mem[92010] = 16'b0000000000000000;
	sram_mem[92011] = 16'b0000000000000000;
	sram_mem[92012] = 16'b0000000000000000;
	sram_mem[92013] = 16'b0000000000000000;
	sram_mem[92014] = 16'b0000000000000000;
	sram_mem[92015] = 16'b0000000000000000;
	sram_mem[92016] = 16'b0000000000000000;
	sram_mem[92017] = 16'b0000000000000000;
	sram_mem[92018] = 16'b0000000000000000;
	sram_mem[92019] = 16'b0000000000000000;
	sram_mem[92020] = 16'b0000000000000000;
	sram_mem[92021] = 16'b0000000000000000;
	sram_mem[92022] = 16'b0000000000000000;
	sram_mem[92023] = 16'b0000000000000000;
	sram_mem[92024] = 16'b0000000000000000;
	sram_mem[92025] = 16'b0000000000000000;
	sram_mem[92026] = 16'b0000000000000000;
	sram_mem[92027] = 16'b0000000000000000;
	sram_mem[92028] = 16'b0000000000000000;
	sram_mem[92029] = 16'b0000000000000000;
	sram_mem[92030] = 16'b0000000000000000;
	sram_mem[92031] = 16'b0000000000000000;
	sram_mem[92032] = 16'b0000000000000000;
	sram_mem[92033] = 16'b0000000000000000;
	sram_mem[92034] = 16'b0000000000000000;
	sram_mem[92035] = 16'b0000000000000000;
	sram_mem[92036] = 16'b0000000000000000;
	sram_mem[92037] = 16'b0000000000000000;
	sram_mem[92038] = 16'b0000000000000000;
	sram_mem[92039] = 16'b0000000000000000;
	sram_mem[92040] = 16'b0000000000000000;
	sram_mem[92041] = 16'b0000000000000000;
	sram_mem[92042] = 16'b0000000000000000;
	sram_mem[92043] = 16'b0000000000000000;
	sram_mem[92044] = 16'b0000000000000000;
	sram_mem[92045] = 16'b0000000000000000;
	sram_mem[92046] = 16'b0000000000000000;
	sram_mem[92047] = 16'b0000000000000000;
	sram_mem[92048] = 16'b0000000000000000;
	sram_mem[92049] = 16'b0000000000000000;
	sram_mem[92050] = 16'b0000000000000000;
	sram_mem[92051] = 16'b0000000000000000;
	sram_mem[92052] = 16'b0000000000000000;
	sram_mem[92053] = 16'b0000000000000000;
	sram_mem[92054] = 16'b0000000000000000;
	sram_mem[92055] = 16'b0000000000000000;
	sram_mem[92056] = 16'b0000000000000000;
	sram_mem[92057] = 16'b0000000000000000;
	sram_mem[92058] = 16'b0000000000000000;
	sram_mem[92059] = 16'b0000000000000000;
	sram_mem[92060] = 16'b0000000000000000;
	sram_mem[92061] = 16'b0000000000000000;
	sram_mem[92062] = 16'b0000000000000000;
	sram_mem[92063] = 16'b0000000000000000;
	sram_mem[92064] = 16'b0000000000000000;
	sram_mem[92065] = 16'b0000000000000000;
	sram_mem[92066] = 16'b0000000000000000;
	sram_mem[92067] = 16'b0000000000000000;
	sram_mem[92068] = 16'b0000000000000000;
	sram_mem[92069] = 16'b0000000000000000;
	sram_mem[92070] = 16'b0000000000000000;
	sram_mem[92071] = 16'b0000000000000000;
	sram_mem[92072] = 16'b0000000000000000;
	sram_mem[92073] = 16'b0000000000000000;
	sram_mem[92074] = 16'b0000000000000000;
	sram_mem[92075] = 16'b0000000000000000;
	sram_mem[92076] = 16'b0000000000000000;
	sram_mem[92077] = 16'b0000000000000000;
	sram_mem[92078] = 16'b0000000000000000;
	sram_mem[92079] = 16'b0000000000000000;
	sram_mem[92080] = 16'b0000000000000000;
	sram_mem[92081] = 16'b0000000000000000;
	sram_mem[92082] = 16'b0000000000000000;
	sram_mem[92083] = 16'b0000000000000000;
	sram_mem[92084] = 16'b0000000000000000;
	sram_mem[92085] = 16'b0000000000000000;
	sram_mem[92086] = 16'b0000000000000000;
	sram_mem[92087] = 16'b0000000000000000;
	sram_mem[92088] = 16'b0000000000000000;
	sram_mem[92089] = 16'b0000000000000000;
	sram_mem[92090] = 16'b0000000000000000;
	sram_mem[92091] = 16'b0000000000000000;
	sram_mem[92092] = 16'b0000000000000000;
	sram_mem[92093] = 16'b0000000000000000;
	sram_mem[92094] = 16'b0000000000000000;
	sram_mem[92095] = 16'b0000000000000000;
	sram_mem[92096] = 16'b0000000000000000;
	sram_mem[92097] = 16'b0000000000000000;
	sram_mem[92098] = 16'b0000000000000000;
	sram_mem[92099] = 16'b0000000000000000;
	sram_mem[92100] = 16'b0000000000000000;
	sram_mem[92101] = 16'b0000000000000000;
	sram_mem[92102] = 16'b0000000000000000;
	sram_mem[92103] = 16'b0000000000000000;
	sram_mem[92104] = 16'b0000000000000000;
	sram_mem[92105] = 16'b0000000000000000;
	sram_mem[92106] = 16'b0000000000000000;
	sram_mem[92107] = 16'b0000000000000000;
	sram_mem[92108] = 16'b0000000000000000;
	sram_mem[92109] = 16'b0000000000000000;
	sram_mem[92110] = 16'b0000000000000000;
	sram_mem[92111] = 16'b0000000000000000;
	sram_mem[92112] = 16'b0000000000000000;
	sram_mem[92113] = 16'b0000000000000000;
	sram_mem[92114] = 16'b0000000000000000;
	sram_mem[92115] = 16'b0000000000000000;
	sram_mem[92116] = 16'b0000000000000000;
	sram_mem[92117] = 16'b0000000000000000;
	sram_mem[92118] = 16'b0000000000000000;
	sram_mem[92119] = 16'b0000000000000000;
	sram_mem[92120] = 16'b0000000000000000;
	sram_mem[92121] = 16'b0000000000000000;
	sram_mem[92122] = 16'b0000000000000000;
	sram_mem[92123] = 16'b0000000000000000;
	sram_mem[92124] = 16'b0000000000000000;
	sram_mem[92125] = 16'b0000000000000000;
	sram_mem[92126] = 16'b0000000000000000;
	sram_mem[92127] = 16'b0000000000000000;
	sram_mem[92128] = 16'b0000000000000000;
	sram_mem[92129] = 16'b0000000000000000;
	sram_mem[92130] = 16'b0000000000000000;
	sram_mem[92131] = 16'b0000000000000000;
	sram_mem[92132] = 16'b0000000000000000;
	sram_mem[92133] = 16'b0000000000000000;
	sram_mem[92134] = 16'b0000000000000000;
	sram_mem[92135] = 16'b0000000000000000;
	sram_mem[92136] = 16'b0000000000000000;
	sram_mem[92137] = 16'b0000000000000000;
	sram_mem[92138] = 16'b0000000000000000;
	sram_mem[92139] = 16'b0000000000000000;
	sram_mem[92140] = 16'b0000000000000000;
	sram_mem[92141] = 16'b0000000000000000;
	sram_mem[92142] = 16'b0000000000000000;
	sram_mem[92143] = 16'b0000000000000000;
	sram_mem[92144] = 16'b0000000000000000;
	sram_mem[92145] = 16'b0000000000000000;
	sram_mem[92146] = 16'b0000000000000000;
	sram_mem[92147] = 16'b0000000000000000;
	sram_mem[92148] = 16'b0000000000000000;
	sram_mem[92149] = 16'b0000000000000000;
	sram_mem[92150] = 16'b0000000000000000;
	sram_mem[92151] = 16'b0000000000000000;
	sram_mem[92152] = 16'b0000000000000000;
	sram_mem[92153] = 16'b0000000000000000;
	sram_mem[92154] = 16'b0000000000000000;
	sram_mem[92155] = 16'b0000000000000000;
	sram_mem[92156] = 16'b0000000000000000;
	sram_mem[92157] = 16'b0000000000000000;
	sram_mem[92158] = 16'b0000000000000000;
	sram_mem[92159] = 16'b0000000000000000;
	sram_mem[92160] = 16'b0000000000000000;
	sram_mem[92161] = 16'b0000000000000000;
	sram_mem[92162] = 16'b0000000000000000;
	sram_mem[92163] = 16'b0000000000000000;
	sram_mem[92164] = 16'b0000000000000000;
	sram_mem[92165] = 16'b0000000000000000;
	sram_mem[92166] = 16'b0000000000000000;
	sram_mem[92167] = 16'b0000000000000000;
	sram_mem[92168] = 16'b0000000000000000;
	sram_mem[92169] = 16'b0000000000000000;
	sram_mem[92170] = 16'b0000000000000000;
	sram_mem[92171] = 16'b0000000000000000;
	sram_mem[92172] = 16'b0000000000000000;
	sram_mem[92173] = 16'b0000000000000000;
	sram_mem[92174] = 16'b0000000000000000;
	sram_mem[92175] = 16'b0000000000000000;
	sram_mem[92176] = 16'b0000000000000000;
	sram_mem[92177] = 16'b0000000000000000;
	sram_mem[92178] = 16'b0000000000000000;
	sram_mem[92179] = 16'b0000000000000000;
	sram_mem[92180] = 16'b0000000000000000;
	sram_mem[92181] = 16'b0000000000000000;
	sram_mem[92182] = 16'b0000000000000000;
	sram_mem[92183] = 16'b0000000000000000;
	sram_mem[92184] = 16'b0000000000000000;
	sram_mem[92185] = 16'b0000000000000000;
	sram_mem[92186] = 16'b0000000000000000;
	sram_mem[92187] = 16'b0000000000000000;
	sram_mem[92188] = 16'b0000000000000000;
	sram_mem[92189] = 16'b0000000000000000;
	sram_mem[92190] = 16'b0000000000000000;
	sram_mem[92191] = 16'b0000000000000000;
	sram_mem[92192] = 16'b0000000000000000;
	sram_mem[92193] = 16'b0000000000000000;
	sram_mem[92194] = 16'b0000000000000000;
	sram_mem[92195] = 16'b0000000000000000;
	sram_mem[92196] = 16'b0000000000000000;
	sram_mem[92197] = 16'b0000000000000000;
	sram_mem[92198] = 16'b0000000000000000;
	sram_mem[92199] = 16'b0000000000000000;
	sram_mem[92200] = 16'b0000000000000000;
	sram_mem[92201] = 16'b0000000000000000;
	sram_mem[92202] = 16'b0000000000000000;
	sram_mem[92203] = 16'b0000000000000000;
	sram_mem[92204] = 16'b0000000000000000;
	sram_mem[92205] = 16'b0000000000000000;
	sram_mem[92206] = 16'b0000000000000000;
	sram_mem[92207] = 16'b0000000000000000;
	sram_mem[92208] = 16'b0000000000000000;
	sram_mem[92209] = 16'b0000000000000000;
	sram_mem[92210] = 16'b0000000000000000;
	sram_mem[92211] = 16'b0000000000000000;
	sram_mem[92212] = 16'b0000000000000000;
	sram_mem[92213] = 16'b0000000000000000;
	sram_mem[92214] = 16'b0000000000000000;
	sram_mem[92215] = 16'b0000000000000000;
	sram_mem[92216] = 16'b0000000000000000;
	sram_mem[92217] = 16'b0000000000000000;
	sram_mem[92218] = 16'b0000000000000000;
	sram_mem[92219] = 16'b0000000000000000;
	sram_mem[92220] = 16'b0000000000000000;
	sram_mem[92221] = 16'b0000000000000000;
	sram_mem[92222] = 16'b0000000000000000;
	sram_mem[92223] = 16'b0000000000000000;
	sram_mem[92224] = 16'b0000000000000000;
	sram_mem[92225] = 16'b0000000000000000;
	sram_mem[92226] = 16'b0000000000000000;
	sram_mem[92227] = 16'b0000000000000000;
	sram_mem[92228] = 16'b0000000000000000;
	sram_mem[92229] = 16'b0000000000000000;
	sram_mem[92230] = 16'b0000000000000000;
	sram_mem[92231] = 16'b0000000000000000;
	sram_mem[92232] = 16'b0000000000000000;
	sram_mem[92233] = 16'b0000000000000000;
	sram_mem[92234] = 16'b0000000000000000;
	sram_mem[92235] = 16'b0000000000000000;
	sram_mem[92236] = 16'b0000000000000000;
	sram_mem[92237] = 16'b0000000000000000;
	sram_mem[92238] = 16'b0000000000000000;
	sram_mem[92239] = 16'b0000000000000000;
	sram_mem[92240] = 16'b0000000000000000;
	sram_mem[92241] = 16'b0000000000000000;
	sram_mem[92242] = 16'b0000000000000000;
	sram_mem[92243] = 16'b0000000000000000;
	sram_mem[92244] = 16'b0000000000000000;
	sram_mem[92245] = 16'b0000000000000000;
	sram_mem[92246] = 16'b0000000000000000;
	sram_mem[92247] = 16'b0000000000000000;
	sram_mem[92248] = 16'b0000000000000000;
	sram_mem[92249] = 16'b0000000000000000;
	sram_mem[92250] = 16'b0000000000000000;
	sram_mem[92251] = 16'b0000000000000000;
	sram_mem[92252] = 16'b0000000000000000;
	sram_mem[92253] = 16'b0000000000000000;
	sram_mem[92254] = 16'b0000000000000000;
	sram_mem[92255] = 16'b0000000000000000;
	sram_mem[92256] = 16'b0000000000000000;
	sram_mem[92257] = 16'b0000000000000000;
	sram_mem[92258] = 16'b0000000000000000;
	sram_mem[92259] = 16'b0000000000000000;
	sram_mem[92260] = 16'b0000000000000000;
	sram_mem[92261] = 16'b0000000000000000;
	sram_mem[92262] = 16'b0000000000000000;
	sram_mem[92263] = 16'b0000000000000000;
	sram_mem[92264] = 16'b0000000000000000;
	sram_mem[92265] = 16'b0000000000000000;
	sram_mem[92266] = 16'b0000000000000000;
	sram_mem[92267] = 16'b0000000000000000;
	sram_mem[92268] = 16'b0000000000000000;
	sram_mem[92269] = 16'b0000000000000000;
	sram_mem[92270] = 16'b0000000000000000;
	sram_mem[92271] = 16'b0000000000000000;
	sram_mem[92272] = 16'b0000000000000000;
	sram_mem[92273] = 16'b0000000000000000;
	sram_mem[92274] = 16'b0000000000000000;
	sram_mem[92275] = 16'b0000000000000000;
	sram_mem[92276] = 16'b0000000000000000;
	sram_mem[92277] = 16'b0000000000000000;
	sram_mem[92278] = 16'b0000000000000000;
	sram_mem[92279] = 16'b0000000000000000;
	sram_mem[92280] = 16'b0000000000000000;
	sram_mem[92281] = 16'b0000000000000000;
	sram_mem[92282] = 16'b0000000000000000;
	sram_mem[92283] = 16'b0000000000000000;
	sram_mem[92284] = 16'b0000000000000000;
	sram_mem[92285] = 16'b0000000000000000;
	sram_mem[92286] = 16'b0000000000000000;
	sram_mem[92287] = 16'b0000000000000000;
	sram_mem[92288] = 16'b0000000000000000;
	sram_mem[92289] = 16'b0000000000000000;
	sram_mem[92290] = 16'b0000000000000000;
	sram_mem[92291] = 16'b0000000000000000;
	sram_mem[92292] = 16'b0000000000000000;
	sram_mem[92293] = 16'b0000000000000000;
	sram_mem[92294] = 16'b0000000000000000;
	sram_mem[92295] = 16'b0000000000000000;
	sram_mem[92296] = 16'b0000000000000000;
	sram_mem[92297] = 16'b0000000000000000;
	sram_mem[92298] = 16'b0000000000000000;
	sram_mem[92299] = 16'b0000000000000000;
	sram_mem[92300] = 16'b0000000000000000;
	sram_mem[92301] = 16'b0000000000000000;
	sram_mem[92302] = 16'b0000000000000000;
	sram_mem[92303] = 16'b0000000000000000;
	sram_mem[92304] = 16'b0000000000000000;
	sram_mem[92305] = 16'b0000000000000000;
	sram_mem[92306] = 16'b0000000000000000;
	sram_mem[92307] = 16'b0000000000000000;
	sram_mem[92308] = 16'b0000000000000000;
	sram_mem[92309] = 16'b0000000000000000;
	sram_mem[92310] = 16'b0000000000000000;
	sram_mem[92311] = 16'b0000000000000000;
	sram_mem[92312] = 16'b0000000000000000;
	sram_mem[92313] = 16'b0000000000000000;
	sram_mem[92314] = 16'b0000000000000000;
	sram_mem[92315] = 16'b0000000000000000;
	sram_mem[92316] = 16'b0000000000000000;
	sram_mem[92317] = 16'b0000000000000000;
	sram_mem[92318] = 16'b0000000000000000;
	sram_mem[92319] = 16'b0000000000000000;
	sram_mem[92320] = 16'b0000000000000000;
	sram_mem[92321] = 16'b0000000000000000;
	sram_mem[92322] = 16'b0000000000000000;
	sram_mem[92323] = 16'b0000000000000000;
	sram_mem[92324] = 16'b0000000000000000;
	sram_mem[92325] = 16'b0000000000000000;
	sram_mem[92326] = 16'b0000000000000000;
	sram_mem[92327] = 16'b0000000000000000;
	sram_mem[92328] = 16'b0000000000000000;
	sram_mem[92329] = 16'b0000000000000000;
	sram_mem[92330] = 16'b0000000000000000;
	sram_mem[92331] = 16'b0000000000000000;
	sram_mem[92332] = 16'b0000000000000000;
	sram_mem[92333] = 16'b0000000000000000;
	sram_mem[92334] = 16'b0000000000000000;
	sram_mem[92335] = 16'b0000000000000000;
	sram_mem[92336] = 16'b0000000000000000;
	sram_mem[92337] = 16'b0000000000000000;
	sram_mem[92338] = 16'b0000000000000000;
	sram_mem[92339] = 16'b0000000000000000;
	sram_mem[92340] = 16'b0000000000000000;
	sram_mem[92341] = 16'b0000000000000000;
	sram_mem[92342] = 16'b0000000000000000;
	sram_mem[92343] = 16'b0000000000000000;
	sram_mem[92344] = 16'b0000000000000000;
	sram_mem[92345] = 16'b0000000000000000;
	sram_mem[92346] = 16'b0000000000000000;
	sram_mem[92347] = 16'b0000000000000000;
	sram_mem[92348] = 16'b0000000000000000;
	sram_mem[92349] = 16'b0000000000000000;
	sram_mem[92350] = 16'b0000000000000000;
	sram_mem[92351] = 16'b0000000000000000;
	sram_mem[92352] = 16'b0000000000000000;
	sram_mem[92353] = 16'b0000000000000000;
	sram_mem[92354] = 16'b0000000000000000;
	sram_mem[92355] = 16'b0000000000000000;
	sram_mem[92356] = 16'b0000000000000000;
	sram_mem[92357] = 16'b0000000000000000;
	sram_mem[92358] = 16'b0000000000000000;
	sram_mem[92359] = 16'b0000000000000000;
	sram_mem[92360] = 16'b0000000000000000;
	sram_mem[92361] = 16'b0000000000000000;
	sram_mem[92362] = 16'b0000000000000000;
	sram_mem[92363] = 16'b0000000000000000;
	sram_mem[92364] = 16'b0000000000000000;
	sram_mem[92365] = 16'b0000000000000000;
	sram_mem[92366] = 16'b0000000000000000;
	sram_mem[92367] = 16'b0000000000000000;
	sram_mem[92368] = 16'b0000000000000000;
	sram_mem[92369] = 16'b0000000000000000;
	sram_mem[92370] = 16'b0000000000000000;
	sram_mem[92371] = 16'b0000000000000000;
	sram_mem[92372] = 16'b0000000000000000;
	sram_mem[92373] = 16'b0000000000000000;
	sram_mem[92374] = 16'b0000000000000000;
	sram_mem[92375] = 16'b0000000000000000;
	sram_mem[92376] = 16'b0000000000000000;
	sram_mem[92377] = 16'b0000000000000000;
	sram_mem[92378] = 16'b0000000000000000;
	sram_mem[92379] = 16'b0000000000000000;
	sram_mem[92380] = 16'b0000000000000000;
	sram_mem[92381] = 16'b0000000000000000;
	sram_mem[92382] = 16'b0000000000000000;
	sram_mem[92383] = 16'b0000000000000000;
	sram_mem[92384] = 16'b0000000000000000;
	sram_mem[92385] = 16'b0000000000000000;
	sram_mem[92386] = 16'b0000000000000000;
	sram_mem[92387] = 16'b0000000000000000;
	sram_mem[92388] = 16'b0000000000000000;
	sram_mem[92389] = 16'b0000000000000000;
	sram_mem[92390] = 16'b0000000000000000;
	sram_mem[92391] = 16'b0000000000000000;
	sram_mem[92392] = 16'b0000000000000000;
	sram_mem[92393] = 16'b0000000000000000;
	sram_mem[92394] = 16'b0000000000000000;
	sram_mem[92395] = 16'b0000000000000000;
	sram_mem[92396] = 16'b0000000000000000;
	sram_mem[92397] = 16'b0000000000000000;
	sram_mem[92398] = 16'b0000000000000000;
	sram_mem[92399] = 16'b0000000000000000;
	sram_mem[92400] = 16'b0000000000000000;
	sram_mem[92401] = 16'b0000000000000000;
	sram_mem[92402] = 16'b0000000000000000;
	sram_mem[92403] = 16'b0000000000000000;
	sram_mem[92404] = 16'b0000000000000000;
	sram_mem[92405] = 16'b0000000000000000;
	sram_mem[92406] = 16'b0000000000000000;
	sram_mem[92407] = 16'b0000000000000000;
	sram_mem[92408] = 16'b0000000000000000;
	sram_mem[92409] = 16'b0000000000000000;
	sram_mem[92410] = 16'b0000000000000000;
	sram_mem[92411] = 16'b0000000000000000;
	sram_mem[92412] = 16'b0000000000000000;
	sram_mem[92413] = 16'b0000000000000000;
	sram_mem[92414] = 16'b0000000000000000;
	sram_mem[92415] = 16'b0000000000000000;
	sram_mem[92416] = 16'b0000000000000000;
	sram_mem[92417] = 16'b0000000000000000;
	sram_mem[92418] = 16'b0000000000000000;
	sram_mem[92419] = 16'b0000000000000000;
	sram_mem[92420] = 16'b0000000000000000;
	sram_mem[92421] = 16'b0000000000000000;
	sram_mem[92422] = 16'b0000000000000000;
	sram_mem[92423] = 16'b0000000000000000;
	sram_mem[92424] = 16'b0000000000000000;
	sram_mem[92425] = 16'b0000000000000000;
	sram_mem[92426] = 16'b0000000000000000;
	sram_mem[92427] = 16'b0000000000000000;
	sram_mem[92428] = 16'b0000000000000000;
	sram_mem[92429] = 16'b0000000000000000;
	sram_mem[92430] = 16'b0000000000000000;
	sram_mem[92431] = 16'b0000000000000000;
	sram_mem[92432] = 16'b0000000000000000;
	sram_mem[92433] = 16'b0000000000000000;
	sram_mem[92434] = 16'b0000000000000000;
	sram_mem[92435] = 16'b0000000000000000;
	sram_mem[92436] = 16'b0000000000000000;
	sram_mem[92437] = 16'b0000000000000000;
	sram_mem[92438] = 16'b0000000000000000;
	sram_mem[92439] = 16'b0000000000000000;
	sram_mem[92440] = 16'b0000000000000000;
	sram_mem[92441] = 16'b0000000000000000;
	sram_mem[92442] = 16'b0000000000000000;
	sram_mem[92443] = 16'b0000000000000000;
	sram_mem[92444] = 16'b0000000000000000;
	sram_mem[92445] = 16'b0000000000000000;
	sram_mem[92446] = 16'b0000000000000000;
	sram_mem[92447] = 16'b0000000000000000;
	sram_mem[92448] = 16'b0000000000000000;
	sram_mem[92449] = 16'b0000000000000000;
	sram_mem[92450] = 16'b0000000000000000;
	sram_mem[92451] = 16'b0000000000000000;
	sram_mem[92452] = 16'b0000000000000000;
	sram_mem[92453] = 16'b0000000000000000;
	sram_mem[92454] = 16'b0000000000000000;
	sram_mem[92455] = 16'b0000000000000000;
	sram_mem[92456] = 16'b0000000000000000;
	sram_mem[92457] = 16'b0000000000000000;
	sram_mem[92458] = 16'b0000000000000000;
	sram_mem[92459] = 16'b0000000000000000;
	sram_mem[92460] = 16'b0000000000000000;
	sram_mem[92461] = 16'b0000000000000000;
	sram_mem[92462] = 16'b0000000000000000;
	sram_mem[92463] = 16'b0000000000000000;
	sram_mem[92464] = 16'b0000000000000000;
	sram_mem[92465] = 16'b0000000000000000;
	sram_mem[92466] = 16'b0000000000000000;
	sram_mem[92467] = 16'b0000000000000000;
	sram_mem[92468] = 16'b0000000000000000;
	sram_mem[92469] = 16'b0000000000000000;
	sram_mem[92470] = 16'b0000000000000000;
	sram_mem[92471] = 16'b0000000000000000;
	sram_mem[92472] = 16'b0000000000000000;
	sram_mem[92473] = 16'b0000000000000000;
	sram_mem[92474] = 16'b0000000000000000;
	sram_mem[92475] = 16'b0000000000000000;
	sram_mem[92476] = 16'b0000000000000000;
	sram_mem[92477] = 16'b0000000000000000;
	sram_mem[92478] = 16'b0000000000000000;
	sram_mem[92479] = 16'b0000000000000000;
	sram_mem[92480] = 16'b0000000000000000;
	sram_mem[92481] = 16'b0000000000000000;
	sram_mem[92482] = 16'b0000000000000000;
	sram_mem[92483] = 16'b0000000000000000;
	sram_mem[92484] = 16'b0000000000000000;
	sram_mem[92485] = 16'b0000000000000000;
	sram_mem[92486] = 16'b0000000000000000;
	sram_mem[92487] = 16'b0000000000000000;
	sram_mem[92488] = 16'b0000000000000000;
	sram_mem[92489] = 16'b0000000000000000;
	sram_mem[92490] = 16'b0000000000000000;
	sram_mem[92491] = 16'b0000000000000000;
	sram_mem[92492] = 16'b0000000000000000;
	sram_mem[92493] = 16'b0000000000000000;
	sram_mem[92494] = 16'b0000000000000000;
	sram_mem[92495] = 16'b0000000000000000;
	sram_mem[92496] = 16'b0000000000000000;
	sram_mem[92497] = 16'b0000000000000000;
	sram_mem[92498] = 16'b0000000000000000;
	sram_mem[92499] = 16'b0000000000000000;
	sram_mem[92500] = 16'b0000000000000000;
	sram_mem[92501] = 16'b0000000000000000;
	sram_mem[92502] = 16'b0000000000000000;
	sram_mem[92503] = 16'b0000000000000000;
	sram_mem[92504] = 16'b0000000000000000;
	sram_mem[92505] = 16'b0000000000000000;
	sram_mem[92506] = 16'b0000000000000000;
	sram_mem[92507] = 16'b0000000000000000;
	sram_mem[92508] = 16'b0000000000000000;
	sram_mem[92509] = 16'b0000000000000000;
	sram_mem[92510] = 16'b0000000000000000;
	sram_mem[92511] = 16'b0000000000000000;
	sram_mem[92512] = 16'b0000000000000000;
	sram_mem[92513] = 16'b0000000000000000;
	sram_mem[92514] = 16'b0000000000000000;
	sram_mem[92515] = 16'b0000000000000000;
	sram_mem[92516] = 16'b0000000000000000;
	sram_mem[92517] = 16'b0000000000000000;
	sram_mem[92518] = 16'b0000000000000000;
	sram_mem[92519] = 16'b0000000000000000;
	sram_mem[92520] = 16'b0000000000000000;
	sram_mem[92521] = 16'b0000000000000000;
	sram_mem[92522] = 16'b0000000000000000;
	sram_mem[92523] = 16'b0000000000000000;
	sram_mem[92524] = 16'b0000000000000000;
	sram_mem[92525] = 16'b0000000000000000;
	sram_mem[92526] = 16'b0000000000000000;
	sram_mem[92527] = 16'b0000000000000000;
	sram_mem[92528] = 16'b0000000000000000;
	sram_mem[92529] = 16'b0000000000000000;
	sram_mem[92530] = 16'b0000000000000000;
	sram_mem[92531] = 16'b0000000000000000;
	sram_mem[92532] = 16'b0000000000000000;
	sram_mem[92533] = 16'b0000000000000000;
	sram_mem[92534] = 16'b0000000000000000;
	sram_mem[92535] = 16'b0000000000000000;
	sram_mem[92536] = 16'b0000000000000000;
	sram_mem[92537] = 16'b0000000000000000;
	sram_mem[92538] = 16'b0000000000000000;
	sram_mem[92539] = 16'b0000000000000000;
	sram_mem[92540] = 16'b0000000000000000;
	sram_mem[92541] = 16'b0000000000000000;
	sram_mem[92542] = 16'b0000000000000000;
	sram_mem[92543] = 16'b0000000000000000;
	sram_mem[92544] = 16'b0000000000000000;
	sram_mem[92545] = 16'b0000000000000000;
	sram_mem[92546] = 16'b0000000000000000;
	sram_mem[92547] = 16'b0000000000000000;
	sram_mem[92548] = 16'b0000000000000000;
	sram_mem[92549] = 16'b0000000000000000;
	sram_mem[92550] = 16'b0000000000000000;
	sram_mem[92551] = 16'b0000000000000000;
	sram_mem[92552] = 16'b0000000000000000;
	sram_mem[92553] = 16'b0000000000000000;
	sram_mem[92554] = 16'b0000000000000000;
	sram_mem[92555] = 16'b0000000000000000;
	sram_mem[92556] = 16'b0000000000000000;
	sram_mem[92557] = 16'b0000000000000000;
	sram_mem[92558] = 16'b0000000000000000;
	sram_mem[92559] = 16'b0000000000000000;
	sram_mem[92560] = 16'b0000000000000000;
	sram_mem[92561] = 16'b0000000000000000;
	sram_mem[92562] = 16'b0000000000000000;
	sram_mem[92563] = 16'b0000000000000000;
	sram_mem[92564] = 16'b0000000000000000;
	sram_mem[92565] = 16'b0000000000000000;
	sram_mem[92566] = 16'b0000000000000000;
	sram_mem[92567] = 16'b0000000000000000;
	sram_mem[92568] = 16'b0000000000000000;
	sram_mem[92569] = 16'b0000000000000000;
	sram_mem[92570] = 16'b0000000000000000;
	sram_mem[92571] = 16'b0000000000000000;
	sram_mem[92572] = 16'b0000000000000000;
	sram_mem[92573] = 16'b0000000000000000;
	sram_mem[92574] = 16'b0000000000000000;
	sram_mem[92575] = 16'b0000000000000000;
	sram_mem[92576] = 16'b0000000000000000;
	sram_mem[92577] = 16'b0000000000000000;
	sram_mem[92578] = 16'b0000000000000000;
	sram_mem[92579] = 16'b0000000000000000;
	sram_mem[92580] = 16'b0000000000000000;
	sram_mem[92581] = 16'b0000000000000000;
	sram_mem[92582] = 16'b0000000000000000;
	sram_mem[92583] = 16'b0000000000000000;
	sram_mem[92584] = 16'b0000000000000000;
	sram_mem[92585] = 16'b0000000000000000;
	sram_mem[92586] = 16'b0000000000000000;
	sram_mem[92587] = 16'b0000000000000000;
	sram_mem[92588] = 16'b0000000000000000;
	sram_mem[92589] = 16'b0000000000000000;
	sram_mem[92590] = 16'b0000000000000000;
	sram_mem[92591] = 16'b0000000000000000;
	sram_mem[92592] = 16'b0000000000000000;
	sram_mem[92593] = 16'b0000000000000000;
	sram_mem[92594] = 16'b0000000000000000;
	sram_mem[92595] = 16'b0000000000000000;
	sram_mem[92596] = 16'b0000000000000000;
	sram_mem[92597] = 16'b0000000000000000;
	sram_mem[92598] = 16'b0000000000000000;
	sram_mem[92599] = 16'b0000000000000000;
	sram_mem[92600] = 16'b0000000000000000;
	sram_mem[92601] = 16'b0000000000000000;
	sram_mem[92602] = 16'b0000000000000000;
	sram_mem[92603] = 16'b0000000000000000;
	sram_mem[92604] = 16'b0000000000000000;
	sram_mem[92605] = 16'b0000000000000000;
	sram_mem[92606] = 16'b0000000000000000;
	sram_mem[92607] = 16'b0000000000000000;
	sram_mem[92608] = 16'b0000000000000000;
	sram_mem[92609] = 16'b0000000000000000;
	sram_mem[92610] = 16'b0000000000000000;
	sram_mem[92611] = 16'b0000000000000000;
	sram_mem[92612] = 16'b0000000000000000;
	sram_mem[92613] = 16'b0000000000000000;
	sram_mem[92614] = 16'b0000000000000000;
	sram_mem[92615] = 16'b0000000000000000;
	sram_mem[92616] = 16'b0000000000000000;
	sram_mem[92617] = 16'b0000000000000000;
	sram_mem[92618] = 16'b0000000000000000;
	sram_mem[92619] = 16'b0000000000000000;
	sram_mem[92620] = 16'b0000000000000000;
	sram_mem[92621] = 16'b0000000000000000;
	sram_mem[92622] = 16'b0000000000000000;
	sram_mem[92623] = 16'b0000000000000000;
	sram_mem[92624] = 16'b0000000000000000;
	sram_mem[92625] = 16'b0000000000000000;
	sram_mem[92626] = 16'b0000000000000000;
	sram_mem[92627] = 16'b0000000000000000;
	sram_mem[92628] = 16'b0000000000000000;
	sram_mem[92629] = 16'b0000000000000000;
	sram_mem[92630] = 16'b0000000000000000;
	sram_mem[92631] = 16'b0000000000000000;
	sram_mem[92632] = 16'b0000000000000000;
	sram_mem[92633] = 16'b0000000000000000;
	sram_mem[92634] = 16'b0000000000000000;
	sram_mem[92635] = 16'b0000000000000000;
	sram_mem[92636] = 16'b0000000000000000;
	sram_mem[92637] = 16'b0000000000000000;
	sram_mem[92638] = 16'b0000000000000000;
	sram_mem[92639] = 16'b0000000000000000;
	sram_mem[92640] = 16'b0000000000000000;
	sram_mem[92641] = 16'b0000000000000000;
	sram_mem[92642] = 16'b0000000000000000;
	sram_mem[92643] = 16'b0000000000000000;
	sram_mem[92644] = 16'b0000000000000000;
	sram_mem[92645] = 16'b0000000000000000;
	sram_mem[92646] = 16'b0000000000000000;
	sram_mem[92647] = 16'b0000000000000000;
	sram_mem[92648] = 16'b0000000000000000;
	sram_mem[92649] = 16'b0000000000000000;
	sram_mem[92650] = 16'b0000000000000000;
	sram_mem[92651] = 16'b0000000000000000;
	sram_mem[92652] = 16'b0000000000000000;
	sram_mem[92653] = 16'b0000000000000000;
	sram_mem[92654] = 16'b0000000000000000;
	sram_mem[92655] = 16'b0000000000000000;
	sram_mem[92656] = 16'b0000000000000000;
	sram_mem[92657] = 16'b0000000000000000;
	sram_mem[92658] = 16'b0000000000000000;
	sram_mem[92659] = 16'b0000000000000000;
	sram_mem[92660] = 16'b0000000000000000;
	sram_mem[92661] = 16'b0000000000000000;
	sram_mem[92662] = 16'b0000000000000000;
	sram_mem[92663] = 16'b0000000000000000;
	sram_mem[92664] = 16'b0000000000000000;
	sram_mem[92665] = 16'b0000000000000000;
	sram_mem[92666] = 16'b0000000000000000;
	sram_mem[92667] = 16'b0000000000000000;
	sram_mem[92668] = 16'b0000000000000000;
	sram_mem[92669] = 16'b0000000000000000;
	sram_mem[92670] = 16'b0000000000000000;
	sram_mem[92671] = 16'b0000000000000000;
	sram_mem[92672] = 16'b0000000000000000;
	sram_mem[92673] = 16'b0000000000000000;
	sram_mem[92674] = 16'b0000000000000000;
	sram_mem[92675] = 16'b0000000000000000;
	sram_mem[92676] = 16'b0000000000000000;
	sram_mem[92677] = 16'b0000000000000000;
	sram_mem[92678] = 16'b0000000000000000;
	sram_mem[92679] = 16'b0000000000000000;
	sram_mem[92680] = 16'b0000000000000000;
	sram_mem[92681] = 16'b0000000000000000;
	sram_mem[92682] = 16'b0000000000000000;
	sram_mem[92683] = 16'b0000000000000000;
	sram_mem[92684] = 16'b0000000000000000;
	sram_mem[92685] = 16'b0000000000000000;
	sram_mem[92686] = 16'b0000000000000000;
	sram_mem[92687] = 16'b0000000000000000;
	sram_mem[92688] = 16'b0000000000000000;
	sram_mem[92689] = 16'b0000000000000000;
	sram_mem[92690] = 16'b0000000000000000;
	sram_mem[92691] = 16'b0000000000000000;
	sram_mem[92692] = 16'b0000000000000000;
	sram_mem[92693] = 16'b0000000000000000;
	sram_mem[92694] = 16'b0000000000000000;
	sram_mem[92695] = 16'b0000000000000000;
	sram_mem[92696] = 16'b0000000000000000;
	sram_mem[92697] = 16'b0000000000000000;
	sram_mem[92698] = 16'b0000000000000000;
	sram_mem[92699] = 16'b0000000000000000;
	sram_mem[92700] = 16'b0000000000000000;
	sram_mem[92701] = 16'b0000000000000000;
	sram_mem[92702] = 16'b0000000000000000;
	sram_mem[92703] = 16'b0000000000000000;
	sram_mem[92704] = 16'b0000000000000000;
	sram_mem[92705] = 16'b0000000000000000;
	sram_mem[92706] = 16'b0000000000000000;
	sram_mem[92707] = 16'b0000000000000000;
	sram_mem[92708] = 16'b0000000000000000;
	sram_mem[92709] = 16'b0000000000000000;
	sram_mem[92710] = 16'b0000000000000000;
	sram_mem[92711] = 16'b0000000000000000;
	sram_mem[92712] = 16'b0000000000000000;
	sram_mem[92713] = 16'b0000000000000000;
	sram_mem[92714] = 16'b0000000000000000;
	sram_mem[92715] = 16'b0000000000000000;
	sram_mem[92716] = 16'b0000000000000000;
	sram_mem[92717] = 16'b0000000000000000;
	sram_mem[92718] = 16'b0000000000000000;
	sram_mem[92719] = 16'b0000000000000000;
	sram_mem[92720] = 16'b0000000000000000;
	sram_mem[92721] = 16'b0000000000000000;
	sram_mem[92722] = 16'b0000000000000000;
	sram_mem[92723] = 16'b0000000000000000;
	sram_mem[92724] = 16'b0000000000000000;
	sram_mem[92725] = 16'b0000000000000000;
	sram_mem[92726] = 16'b0000000000000000;
	sram_mem[92727] = 16'b0000000000000000;
	sram_mem[92728] = 16'b0000000000000000;
	sram_mem[92729] = 16'b0000000000000000;
	sram_mem[92730] = 16'b0000000000000000;
	sram_mem[92731] = 16'b0000000000000000;
	sram_mem[92732] = 16'b0000000000000000;
	sram_mem[92733] = 16'b0000000000000000;
	sram_mem[92734] = 16'b0000000000000000;
	sram_mem[92735] = 16'b0000000000000000;
	sram_mem[92736] = 16'b0000000000000000;
	sram_mem[92737] = 16'b0000000000000000;
	sram_mem[92738] = 16'b0000000000000000;
	sram_mem[92739] = 16'b0000000000000000;
	sram_mem[92740] = 16'b0000000000000000;
	sram_mem[92741] = 16'b0000000000000000;
	sram_mem[92742] = 16'b0000000000000000;
	sram_mem[92743] = 16'b0000000000000000;
	sram_mem[92744] = 16'b0000000000000000;
	sram_mem[92745] = 16'b0000000000000000;
	sram_mem[92746] = 16'b0000000000000000;
	sram_mem[92747] = 16'b0000000000000000;
	sram_mem[92748] = 16'b0000000000000000;
	sram_mem[92749] = 16'b0000000000000000;
	sram_mem[92750] = 16'b0000000000000000;
	sram_mem[92751] = 16'b0000000000000000;
	sram_mem[92752] = 16'b0000000000000000;
	sram_mem[92753] = 16'b0000000000000000;
	sram_mem[92754] = 16'b0000000000000000;
	sram_mem[92755] = 16'b0000000000000000;
	sram_mem[92756] = 16'b0000000000000000;
	sram_mem[92757] = 16'b0000000000000000;
	sram_mem[92758] = 16'b0000000000000000;
	sram_mem[92759] = 16'b0000000000000000;
	sram_mem[92760] = 16'b0000000000000000;
	sram_mem[92761] = 16'b0000000000000000;
	sram_mem[92762] = 16'b0000000000000000;
	sram_mem[92763] = 16'b0000000000000000;
	sram_mem[92764] = 16'b0000000000000000;
	sram_mem[92765] = 16'b0000000000000000;
	sram_mem[92766] = 16'b0000000000000000;
	sram_mem[92767] = 16'b0000000000000000;
	sram_mem[92768] = 16'b0000000000000000;
	sram_mem[92769] = 16'b0000000000000000;
	sram_mem[92770] = 16'b0000000000000000;
	sram_mem[92771] = 16'b0000000000000000;
	sram_mem[92772] = 16'b0000000000000000;
	sram_mem[92773] = 16'b0000000000000000;
	sram_mem[92774] = 16'b0000000000000000;
	sram_mem[92775] = 16'b0000000000000000;
	sram_mem[92776] = 16'b0000000000000000;
	sram_mem[92777] = 16'b0000000000000000;
	sram_mem[92778] = 16'b0000000000000000;
	sram_mem[92779] = 16'b0000000000000000;
	sram_mem[92780] = 16'b0000000000000000;
	sram_mem[92781] = 16'b0000000000000000;
	sram_mem[92782] = 16'b0000000000000000;
	sram_mem[92783] = 16'b0000000000000000;
	sram_mem[92784] = 16'b0000000000000000;
	sram_mem[92785] = 16'b0000000000000000;
	sram_mem[92786] = 16'b0000000000000000;
	sram_mem[92787] = 16'b0000000000000000;
	sram_mem[92788] = 16'b0000000000000000;
	sram_mem[92789] = 16'b0000000000000000;
	sram_mem[92790] = 16'b0000000000000000;
	sram_mem[92791] = 16'b0000000000000000;
	sram_mem[92792] = 16'b0000000000000000;
	sram_mem[92793] = 16'b0000000000000000;
	sram_mem[92794] = 16'b0000000000000000;
	sram_mem[92795] = 16'b0000000000000000;
	sram_mem[92796] = 16'b0000000000000000;
	sram_mem[92797] = 16'b0000000000000000;
	sram_mem[92798] = 16'b0000000000000000;
	sram_mem[92799] = 16'b0000000000000000;
	sram_mem[92800] = 16'b0000000000000000;
	sram_mem[92801] = 16'b0000000000000000;
	sram_mem[92802] = 16'b0000000000000000;
	sram_mem[92803] = 16'b0000000000000000;
	sram_mem[92804] = 16'b0000000000000000;
	sram_mem[92805] = 16'b0000000000000000;
	sram_mem[92806] = 16'b0000000000000000;
	sram_mem[92807] = 16'b0000000000000000;
	sram_mem[92808] = 16'b0000000000000000;
	sram_mem[92809] = 16'b0000000000000000;
	sram_mem[92810] = 16'b0000000000000000;
	sram_mem[92811] = 16'b0000000000000000;
	sram_mem[92812] = 16'b0000000000000000;
	sram_mem[92813] = 16'b0000000000000000;
	sram_mem[92814] = 16'b0000000000000000;
	sram_mem[92815] = 16'b0000000000000000;
	sram_mem[92816] = 16'b0000000000000000;
	sram_mem[92817] = 16'b0000000000000000;
	sram_mem[92818] = 16'b0000000000000000;
	sram_mem[92819] = 16'b0000000000000000;
	sram_mem[92820] = 16'b0000000000000000;
	sram_mem[92821] = 16'b0000000000000000;
	sram_mem[92822] = 16'b0000000000000000;
	sram_mem[92823] = 16'b0000000000000000;
	sram_mem[92824] = 16'b0000000000000000;
	sram_mem[92825] = 16'b0000000000000000;
	sram_mem[92826] = 16'b0000000000000000;
	sram_mem[92827] = 16'b0000000000000000;
	sram_mem[92828] = 16'b0000000000000000;
	sram_mem[92829] = 16'b0000000000000000;
	sram_mem[92830] = 16'b0000000000000000;
	sram_mem[92831] = 16'b0000000000000000;
	sram_mem[92832] = 16'b0000000000000000;
	sram_mem[92833] = 16'b0000000000000000;
	sram_mem[92834] = 16'b0000000000000000;
	sram_mem[92835] = 16'b0000000000000000;
	sram_mem[92836] = 16'b0000000000000000;
	sram_mem[92837] = 16'b0000000000000000;
	sram_mem[92838] = 16'b0000000000000000;
	sram_mem[92839] = 16'b0000000000000000;
	sram_mem[92840] = 16'b0000000000000000;
	sram_mem[92841] = 16'b0000000000000000;
	sram_mem[92842] = 16'b0000000000000000;
	sram_mem[92843] = 16'b0000000000000000;
	sram_mem[92844] = 16'b0000000000000000;
	sram_mem[92845] = 16'b0000000000000000;
	sram_mem[92846] = 16'b0000000000000000;
	sram_mem[92847] = 16'b0000000000000000;
	sram_mem[92848] = 16'b0000000000000000;
	sram_mem[92849] = 16'b0000000000000000;
	sram_mem[92850] = 16'b0000000000000000;
	sram_mem[92851] = 16'b0000000000000000;
	sram_mem[92852] = 16'b0000000000000000;
	sram_mem[92853] = 16'b0000000000000000;
	sram_mem[92854] = 16'b0000000000000000;
	sram_mem[92855] = 16'b0000000000000000;
	sram_mem[92856] = 16'b0000000000000000;
	sram_mem[92857] = 16'b0000000000000000;
	sram_mem[92858] = 16'b0000000000000000;
	sram_mem[92859] = 16'b0000000000000000;
	sram_mem[92860] = 16'b0000000000000000;
	sram_mem[92861] = 16'b0000000000000000;
	sram_mem[92862] = 16'b0000000000000000;
	sram_mem[92863] = 16'b0000000000000000;
	sram_mem[92864] = 16'b0000000000000000;
	sram_mem[92865] = 16'b0000000000000000;
	sram_mem[92866] = 16'b0000000000000000;
	sram_mem[92867] = 16'b0000000000000000;
	sram_mem[92868] = 16'b0000000000000000;
	sram_mem[92869] = 16'b0000000000000000;
	sram_mem[92870] = 16'b0000000000000000;
	sram_mem[92871] = 16'b0000000000000000;
	sram_mem[92872] = 16'b0000000000000000;
	sram_mem[92873] = 16'b0000000000000000;
	sram_mem[92874] = 16'b0000000000000000;
	sram_mem[92875] = 16'b0000000000000000;
	sram_mem[92876] = 16'b0000000000000000;
	sram_mem[92877] = 16'b0000000000000000;
	sram_mem[92878] = 16'b0000000000000000;
	sram_mem[92879] = 16'b0000000000000000;
	sram_mem[92880] = 16'b0000000000000000;
	sram_mem[92881] = 16'b0000000000000000;
	sram_mem[92882] = 16'b0000000000000000;
	sram_mem[92883] = 16'b0000000000000000;
	sram_mem[92884] = 16'b0000000000000000;
	sram_mem[92885] = 16'b0000000000000000;
	sram_mem[92886] = 16'b0000000000000000;
	sram_mem[92887] = 16'b0000000000000000;
	sram_mem[92888] = 16'b0000000000000000;
	sram_mem[92889] = 16'b0000000000000000;
	sram_mem[92890] = 16'b0000000000000000;
	sram_mem[92891] = 16'b0000000000000000;
	sram_mem[92892] = 16'b0000000000000000;
	sram_mem[92893] = 16'b0000000000000000;
	sram_mem[92894] = 16'b0000000000000000;
	sram_mem[92895] = 16'b0000000000000000;
	sram_mem[92896] = 16'b0000000000000000;
	sram_mem[92897] = 16'b0000000000000000;
	sram_mem[92898] = 16'b0000000000000000;
	sram_mem[92899] = 16'b0000000000000000;
	sram_mem[92900] = 16'b0000000000000000;
	sram_mem[92901] = 16'b0000000000000000;
	sram_mem[92902] = 16'b0000000000000000;
	sram_mem[92903] = 16'b0000000000000000;
	sram_mem[92904] = 16'b0000000000000000;
	sram_mem[92905] = 16'b0000000000000000;
	sram_mem[92906] = 16'b0000000000000000;
	sram_mem[92907] = 16'b0000000000000000;
	sram_mem[92908] = 16'b0000000000000000;
	sram_mem[92909] = 16'b0000000000000000;
	sram_mem[92910] = 16'b0000000000000000;
	sram_mem[92911] = 16'b0000000000000000;
	sram_mem[92912] = 16'b0000000000000000;
	sram_mem[92913] = 16'b0000000000000000;
	sram_mem[92914] = 16'b0000000000000000;
	sram_mem[92915] = 16'b0000000000000000;
	sram_mem[92916] = 16'b0000000000000000;
	sram_mem[92917] = 16'b0000000000000000;
	sram_mem[92918] = 16'b0000000000000000;
	sram_mem[92919] = 16'b0000000000000000;
	sram_mem[92920] = 16'b0000000000000000;
	sram_mem[92921] = 16'b0000000000000000;
	sram_mem[92922] = 16'b0000000000000000;
	sram_mem[92923] = 16'b0000000000000000;
	sram_mem[92924] = 16'b0000000000000000;
	sram_mem[92925] = 16'b0000000000000000;
	sram_mem[92926] = 16'b0000000000000000;
	sram_mem[92927] = 16'b0000000000000000;
	sram_mem[92928] = 16'b0000000000000000;
	sram_mem[92929] = 16'b0000000000000000;
	sram_mem[92930] = 16'b0000000000000000;
	sram_mem[92931] = 16'b0000000000000000;
	sram_mem[92932] = 16'b0000000000000000;
	sram_mem[92933] = 16'b0000000000000000;
	sram_mem[92934] = 16'b0000000000000000;
	sram_mem[92935] = 16'b0000000000000000;
	sram_mem[92936] = 16'b0000000000000000;
	sram_mem[92937] = 16'b0000000000000000;
	sram_mem[92938] = 16'b0000000000000000;
	sram_mem[92939] = 16'b0000000000000000;
	sram_mem[92940] = 16'b0000000000000000;
	sram_mem[92941] = 16'b0000000000000000;
	sram_mem[92942] = 16'b0000000000000000;
	sram_mem[92943] = 16'b0000000000000000;
	sram_mem[92944] = 16'b0000000000000000;
	sram_mem[92945] = 16'b0000000000000000;
	sram_mem[92946] = 16'b0000000000000000;
	sram_mem[92947] = 16'b0000000000000000;
	sram_mem[92948] = 16'b0000000000000000;
	sram_mem[92949] = 16'b0000000000000000;
	sram_mem[92950] = 16'b0000000000000000;
	sram_mem[92951] = 16'b0000000000000000;
	sram_mem[92952] = 16'b0000000000000000;
	sram_mem[92953] = 16'b0000000000000000;
	sram_mem[92954] = 16'b0000000000000000;
	sram_mem[92955] = 16'b0000000000000000;
	sram_mem[92956] = 16'b0000000000000000;
	sram_mem[92957] = 16'b0000000000000000;
	sram_mem[92958] = 16'b0000000000000000;
	sram_mem[92959] = 16'b0000000000000000;
	sram_mem[92960] = 16'b0000000000000000;
	sram_mem[92961] = 16'b0000000000000000;
	sram_mem[92962] = 16'b0000000000000000;
	sram_mem[92963] = 16'b0000000000000000;
	sram_mem[92964] = 16'b0000000000000000;
	sram_mem[92965] = 16'b0000000000000000;
	sram_mem[92966] = 16'b0000000000000000;
	sram_mem[92967] = 16'b0000000000000000;
	sram_mem[92968] = 16'b0000000000000000;
	sram_mem[92969] = 16'b0000000000000000;
	sram_mem[92970] = 16'b0000000000000000;
	sram_mem[92971] = 16'b0000000000000000;
	sram_mem[92972] = 16'b0000000000000000;
	sram_mem[92973] = 16'b0000000000000000;
	sram_mem[92974] = 16'b0000000000000000;
	sram_mem[92975] = 16'b0000000000000000;
	sram_mem[92976] = 16'b0000000000000000;
	sram_mem[92977] = 16'b0000000000000000;
	sram_mem[92978] = 16'b0000000000000000;
	sram_mem[92979] = 16'b0000000000000000;
	sram_mem[92980] = 16'b0000000000000000;
	sram_mem[92981] = 16'b0000000000000000;
	sram_mem[92982] = 16'b0000000000000000;
	sram_mem[92983] = 16'b0000000000000000;
	sram_mem[92984] = 16'b0000000000000000;
	sram_mem[92985] = 16'b0000000000000000;
	sram_mem[92986] = 16'b0000000000000000;
	sram_mem[92987] = 16'b0000000000000000;
	sram_mem[92988] = 16'b0000000000000000;
	sram_mem[92989] = 16'b0000000000000000;
	sram_mem[92990] = 16'b0000000000000000;
	sram_mem[92991] = 16'b0000000000000000;
	sram_mem[92992] = 16'b0000000000000000;
	sram_mem[92993] = 16'b0000000000000000;
	sram_mem[92994] = 16'b0000000000000000;
	sram_mem[92995] = 16'b0000000000000000;
	sram_mem[92996] = 16'b0000000000000000;
	sram_mem[92997] = 16'b0000000000000000;
	sram_mem[92998] = 16'b0000000000000000;
	sram_mem[92999] = 16'b0000000000000000;
	sram_mem[93000] = 16'b0000000000000000;
	sram_mem[93001] = 16'b0000000000000000;
	sram_mem[93002] = 16'b0000000000000000;
	sram_mem[93003] = 16'b0000000000000000;
	sram_mem[93004] = 16'b0000000000000000;
	sram_mem[93005] = 16'b0000000000000000;
	sram_mem[93006] = 16'b0000000000000000;
	sram_mem[93007] = 16'b0000000000000000;
	sram_mem[93008] = 16'b0000000000000000;
	sram_mem[93009] = 16'b0000000000000000;
	sram_mem[93010] = 16'b0000000000000000;
	sram_mem[93011] = 16'b0000000000000000;
	sram_mem[93012] = 16'b0000000000000000;
	sram_mem[93013] = 16'b0000000000000000;
	sram_mem[93014] = 16'b0000000000000000;
	sram_mem[93015] = 16'b0000000000000000;
	sram_mem[93016] = 16'b0000000000000000;
	sram_mem[93017] = 16'b0000000000000000;
	sram_mem[93018] = 16'b0000000000000000;
	sram_mem[93019] = 16'b0000000000000000;
	sram_mem[93020] = 16'b0000000000000000;
	sram_mem[93021] = 16'b0000000000000000;
	sram_mem[93022] = 16'b0000000000000000;
	sram_mem[93023] = 16'b0000000000000000;
	sram_mem[93024] = 16'b0000000000000000;
	sram_mem[93025] = 16'b0000000000000000;
	sram_mem[93026] = 16'b0000000000000000;
	sram_mem[93027] = 16'b0000000000000000;
	sram_mem[93028] = 16'b0000000000000000;
	sram_mem[93029] = 16'b0000000000000000;
	sram_mem[93030] = 16'b0000000000000000;
	sram_mem[93031] = 16'b0000000000000000;
	sram_mem[93032] = 16'b0000000000000000;
	sram_mem[93033] = 16'b0000000000000000;
	sram_mem[93034] = 16'b0000000000000000;
	sram_mem[93035] = 16'b0000000000000000;
	sram_mem[93036] = 16'b0000000000000000;
	sram_mem[93037] = 16'b0000000000000000;
	sram_mem[93038] = 16'b0000000000000000;
	sram_mem[93039] = 16'b0000000000000000;
	sram_mem[93040] = 16'b0000000000000000;
	sram_mem[93041] = 16'b0000000000000000;
	sram_mem[93042] = 16'b0000000000000000;
	sram_mem[93043] = 16'b0000000000000000;
	sram_mem[93044] = 16'b0000000000000000;
	sram_mem[93045] = 16'b0000000000000000;
	sram_mem[93046] = 16'b0000000000000000;
	sram_mem[93047] = 16'b0000000000000000;
	sram_mem[93048] = 16'b0000000000000000;
	sram_mem[93049] = 16'b0000000000000000;
	sram_mem[93050] = 16'b0000000000000000;
	sram_mem[93051] = 16'b0000000000000000;
	sram_mem[93052] = 16'b0000000000000000;
	sram_mem[93053] = 16'b0000000000000000;
	sram_mem[93054] = 16'b0000000000000000;
	sram_mem[93055] = 16'b0000000000000000;
	sram_mem[93056] = 16'b0000000000000000;
	sram_mem[93057] = 16'b0000000000000000;
	sram_mem[93058] = 16'b0000000000000000;
	sram_mem[93059] = 16'b0000000000000000;
	sram_mem[93060] = 16'b0000000000000000;
	sram_mem[93061] = 16'b0000000000000000;
	sram_mem[93062] = 16'b0000000000000000;
	sram_mem[93063] = 16'b0000000000000000;
	sram_mem[93064] = 16'b0000000000000000;
	sram_mem[93065] = 16'b0000000000000000;
	sram_mem[93066] = 16'b0000000000000000;
	sram_mem[93067] = 16'b0000000000000000;
	sram_mem[93068] = 16'b0000000000000000;
	sram_mem[93069] = 16'b0000000000000000;
	sram_mem[93070] = 16'b0000000000000000;
	sram_mem[93071] = 16'b0000000000000000;
	sram_mem[93072] = 16'b0000000000000000;
	sram_mem[93073] = 16'b0000000000000000;
	sram_mem[93074] = 16'b0000000000000000;
	sram_mem[93075] = 16'b0000000000000000;
	sram_mem[93076] = 16'b0000000000000000;
	sram_mem[93077] = 16'b0000000000000000;
	sram_mem[93078] = 16'b0000000000000000;
	sram_mem[93079] = 16'b0000000000000000;
	sram_mem[93080] = 16'b0000000000000000;
	sram_mem[93081] = 16'b0000000000000000;
	sram_mem[93082] = 16'b0000000000000000;
	sram_mem[93083] = 16'b0000000000000000;
	sram_mem[93084] = 16'b0000000000000000;
	sram_mem[93085] = 16'b0000000000000000;
	sram_mem[93086] = 16'b0000000000000000;
	sram_mem[93087] = 16'b0000000000000000;
	sram_mem[93088] = 16'b0000000000000000;
	sram_mem[93089] = 16'b0000000000000000;
	sram_mem[93090] = 16'b0000000000000000;
	sram_mem[93091] = 16'b0000000000000000;
	sram_mem[93092] = 16'b0000000000000000;
	sram_mem[93093] = 16'b0000000000000000;
	sram_mem[93094] = 16'b0000000000000000;
	sram_mem[93095] = 16'b0000000000000000;
	sram_mem[93096] = 16'b0000000000000000;
	sram_mem[93097] = 16'b0000000000000000;
	sram_mem[93098] = 16'b0000000000000000;
	sram_mem[93099] = 16'b0000000000000000;
	sram_mem[93100] = 16'b0000000000000000;
	sram_mem[93101] = 16'b0000000000000000;
	sram_mem[93102] = 16'b0000000000000000;
	sram_mem[93103] = 16'b0000000000000000;
	sram_mem[93104] = 16'b0000000000000000;
	sram_mem[93105] = 16'b0000000000000000;
	sram_mem[93106] = 16'b0000000000000000;
	sram_mem[93107] = 16'b0000000000000000;
	sram_mem[93108] = 16'b0000000000000000;
	sram_mem[93109] = 16'b0000000000000000;
	sram_mem[93110] = 16'b0000000000000000;
	sram_mem[93111] = 16'b0000000000000000;
	sram_mem[93112] = 16'b0000000000000000;
	sram_mem[93113] = 16'b0000000000000000;
	sram_mem[93114] = 16'b0000000000000000;
	sram_mem[93115] = 16'b0000000000000000;
	sram_mem[93116] = 16'b0000000000000000;
	sram_mem[93117] = 16'b0000000000000000;
	sram_mem[93118] = 16'b0000000000000000;
	sram_mem[93119] = 16'b0000000000000000;
	sram_mem[93120] = 16'b0000000000000000;
	sram_mem[93121] = 16'b0000000000000000;
	sram_mem[93122] = 16'b0000000000000000;
	sram_mem[93123] = 16'b0000000000000000;
	sram_mem[93124] = 16'b0000000000000000;
	sram_mem[93125] = 16'b0000000000000000;
	sram_mem[93126] = 16'b0000000000000000;
	sram_mem[93127] = 16'b0000000000000000;
	sram_mem[93128] = 16'b0000000000000000;
	sram_mem[93129] = 16'b0000000000000000;
	sram_mem[93130] = 16'b0000000000000000;
	sram_mem[93131] = 16'b0000000000000000;
	sram_mem[93132] = 16'b0000000000000000;
	sram_mem[93133] = 16'b0000000000000000;
	sram_mem[93134] = 16'b0000000000000000;
	sram_mem[93135] = 16'b0000000000000000;
	sram_mem[93136] = 16'b0000000000000000;
	sram_mem[93137] = 16'b0000000000000000;
	sram_mem[93138] = 16'b0000000000000000;
	sram_mem[93139] = 16'b0000000000000000;
	sram_mem[93140] = 16'b0000000000000000;
	sram_mem[93141] = 16'b0000000000000000;
	sram_mem[93142] = 16'b0000000000000000;
	sram_mem[93143] = 16'b0000000000000000;
	sram_mem[93144] = 16'b0000000000000000;
	sram_mem[93145] = 16'b0000000000000000;
	sram_mem[93146] = 16'b0000000000000000;
	sram_mem[93147] = 16'b0000000000000000;
	sram_mem[93148] = 16'b0000000000000000;
	sram_mem[93149] = 16'b0000000000000000;
	sram_mem[93150] = 16'b0000000000000000;
	sram_mem[93151] = 16'b0000000000000000;
	sram_mem[93152] = 16'b0000000000000000;
	sram_mem[93153] = 16'b0000000000000000;
	sram_mem[93154] = 16'b0000000000000000;
	sram_mem[93155] = 16'b0000000000000000;
	sram_mem[93156] = 16'b0000000000000000;
	sram_mem[93157] = 16'b0000000000000000;
	sram_mem[93158] = 16'b0000000000000000;
	sram_mem[93159] = 16'b0000000000000000;
	sram_mem[93160] = 16'b0000000000000000;
	sram_mem[93161] = 16'b0000000000000000;
	sram_mem[93162] = 16'b0000000000000000;
	sram_mem[93163] = 16'b0000000000000000;
	sram_mem[93164] = 16'b0000000000000000;
	sram_mem[93165] = 16'b0000000000000000;
	sram_mem[93166] = 16'b0000000000000000;
	sram_mem[93167] = 16'b0000000000000000;
	sram_mem[93168] = 16'b0000000000000000;
	sram_mem[93169] = 16'b0000000000000000;
	sram_mem[93170] = 16'b0000000000000000;
	sram_mem[93171] = 16'b0000000000000000;
	sram_mem[93172] = 16'b0000000000000000;
	sram_mem[93173] = 16'b0000000000000000;
	sram_mem[93174] = 16'b0000000000000000;
	sram_mem[93175] = 16'b0000000000000000;
	sram_mem[93176] = 16'b0000000000000000;
	sram_mem[93177] = 16'b0000000000000000;
	sram_mem[93178] = 16'b0000000000000000;
	sram_mem[93179] = 16'b0000000000000000;
	sram_mem[93180] = 16'b0000000000000000;
	sram_mem[93181] = 16'b0000000000000000;
	sram_mem[93182] = 16'b0000000000000000;
	sram_mem[93183] = 16'b0000000000000000;
	sram_mem[93184] = 16'b0000000000000000;
	sram_mem[93185] = 16'b0000000000000000;
	sram_mem[93186] = 16'b0000000000000000;
	sram_mem[93187] = 16'b0000000000000000;
	sram_mem[93188] = 16'b0000000000000000;
	sram_mem[93189] = 16'b0000000000000000;
	sram_mem[93190] = 16'b0000000000000000;
	sram_mem[93191] = 16'b0000000000000000;
	sram_mem[93192] = 16'b0000000000000000;
	sram_mem[93193] = 16'b0000000000000000;
	sram_mem[93194] = 16'b0000000000000000;
	sram_mem[93195] = 16'b0000000000000000;
	sram_mem[93196] = 16'b0000000000000000;
	sram_mem[93197] = 16'b0000000000000000;
	sram_mem[93198] = 16'b0000000000000000;
	sram_mem[93199] = 16'b0000000000000000;
	sram_mem[93200] = 16'b0000000000000000;
	sram_mem[93201] = 16'b0000000000000000;
	sram_mem[93202] = 16'b0000000000000000;
	sram_mem[93203] = 16'b0000000000000000;
	sram_mem[93204] = 16'b0000000000000000;
	sram_mem[93205] = 16'b0000000000000000;
	sram_mem[93206] = 16'b0000000000000000;
	sram_mem[93207] = 16'b0000000000000000;
	sram_mem[93208] = 16'b0000000000000000;
	sram_mem[93209] = 16'b0000000000000000;
	sram_mem[93210] = 16'b0000000000000000;
	sram_mem[93211] = 16'b0000000000000000;
	sram_mem[93212] = 16'b0000000000000000;
	sram_mem[93213] = 16'b0000000000000000;
	sram_mem[93214] = 16'b0000000000000000;
	sram_mem[93215] = 16'b0000000000000000;
	sram_mem[93216] = 16'b0000000000000000;
	sram_mem[93217] = 16'b0000000000000000;
	sram_mem[93218] = 16'b0000000000000000;
	sram_mem[93219] = 16'b0000000000000000;
	sram_mem[93220] = 16'b0000000000000000;
	sram_mem[93221] = 16'b0000000000000000;
	sram_mem[93222] = 16'b0000000000000000;
	sram_mem[93223] = 16'b0000000000000000;
	sram_mem[93224] = 16'b0000000000000000;
	sram_mem[93225] = 16'b0000000000000000;
	sram_mem[93226] = 16'b0000000000000000;
	sram_mem[93227] = 16'b0000000000000000;
	sram_mem[93228] = 16'b0000000000000000;
	sram_mem[93229] = 16'b0000000000000000;
	sram_mem[93230] = 16'b0000000000000000;
	sram_mem[93231] = 16'b0000000000000000;
	sram_mem[93232] = 16'b0000000000000000;
	sram_mem[93233] = 16'b0000000000000000;
	sram_mem[93234] = 16'b0000000000000000;
	sram_mem[93235] = 16'b0000000000000000;
	sram_mem[93236] = 16'b0000000000000000;
	sram_mem[93237] = 16'b0000000000000000;
	sram_mem[93238] = 16'b0000000000000000;
	sram_mem[93239] = 16'b0000000000000000;
	sram_mem[93240] = 16'b0000000000000000;
	sram_mem[93241] = 16'b0000000000000000;
	sram_mem[93242] = 16'b0000000000000000;
	sram_mem[93243] = 16'b0000000000000000;
	sram_mem[93244] = 16'b0000000000000000;
	sram_mem[93245] = 16'b0000000000000000;
	sram_mem[93246] = 16'b0000000000000000;
	sram_mem[93247] = 16'b0000000000000000;
	sram_mem[93248] = 16'b0000000000000000;
	sram_mem[93249] = 16'b0000000000000000;
	sram_mem[93250] = 16'b0000000000000000;
	sram_mem[93251] = 16'b0000000000000000;
	sram_mem[93252] = 16'b0000000000000000;
	sram_mem[93253] = 16'b0000000000000000;
	sram_mem[93254] = 16'b0000000000000000;
	sram_mem[93255] = 16'b0000000000000000;
	sram_mem[93256] = 16'b0000000000000000;
	sram_mem[93257] = 16'b0000000000000000;
	sram_mem[93258] = 16'b0000000000000000;
	sram_mem[93259] = 16'b0000000000000000;
	sram_mem[93260] = 16'b0000000000000000;
	sram_mem[93261] = 16'b0000000000000000;
	sram_mem[93262] = 16'b0000000000000000;
	sram_mem[93263] = 16'b0000000000000000;
	sram_mem[93264] = 16'b0000000000000000;
	sram_mem[93265] = 16'b0000000000000000;
	sram_mem[93266] = 16'b0000000000000000;
	sram_mem[93267] = 16'b0000000000000000;
	sram_mem[93268] = 16'b0000000000000000;
	sram_mem[93269] = 16'b0000000000000000;
	sram_mem[93270] = 16'b0000000000000000;
	sram_mem[93271] = 16'b0000000000000000;
	sram_mem[93272] = 16'b0000000000000000;
	sram_mem[93273] = 16'b0000000000000000;
	sram_mem[93274] = 16'b0000000000000000;
	sram_mem[93275] = 16'b0000000000000000;
	sram_mem[93276] = 16'b0000000000000000;
	sram_mem[93277] = 16'b0000000000000000;
	sram_mem[93278] = 16'b0000000000000000;
	sram_mem[93279] = 16'b0000000000000000;
	sram_mem[93280] = 16'b0000000000000000;
	sram_mem[93281] = 16'b0000000000000000;
	sram_mem[93282] = 16'b0000000000000000;
	sram_mem[93283] = 16'b0000000000000000;
	sram_mem[93284] = 16'b0000000000000000;
	sram_mem[93285] = 16'b0000000000000000;
	sram_mem[93286] = 16'b0000000000000000;
	sram_mem[93287] = 16'b0000000000000000;
	sram_mem[93288] = 16'b0000000000000000;
	sram_mem[93289] = 16'b0000000000000000;
	sram_mem[93290] = 16'b0000000000000000;
	sram_mem[93291] = 16'b0000000000000000;
	sram_mem[93292] = 16'b0000000000000000;
	sram_mem[93293] = 16'b0000000000000000;
	sram_mem[93294] = 16'b0000000000000000;
	sram_mem[93295] = 16'b0000000000000000;
	sram_mem[93296] = 16'b0000000000000000;
	sram_mem[93297] = 16'b0000000000000000;
	sram_mem[93298] = 16'b0000000000000000;
	sram_mem[93299] = 16'b0000000000000000;
	sram_mem[93300] = 16'b0000000000000000;
	sram_mem[93301] = 16'b0000000000000000;
	sram_mem[93302] = 16'b0000000000000000;
	sram_mem[93303] = 16'b0000000000000000;
	sram_mem[93304] = 16'b0000000000000000;
	sram_mem[93305] = 16'b0000000000000000;
	sram_mem[93306] = 16'b0000000000000000;
	sram_mem[93307] = 16'b0000000000000000;
	sram_mem[93308] = 16'b0000000000000000;
	sram_mem[93309] = 16'b0000000000000000;
	sram_mem[93310] = 16'b0000000000000000;
	sram_mem[93311] = 16'b0000000000000000;
	sram_mem[93312] = 16'b0000000000000000;
	sram_mem[93313] = 16'b0000000000000000;
	sram_mem[93314] = 16'b0000000000000000;
	sram_mem[93315] = 16'b0000000000000000;
	sram_mem[93316] = 16'b0000000000000000;
	sram_mem[93317] = 16'b0000000000000000;
	sram_mem[93318] = 16'b0000000000000000;
	sram_mem[93319] = 16'b0000000000000000;
	sram_mem[93320] = 16'b0000000000000000;
	sram_mem[93321] = 16'b0000000000000000;
	sram_mem[93322] = 16'b0000000000000000;
	sram_mem[93323] = 16'b0000000000000000;
	sram_mem[93324] = 16'b0000000000000000;
	sram_mem[93325] = 16'b0000000000000000;
	sram_mem[93326] = 16'b0000000000000000;
	sram_mem[93327] = 16'b0000000000000000;
	sram_mem[93328] = 16'b0000000000000000;
	sram_mem[93329] = 16'b0000000000000000;
	sram_mem[93330] = 16'b0000000000000000;
	sram_mem[93331] = 16'b0000000000000000;
	sram_mem[93332] = 16'b0000000000000000;
	sram_mem[93333] = 16'b0000000000000000;
	sram_mem[93334] = 16'b0000000000000000;
	sram_mem[93335] = 16'b0000000000000000;
	sram_mem[93336] = 16'b0000000000000000;
	sram_mem[93337] = 16'b0000000000000000;
	sram_mem[93338] = 16'b0000000000000000;
	sram_mem[93339] = 16'b0000000000000000;
	sram_mem[93340] = 16'b0000000000000000;
	sram_mem[93341] = 16'b0000000000000000;
	sram_mem[93342] = 16'b0000000000000000;
	sram_mem[93343] = 16'b0000000000000000;
	sram_mem[93344] = 16'b0000000000000000;
	sram_mem[93345] = 16'b0000000000000000;
	sram_mem[93346] = 16'b0000000000000000;
	sram_mem[93347] = 16'b0000000000000000;
	sram_mem[93348] = 16'b0000000000000000;
	sram_mem[93349] = 16'b0000000000000000;
	sram_mem[93350] = 16'b0000000000000000;
	sram_mem[93351] = 16'b0000000000000000;
	sram_mem[93352] = 16'b0000000000000000;
	sram_mem[93353] = 16'b0000000000000000;
	sram_mem[93354] = 16'b0000000000000000;
	sram_mem[93355] = 16'b0000000000000000;
	sram_mem[93356] = 16'b0000000000000000;
	sram_mem[93357] = 16'b0000000000000000;
	sram_mem[93358] = 16'b0000000000000000;
	sram_mem[93359] = 16'b0000000000000000;
	sram_mem[93360] = 16'b0000000000000000;
	sram_mem[93361] = 16'b0000000000000000;
	sram_mem[93362] = 16'b0000000000000000;
	sram_mem[93363] = 16'b0000000000000000;
	sram_mem[93364] = 16'b0000000000000000;
	sram_mem[93365] = 16'b0000000000000000;
	sram_mem[93366] = 16'b0000000000000000;
	sram_mem[93367] = 16'b0000000000000000;
	sram_mem[93368] = 16'b0000000000000000;
	sram_mem[93369] = 16'b0000000000000000;
	sram_mem[93370] = 16'b0000000000000000;
	sram_mem[93371] = 16'b0000000000000000;
	sram_mem[93372] = 16'b0000000000000000;
	sram_mem[93373] = 16'b0000000000000000;
	sram_mem[93374] = 16'b0000000000000000;
	sram_mem[93375] = 16'b0000000000000000;
	sram_mem[93376] = 16'b0000000000000000;
	sram_mem[93377] = 16'b0000000000000000;
	sram_mem[93378] = 16'b0000000000000000;
	sram_mem[93379] = 16'b0000000000000000;
	sram_mem[93380] = 16'b0000000000000000;
	sram_mem[93381] = 16'b0000000000000000;
	sram_mem[93382] = 16'b0000000000000000;
	sram_mem[93383] = 16'b0000000000000000;
	sram_mem[93384] = 16'b0000000000000000;
	sram_mem[93385] = 16'b0000000000000000;
	sram_mem[93386] = 16'b0000000000000000;
	sram_mem[93387] = 16'b0000000000000000;
	sram_mem[93388] = 16'b0000000000000000;
	sram_mem[93389] = 16'b0000000000000000;
	sram_mem[93390] = 16'b0000000000000000;
	sram_mem[93391] = 16'b0000000000000000;
	sram_mem[93392] = 16'b0000000000000000;
	sram_mem[93393] = 16'b0000000000000000;
	sram_mem[93394] = 16'b0000000000000000;
	sram_mem[93395] = 16'b0000000000000000;
	sram_mem[93396] = 16'b0000000000000000;
	sram_mem[93397] = 16'b0000000000000000;
	sram_mem[93398] = 16'b0000000000000000;
	sram_mem[93399] = 16'b0000000000000000;
	sram_mem[93400] = 16'b0000000000000000;
	sram_mem[93401] = 16'b0000000000000000;
	sram_mem[93402] = 16'b0000000000000000;
	sram_mem[93403] = 16'b0000000000000000;
	sram_mem[93404] = 16'b0000000000000000;
	sram_mem[93405] = 16'b0000000000000000;
	sram_mem[93406] = 16'b0000000000000000;
	sram_mem[93407] = 16'b0000000000000000;
	sram_mem[93408] = 16'b0000000000000000;
	sram_mem[93409] = 16'b0000000000000000;
	sram_mem[93410] = 16'b0000000000000000;
	sram_mem[93411] = 16'b0000000000000000;
	sram_mem[93412] = 16'b0000000000000000;
	sram_mem[93413] = 16'b0000000000000000;
	sram_mem[93414] = 16'b0000000000000000;
	sram_mem[93415] = 16'b0000000000000000;
	sram_mem[93416] = 16'b0000000000000000;
	sram_mem[93417] = 16'b0000000000000000;
	sram_mem[93418] = 16'b0000000000000000;
	sram_mem[93419] = 16'b0000000000000000;
	sram_mem[93420] = 16'b0000000000000000;
	sram_mem[93421] = 16'b0000000000000000;
	sram_mem[93422] = 16'b0000000000000000;
	sram_mem[93423] = 16'b0000000000000000;
	sram_mem[93424] = 16'b0000000000000000;
	sram_mem[93425] = 16'b0000000000000000;
	sram_mem[93426] = 16'b0000000000000000;
	sram_mem[93427] = 16'b0000000000000000;
	sram_mem[93428] = 16'b0000000000000000;
	sram_mem[93429] = 16'b0000000000000000;
	sram_mem[93430] = 16'b0000000000000000;
	sram_mem[93431] = 16'b0000000000000000;
	sram_mem[93432] = 16'b0000000000000000;
	sram_mem[93433] = 16'b0000000000000000;
	sram_mem[93434] = 16'b0000000000000000;
	sram_mem[93435] = 16'b0000000000000000;
	sram_mem[93436] = 16'b0000000000000000;
	sram_mem[93437] = 16'b0000000000000000;
	sram_mem[93438] = 16'b0000000000000000;
	sram_mem[93439] = 16'b0000000000000000;
	sram_mem[93440] = 16'b0000000000000000;
	sram_mem[93441] = 16'b0000000000000000;
	sram_mem[93442] = 16'b0000000000000000;
	sram_mem[93443] = 16'b0000000000000000;
	sram_mem[93444] = 16'b0000000000000000;
	sram_mem[93445] = 16'b0000000000000000;
	sram_mem[93446] = 16'b0000000000000000;
	sram_mem[93447] = 16'b0000000000000000;
	sram_mem[93448] = 16'b0000000000000000;
	sram_mem[93449] = 16'b0000000000000000;
	sram_mem[93450] = 16'b0000000000000000;
	sram_mem[93451] = 16'b0000000000000000;
	sram_mem[93452] = 16'b0000000000000000;
	sram_mem[93453] = 16'b0000000000000000;
	sram_mem[93454] = 16'b0000000000000000;
	sram_mem[93455] = 16'b0000000000000000;
	sram_mem[93456] = 16'b0000000000000000;
	sram_mem[93457] = 16'b0000000000000000;
	sram_mem[93458] = 16'b0000000000000000;
	sram_mem[93459] = 16'b0000000000000000;
	sram_mem[93460] = 16'b0000000000000000;
	sram_mem[93461] = 16'b0000000000000000;
	sram_mem[93462] = 16'b0000000000000000;
	sram_mem[93463] = 16'b0000000000000000;
	sram_mem[93464] = 16'b0000000000000000;
	sram_mem[93465] = 16'b0000000000000000;
	sram_mem[93466] = 16'b0000000000000000;
	sram_mem[93467] = 16'b0000000000000000;
	sram_mem[93468] = 16'b0000000000000000;
	sram_mem[93469] = 16'b0000000000000000;
	sram_mem[93470] = 16'b0000000000000000;
	sram_mem[93471] = 16'b0000000000000000;
	sram_mem[93472] = 16'b0000000000000000;
	sram_mem[93473] = 16'b0000000000000000;
	sram_mem[93474] = 16'b0000000000000000;
	sram_mem[93475] = 16'b0000000000000000;
	sram_mem[93476] = 16'b0000000000000000;
	sram_mem[93477] = 16'b0000000000000000;
	sram_mem[93478] = 16'b0000000000000000;
	sram_mem[93479] = 16'b0000000000000000;
	sram_mem[93480] = 16'b0000000000000000;
	sram_mem[93481] = 16'b0000000000000000;
	sram_mem[93482] = 16'b0000000000000000;
	sram_mem[93483] = 16'b0000000000000000;
	sram_mem[93484] = 16'b0000000000000000;
	sram_mem[93485] = 16'b0000000000000000;
	sram_mem[93486] = 16'b0000000000000000;
	sram_mem[93487] = 16'b0000000000000000;
	sram_mem[93488] = 16'b0000000000000000;
	sram_mem[93489] = 16'b0000000000000000;
	sram_mem[93490] = 16'b0000000000000000;
	sram_mem[93491] = 16'b0000000000000000;
	sram_mem[93492] = 16'b0000000000000000;
	sram_mem[93493] = 16'b0000000000000000;
	sram_mem[93494] = 16'b0000000000000000;
	sram_mem[93495] = 16'b0000000000000000;
	sram_mem[93496] = 16'b0000000000000000;
	sram_mem[93497] = 16'b0000000000000000;
	sram_mem[93498] = 16'b0000000000000000;
	sram_mem[93499] = 16'b0000000000000000;
	sram_mem[93500] = 16'b0000000000000000;
	sram_mem[93501] = 16'b0000000000000000;
	sram_mem[93502] = 16'b0000000000000000;
	sram_mem[93503] = 16'b0000000000000000;
	sram_mem[93504] = 16'b0000000000000000;
	sram_mem[93505] = 16'b0000000000000000;
	sram_mem[93506] = 16'b0000000000000000;
	sram_mem[93507] = 16'b0000000000000000;
	sram_mem[93508] = 16'b0000000000000000;
	sram_mem[93509] = 16'b0000000000000000;
	sram_mem[93510] = 16'b0000000000000000;
	sram_mem[93511] = 16'b0000000000000000;
	sram_mem[93512] = 16'b0000000000000000;
	sram_mem[93513] = 16'b0000000000000000;
	sram_mem[93514] = 16'b0000000000000000;
	sram_mem[93515] = 16'b0000000000000000;
	sram_mem[93516] = 16'b0000000000000000;
	sram_mem[93517] = 16'b0000000000000000;
	sram_mem[93518] = 16'b0000000000000000;
	sram_mem[93519] = 16'b0000000000000000;
	sram_mem[93520] = 16'b0000000000000000;
	sram_mem[93521] = 16'b0000000000000000;
	sram_mem[93522] = 16'b0000000000000000;
	sram_mem[93523] = 16'b0000000000000000;
	sram_mem[93524] = 16'b0000000000000000;
	sram_mem[93525] = 16'b0000000000000000;
	sram_mem[93526] = 16'b0000000000000000;
	sram_mem[93527] = 16'b0000000000000000;
	sram_mem[93528] = 16'b0000000000000000;
	sram_mem[93529] = 16'b0000000000000000;
	sram_mem[93530] = 16'b0000000000000000;
	sram_mem[93531] = 16'b0000000000000000;
	sram_mem[93532] = 16'b0000000000000000;
	sram_mem[93533] = 16'b0000000000000000;
	sram_mem[93534] = 16'b0000000000000000;
	sram_mem[93535] = 16'b0000000000000000;
	sram_mem[93536] = 16'b0000000000000000;
	sram_mem[93537] = 16'b0000000000000000;
	sram_mem[93538] = 16'b0000000000000000;
	sram_mem[93539] = 16'b0000000000000000;
	sram_mem[93540] = 16'b0000000000000000;
	sram_mem[93541] = 16'b0000000000000000;
	sram_mem[93542] = 16'b0000000000000000;
	sram_mem[93543] = 16'b0000000000000000;
	sram_mem[93544] = 16'b0000000000000000;
	sram_mem[93545] = 16'b0000000000000000;
	sram_mem[93546] = 16'b0000000000000000;
	sram_mem[93547] = 16'b0000000000000000;
	sram_mem[93548] = 16'b0000000000000000;
	sram_mem[93549] = 16'b0000000000000000;
	sram_mem[93550] = 16'b0000000000000000;
	sram_mem[93551] = 16'b0000000000000000;
	sram_mem[93552] = 16'b0000000000000000;
	sram_mem[93553] = 16'b0000000000000000;
	sram_mem[93554] = 16'b0000000000000000;
	sram_mem[93555] = 16'b0000000000000000;
	sram_mem[93556] = 16'b0000000000000000;
	sram_mem[93557] = 16'b0000000000000000;
	sram_mem[93558] = 16'b0000000000000000;
	sram_mem[93559] = 16'b0000000000000000;
	sram_mem[93560] = 16'b0000000000000000;
	sram_mem[93561] = 16'b0000000000000000;
	sram_mem[93562] = 16'b0000000000000000;
	sram_mem[93563] = 16'b0000000000000000;
	sram_mem[93564] = 16'b0000000000000000;
	sram_mem[93565] = 16'b0000000000000000;
	sram_mem[93566] = 16'b0000000000000000;
	sram_mem[93567] = 16'b0000000000000000;
	sram_mem[93568] = 16'b0000000000000000;
	sram_mem[93569] = 16'b0000000000000000;
	sram_mem[93570] = 16'b0000000000000000;
	sram_mem[93571] = 16'b0000000000000000;
	sram_mem[93572] = 16'b0000000000000000;
	sram_mem[93573] = 16'b0000000000000000;
	sram_mem[93574] = 16'b0000000000000000;
	sram_mem[93575] = 16'b0000000000000000;
	sram_mem[93576] = 16'b0000000000000000;
	sram_mem[93577] = 16'b0000000000000000;
	sram_mem[93578] = 16'b0000000000000000;
	sram_mem[93579] = 16'b0000000000000000;
	sram_mem[93580] = 16'b0000000000000000;
	sram_mem[93581] = 16'b0000000000000000;
	sram_mem[93582] = 16'b0000000000000000;
	sram_mem[93583] = 16'b0000000000000000;
	sram_mem[93584] = 16'b0000000000000000;
	sram_mem[93585] = 16'b0000000000000000;
	sram_mem[93586] = 16'b0000000000000000;
	sram_mem[93587] = 16'b0000000000000000;
	sram_mem[93588] = 16'b0000000000000000;
	sram_mem[93589] = 16'b0000000000000000;
	sram_mem[93590] = 16'b0000000000000000;
	sram_mem[93591] = 16'b0000000000000000;
	sram_mem[93592] = 16'b0000000000000000;
	sram_mem[93593] = 16'b0000000000000000;
	sram_mem[93594] = 16'b0000000000000000;
	sram_mem[93595] = 16'b0000000000000000;
	sram_mem[93596] = 16'b0000000000000000;
	sram_mem[93597] = 16'b0000000000000000;
	sram_mem[93598] = 16'b0000000000000000;
	sram_mem[93599] = 16'b0000000000000000;
	sram_mem[93600] = 16'b0000000000000000;
	sram_mem[93601] = 16'b0000000000000000;
	sram_mem[93602] = 16'b0000000000000000;
	sram_mem[93603] = 16'b0000000000000000;
	sram_mem[93604] = 16'b0000000000000000;
	sram_mem[93605] = 16'b0000000000000000;
	sram_mem[93606] = 16'b0000000000000000;
	sram_mem[93607] = 16'b0000000000000000;
	sram_mem[93608] = 16'b0000000000000000;
	sram_mem[93609] = 16'b0000000000000000;
	sram_mem[93610] = 16'b0000000000000000;
	sram_mem[93611] = 16'b0000000000000000;
	sram_mem[93612] = 16'b0000000000000000;
	sram_mem[93613] = 16'b0000000000000000;
	sram_mem[93614] = 16'b0000000000000000;
	sram_mem[93615] = 16'b0000000000000000;
	sram_mem[93616] = 16'b0000000000000000;
	sram_mem[93617] = 16'b0000000000000000;
	sram_mem[93618] = 16'b0000000000000000;
	sram_mem[93619] = 16'b0000000000000000;
	sram_mem[93620] = 16'b0000000000000000;
	sram_mem[93621] = 16'b0000000000000000;
	sram_mem[93622] = 16'b0000000000000000;
	sram_mem[93623] = 16'b0000000000000000;
	sram_mem[93624] = 16'b0000000000000000;
	sram_mem[93625] = 16'b0000000000000000;
	sram_mem[93626] = 16'b0000000000000000;
	sram_mem[93627] = 16'b0000000000000000;
	sram_mem[93628] = 16'b0000000000000000;
	sram_mem[93629] = 16'b0000000000000000;
	sram_mem[93630] = 16'b0000000000000000;
	sram_mem[93631] = 16'b0000000000000000;
	sram_mem[93632] = 16'b0000000000000000;
	sram_mem[93633] = 16'b0000000000000000;
	sram_mem[93634] = 16'b0000000000000000;
	sram_mem[93635] = 16'b0000000000000000;
	sram_mem[93636] = 16'b0000000000000000;
	sram_mem[93637] = 16'b0000000000000000;
	sram_mem[93638] = 16'b0000000000000000;
	sram_mem[93639] = 16'b0000000000000000;
	sram_mem[93640] = 16'b0000000000000000;
	sram_mem[93641] = 16'b0000000000000000;
	sram_mem[93642] = 16'b0000000000000000;
	sram_mem[93643] = 16'b0000000000000000;
	sram_mem[93644] = 16'b0000000000000000;
	sram_mem[93645] = 16'b0000000000000000;
	sram_mem[93646] = 16'b0000000000000000;
	sram_mem[93647] = 16'b0000000000000000;
	sram_mem[93648] = 16'b0000000000000000;
	sram_mem[93649] = 16'b0000000000000000;
	sram_mem[93650] = 16'b0000000000000000;
	sram_mem[93651] = 16'b0000000000000000;
	sram_mem[93652] = 16'b0000000000000000;
	sram_mem[93653] = 16'b0000000000000000;
	sram_mem[93654] = 16'b0000000000000000;
	sram_mem[93655] = 16'b0000000000000000;
	sram_mem[93656] = 16'b0000000000000000;
	sram_mem[93657] = 16'b0000000000000000;
	sram_mem[93658] = 16'b0000000000000000;
	sram_mem[93659] = 16'b0000000000000000;
	sram_mem[93660] = 16'b0000000000000000;
	sram_mem[93661] = 16'b0000000000000000;
	sram_mem[93662] = 16'b0000000000000000;
	sram_mem[93663] = 16'b0000000000000000;
	sram_mem[93664] = 16'b0000000000000000;
	sram_mem[93665] = 16'b0000000000000000;
	sram_mem[93666] = 16'b0000000000000000;
	sram_mem[93667] = 16'b0000000000000000;
	sram_mem[93668] = 16'b0000000000000000;
	sram_mem[93669] = 16'b0000000000000000;
	sram_mem[93670] = 16'b0000000000000000;
	sram_mem[93671] = 16'b0000000000000000;
	sram_mem[93672] = 16'b0000000000000000;
	sram_mem[93673] = 16'b0000000000000000;
	sram_mem[93674] = 16'b0000000000000000;
	sram_mem[93675] = 16'b0000000000000000;
	sram_mem[93676] = 16'b0000000000000000;
	sram_mem[93677] = 16'b0000000000000000;
	sram_mem[93678] = 16'b0000000000000000;
	sram_mem[93679] = 16'b0000000000000000;
	sram_mem[93680] = 16'b0000000000000000;
	sram_mem[93681] = 16'b0000000000000000;
	sram_mem[93682] = 16'b0000000000000000;
	sram_mem[93683] = 16'b0000000000000000;
	sram_mem[93684] = 16'b0000000000000000;
	sram_mem[93685] = 16'b0000000000000000;
	sram_mem[93686] = 16'b0000000000000000;
	sram_mem[93687] = 16'b0000000000000000;
	sram_mem[93688] = 16'b0000000000000000;
	sram_mem[93689] = 16'b0000000000000000;
	sram_mem[93690] = 16'b0000000000000000;
	sram_mem[93691] = 16'b0000000000000000;
	sram_mem[93692] = 16'b0000000000000000;
	sram_mem[93693] = 16'b0000000000000000;
	sram_mem[93694] = 16'b0000000000000000;
	sram_mem[93695] = 16'b0000000000000000;
	sram_mem[93696] = 16'b0000000000000000;
	sram_mem[93697] = 16'b0000000000000000;
	sram_mem[93698] = 16'b0000000000000000;
	sram_mem[93699] = 16'b0000000000000000;
	sram_mem[93700] = 16'b0000000000000000;
	sram_mem[93701] = 16'b0000000000000000;
	sram_mem[93702] = 16'b0000000000000000;
	sram_mem[93703] = 16'b0000000000000000;
	sram_mem[93704] = 16'b0000000000000000;
	sram_mem[93705] = 16'b0000000000000000;
	sram_mem[93706] = 16'b0000000000000000;
	sram_mem[93707] = 16'b0000000000000000;
	sram_mem[93708] = 16'b0000000000000000;
	sram_mem[93709] = 16'b0000000000000000;
	sram_mem[93710] = 16'b0000000000000000;
	sram_mem[93711] = 16'b0000000000000000;
	sram_mem[93712] = 16'b0000000000000000;
	sram_mem[93713] = 16'b0000000000000000;
	sram_mem[93714] = 16'b0000000000000000;
	sram_mem[93715] = 16'b0000000000000000;
	sram_mem[93716] = 16'b0000000000000000;
	sram_mem[93717] = 16'b0000000000000000;
	sram_mem[93718] = 16'b0000000000000000;
	sram_mem[93719] = 16'b0000000000000000;
	sram_mem[93720] = 16'b0000000000000000;
	sram_mem[93721] = 16'b0000000000000000;
	sram_mem[93722] = 16'b0000000000000000;
	sram_mem[93723] = 16'b0000000000000000;
	sram_mem[93724] = 16'b0000000000000000;
	sram_mem[93725] = 16'b0000000000000000;
	sram_mem[93726] = 16'b0000000000000000;
	sram_mem[93727] = 16'b0000000000000000;
	sram_mem[93728] = 16'b0000000000000000;
	sram_mem[93729] = 16'b0000000000000000;
	sram_mem[93730] = 16'b0000000000000000;
	sram_mem[93731] = 16'b0000000000000000;
	sram_mem[93732] = 16'b0000000000000000;
	sram_mem[93733] = 16'b0000000000000000;
	sram_mem[93734] = 16'b0000000000000000;
	sram_mem[93735] = 16'b0000000000000000;
	sram_mem[93736] = 16'b0000000000000000;
	sram_mem[93737] = 16'b0000000000000000;
	sram_mem[93738] = 16'b0000000000000000;
	sram_mem[93739] = 16'b0000000000000000;
	sram_mem[93740] = 16'b0000000000000000;
	sram_mem[93741] = 16'b0000000000000000;
	sram_mem[93742] = 16'b0000000000000000;
	sram_mem[93743] = 16'b0000000000000000;
	sram_mem[93744] = 16'b0000000000000000;
	sram_mem[93745] = 16'b0000000000000000;
	sram_mem[93746] = 16'b0000000000000000;
	sram_mem[93747] = 16'b0000000000000000;
	sram_mem[93748] = 16'b0000000000000000;
	sram_mem[93749] = 16'b0000000000000000;
	sram_mem[93750] = 16'b0000000000000000;
	sram_mem[93751] = 16'b0000000000000000;
	sram_mem[93752] = 16'b0000000000000000;
	sram_mem[93753] = 16'b0000000000000000;
	sram_mem[93754] = 16'b0000000000000000;
	sram_mem[93755] = 16'b0000000000000000;
	sram_mem[93756] = 16'b0000000000000000;
	sram_mem[93757] = 16'b0000000000000000;
	sram_mem[93758] = 16'b0000000000000000;
	sram_mem[93759] = 16'b0000000000000000;
	sram_mem[93760] = 16'b0000000000000000;
	sram_mem[93761] = 16'b0000000000000000;
	sram_mem[93762] = 16'b0000000000000000;
	sram_mem[93763] = 16'b0000000000000000;
	sram_mem[93764] = 16'b0000000000000000;
	sram_mem[93765] = 16'b0000000000000000;
	sram_mem[93766] = 16'b0000000000000000;
	sram_mem[93767] = 16'b0000000000000000;
	sram_mem[93768] = 16'b0000000000000000;
	sram_mem[93769] = 16'b0000000000000000;
	sram_mem[93770] = 16'b0000000000000000;
	sram_mem[93771] = 16'b0000000000000000;
	sram_mem[93772] = 16'b0000000000000000;
	sram_mem[93773] = 16'b0000000000000000;
	sram_mem[93774] = 16'b0000000000000000;
	sram_mem[93775] = 16'b0000000000000000;
	sram_mem[93776] = 16'b0000000000000000;
	sram_mem[93777] = 16'b0000000000000000;
	sram_mem[93778] = 16'b0000000000000000;
	sram_mem[93779] = 16'b0000000000000000;
	sram_mem[93780] = 16'b0000000000000000;
	sram_mem[93781] = 16'b0000000000000000;
	sram_mem[93782] = 16'b0000000000000000;
	sram_mem[93783] = 16'b0000000000000000;
	sram_mem[93784] = 16'b0000000000000000;
	sram_mem[93785] = 16'b0000000000000000;
	sram_mem[93786] = 16'b0000000000000000;
	sram_mem[93787] = 16'b0000000000000000;
	sram_mem[93788] = 16'b0000000000000000;
	sram_mem[93789] = 16'b0000000000000000;
	sram_mem[93790] = 16'b0000000000000000;
	sram_mem[93791] = 16'b0000000000000000;
	sram_mem[93792] = 16'b0000000000000000;
	sram_mem[93793] = 16'b0000000000000000;
	sram_mem[93794] = 16'b0000000000000000;
	sram_mem[93795] = 16'b0000000000000000;
	sram_mem[93796] = 16'b0000000000000000;
	sram_mem[93797] = 16'b0000000000000000;
	sram_mem[93798] = 16'b0000000000000000;
	sram_mem[93799] = 16'b0000000000000000;
	sram_mem[93800] = 16'b0000000000000000;
	sram_mem[93801] = 16'b0000000000000000;
	sram_mem[93802] = 16'b0000000000000000;
	sram_mem[93803] = 16'b0000000000000000;
	sram_mem[93804] = 16'b0000000000000000;
	sram_mem[93805] = 16'b0000000000000000;
	sram_mem[93806] = 16'b0000000000000000;
	sram_mem[93807] = 16'b0000000000000000;
	sram_mem[93808] = 16'b0000000000000000;
	sram_mem[93809] = 16'b0000000000000000;
	sram_mem[93810] = 16'b0000000000000000;
	sram_mem[93811] = 16'b0000000000000000;
	sram_mem[93812] = 16'b0000000000000000;
	sram_mem[93813] = 16'b0000000000000000;
	sram_mem[93814] = 16'b0000000000000000;
	sram_mem[93815] = 16'b0000000000000000;
	sram_mem[93816] = 16'b0000000000000000;
	sram_mem[93817] = 16'b0000000000000000;
	sram_mem[93818] = 16'b0000000000000000;
	sram_mem[93819] = 16'b0000000000000000;
	sram_mem[93820] = 16'b0000000000000000;
	sram_mem[93821] = 16'b0000000000000000;
	sram_mem[93822] = 16'b0000000000000000;
	sram_mem[93823] = 16'b0000000000000000;
	sram_mem[93824] = 16'b0000000000000000;
	sram_mem[93825] = 16'b0000000000000000;
	sram_mem[93826] = 16'b0000000000000000;
	sram_mem[93827] = 16'b0000000000000000;
	sram_mem[93828] = 16'b0000000000000000;
	sram_mem[93829] = 16'b0000000000000000;
	sram_mem[93830] = 16'b0000000000000000;
	sram_mem[93831] = 16'b0000000000000000;
	sram_mem[93832] = 16'b0000000000000000;
	sram_mem[93833] = 16'b0000000000000000;
	sram_mem[93834] = 16'b0000000000000000;
	sram_mem[93835] = 16'b0000000000000000;
	sram_mem[93836] = 16'b0000000000000000;
	sram_mem[93837] = 16'b0000000000000000;
	sram_mem[93838] = 16'b0000000000000000;
	sram_mem[93839] = 16'b0000000000000000;
	sram_mem[93840] = 16'b0000000000000000;
	sram_mem[93841] = 16'b0000000000000000;
	sram_mem[93842] = 16'b0000000000000000;
	sram_mem[93843] = 16'b0000000000000000;
	sram_mem[93844] = 16'b0000000000000000;
	sram_mem[93845] = 16'b0000000000000000;
	sram_mem[93846] = 16'b0000000000000000;
	sram_mem[93847] = 16'b0000000000000000;
	sram_mem[93848] = 16'b0000000000000000;
	sram_mem[93849] = 16'b0000000000000000;
	sram_mem[93850] = 16'b0000000000000000;
	sram_mem[93851] = 16'b0000000000000000;
	sram_mem[93852] = 16'b0000000000000000;
	sram_mem[93853] = 16'b0000000000000000;
	sram_mem[93854] = 16'b0000000000000000;
	sram_mem[93855] = 16'b0000000000000000;
	sram_mem[93856] = 16'b0000000000000000;
	sram_mem[93857] = 16'b0000000000000000;
	sram_mem[93858] = 16'b0000000000000000;
	sram_mem[93859] = 16'b0000000000000000;
	sram_mem[93860] = 16'b0000000000000000;
	sram_mem[93861] = 16'b0000000000000000;
	sram_mem[93862] = 16'b0000000000000000;
	sram_mem[93863] = 16'b0000000000000000;
	sram_mem[93864] = 16'b0000000000000000;
	sram_mem[93865] = 16'b0000000000000000;
	sram_mem[93866] = 16'b0000000000000000;
	sram_mem[93867] = 16'b0000000000000000;
	sram_mem[93868] = 16'b0000000000000000;
	sram_mem[93869] = 16'b0000000000000000;
	sram_mem[93870] = 16'b0000000000000000;
	sram_mem[93871] = 16'b0000000000000000;
	sram_mem[93872] = 16'b0000000000000000;
	sram_mem[93873] = 16'b0000000000000000;
	sram_mem[93874] = 16'b0000000000000000;
	sram_mem[93875] = 16'b0000000000000000;
	sram_mem[93876] = 16'b0000000000000000;
	sram_mem[93877] = 16'b0000000000000000;
	sram_mem[93878] = 16'b0000000000000000;
	sram_mem[93879] = 16'b0000000000000000;
	sram_mem[93880] = 16'b0000000000000000;
	sram_mem[93881] = 16'b0000000000000000;
	sram_mem[93882] = 16'b0000000000000000;
	sram_mem[93883] = 16'b0000000000000000;
	sram_mem[93884] = 16'b0000000000000000;
	sram_mem[93885] = 16'b0000000000000000;
	sram_mem[93886] = 16'b0000000000000000;
	sram_mem[93887] = 16'b0000000000000000;
	sram_mem[93888] = 16'b0000000000000000;
	sram_mem[93889] = 16'b0000000000000000;
	sram_mem[93890] = 16'b0000000000000000;
	sram_mem[93891] = 16'b0000000000000000;
	sram_mem[93892] = 16'b0000000000000000;
	sram_mem[93893] = 16'b0000000000000000;
	sram_mem[93894] = 16'b0000000000000000;
	sram_mem[93895] = 16'b0000000000000000;
	sram_mem[93896] = 16'b0000000000000000;
	sram_mem[93897] = 16'b0000000000000000;
	sram_mem[93898] = 16'b0000000000000000;
	sram_mem[93899] = 16'b0000000000000000;
	sram_mem[93900] = 16'b0000000000000000;
	sram_mem[93901] = 16'b0000000000000000;
	sram_mem[93902] = 16'b0000000000000000;
	sram_mem[93903] = 16'b0000000000000000;
	sram_mem[93904] = 16'b0000000000000000;
	sram_mem[93905] = 16'b0000000000000000;
	sram_mem[93906] = 16'b0000000000000000;
	sram_mem[93907] = 16'b0000000000000000;
	sram_mem[93908] = 16'b0000000000000000;
	sram_mem[93909] = 16'b0000000000000000;
	sram_mem[93910] = 16'b0000000000000000;
	sram_mem[93911] = 16'b0000000000000000;
	sram_mem[93912] = 16'b0000000000000000;
	sram_mem[93913] = 16'b0000000000000000;
	sram_mem[93914] = 16'b0000000000000000;
	sram_mem[93915] = 16'b0000000000000000;
	sram_mem[93916] = 16'b0000000000000000;
	sram_mem[93917] = 16'b0000000000000000;
	sram_mem[93918] = 16'b0000000000000000;
	sram_mem[93919] = 16'b0000000000000000;
	sram_mem[93920] = 16'b0000000000000000;
	sram_mem[93921] = 16'b0000000000000000;
	sram_mem[93922] = 16'b0000000000000000;
	sram_mem[93923] = 16'b0000000000000000;
	sram_mem[93924] = 16'b0000000000000000;
	sram_mem[93925] = 16'b0000000000000000;
	sram_mem[93926] = 16'b0000000000000000;
	sram_mem[93927] = 16'b0000000000000000;
	sram_mem[93928] = 16'b0000000000000000;
	sram_mem[93929] = 16'b0000000000000000;
	sram_mem[93930] = 16'b0000000000000000;
	sram_mem[93931] = 16'b0000000000000000;
	sram_mem[93932] = 16'b0000000000000000;
	sram_mem[93933] = 16'b0000000000000000;
	sram_mem[93934] = 16'b0000000000000000;
	sram_mem[93935] = 16'b0000000000000000;
	sram_mem[93936] = 16'b0000000000000000;
	sram_mem[93937] = 16'b0000000000000000;
	sram_mem[93938] = 16'b0000000000000000;
	sram_mem[93939] = 16'b0000000000000000;
	sram_mem[93940] = 16'b0000000000000000;
	sram_mem[93941] = 16'b0000000000000000;
	sram_mem[93942] = 16'b0000000000000000;
	sram_mem[93943] = 16'b0000000000000000;
	sram_mem[93944] = 16'b0000000000000000;
	sram_mem[93945] = 16'b0000000000000000;
	sram_mem[93946] = 16'b0000000000000000;
	sram_mem[93947] = 16'b0000000000000000;
	sram_mem[93948] = 16'b0000000000000000;
	sram_mem[93949] = 16'b0000000000000000;
	sram_mem[93950] = 16'b0000000000000000;
	sram_mem[93951] = 16'b0000000000000000;
	sram_mem[93952] = 16'b0000000000000000;
	sram_mem[93953] = 16'b0000000000000000;
	sram_mem[93954] = 16'b0000000000000000;
	sram_mem[93955] = 16'b0000000000000000;
	sram_mem[93956] = 16'b0000000000000000;
	sram_mem[93957] = 16'b0000000000000000;
	sram_mem[93958] = 16'b0000000000000000;
	sram_mem[93959] = 16'b0000000000000000;
	sram_mem[93960] = 16'b0000000000000000;
	sram_mem[93961] = 16'b0000000000000000;
	sram_mem[93962] = 16'b0000000000000000;
	sram_mem[93963] = 16'b0000000000000000;
	sram_mem[93964] = 16'b0000000000000000;
	sram_mem[93965] = 16'b0000000000000000;
	sram_mem[93966] = 16'b0000000000000000;
	sram_mem[93967] = 16'b0000000000000000;
	sram_mem[93968] = 16'b0000000000000000;
	sram_mem[93969] = 16'b0000000000000000;
	sram_mem[93970] = 16'b0000000000000000;
	sram_mem[93971] = 16'b0000000000000000;
	sram_mem[93972] = 16'b0000000000000000;
	sram_mem[93973] = 16'b0000000000000000;
	sram_mem[93974] = 16'b0000000000000000;
	sram_mem[93975] = 16'b0000000000000000;
	sram_mem[93976] = 16'b0000000000000000;
	sram_mem[93977] = 16'b0000000000000000;
	sram_mem[93978] = 16'b0000000000000000;
	sram_mem[93979] = 16'b0000000000000000;
	sram_mem[93980] = 16'b0000000000000000;
	sram_mem[93981] = 16'b0000000000000000;
	sram_mem[93982] = 16'b0000000000000000;
	sram_mem[93983] = 16'b0000000000000000;
	sram_mem[93984] = 16'b0000000000000000;
	sram_mem[93985] = 16'b0000000000000000;
	sram_mem[93986] = 16'b0000000000000000;
	sram_mem[93987] = 16'b0000000000000000;
	sram_mem[93988] = 16'b0000000000000000;
	sram_mem[93989] = 16'b0000000000000000;
	sram_mem[93990] = 16'b0000000000000000;
	sram_mem[93991] = 16'b0000000000000000;
	sram_mem[93992] = 16'b0000000000000000;
	sram_mem[93993] = 16'b0000000000000000;
	sram_mem[93994] = 16'b0000000000000000;
	sram_mem[93995] = 16'b0000000000000000;
	sram_mem[93996] = 16'b0000000000000000;
	sram_mem[93997] = 16'b0000000000000000;
	sram_mem[93998] = 16'b0000000000000000;
	sram_mem[93999] = 16'b0000000000000000;
	sram_mem[94000] = 16'b0000000000000000;
	sram_mem[94001] = 16'b0000000000000000;
	sram_mem[94002] = 16'b0000000000000000;
	sram_mem[94003] = 16'b0000000000000000;
	sram_mem[94004] = 16'b0000000000000000;
	sram_mem[94005] = 16'b0000000000000000;
	sram_mem[94006] = 16'b0000000000000000;
	sram_mem[94007] = 16'b0000000000000000;
	sram_mem[94008] = 16'b0000000000000000;
	sram_mem[94009] = 16'b0000000000000000;
	sram_mem[94010] = 16'b0000000000000000;
	sram_mem[94011] = 16'b0000000000000000;
	sram_mem[94012] = 16'b0000000000000000;
	sram_mem[94013] = 16'b0000000000000000;
	sram_mem[94014] = 16'b0000000000000000;
	sram_mem[94015] = 16'b0000000000000000;
	sram_mem[94016] = 16'b0000000000000000;
	sram_mem[94017] = 16'b0000000000000000;
	sram_mem[94018] = 16'b0000000000000000;
	sram_mem[94019] = 16'b0000000000000000;
	sram_mem[94020] = 16'b0000000000000000;
	sram_mem[94021] = 16'b0000000000000000;
	sram_mem[94022] = 16'b0000000000000000;
	sram_mem[94023] = 16'b0000000000000000;
	sram_mem[94024] = 16'b0000000000000000;
	sram_mem[94025] = 16'b0000000000000000;
	sram_mem[94026] = 16'b0000000000000000;
	sram_mem[94027] = 16'b0000000000000000;
	sram_mem[94028] = 16'b0000000000000000;
	sram_mem[94029] = 16'b0000000000000000;
	sram_mem[94030] = 16'b0000000000000000;
	sram_mem[94031] = 16'b0000000000000000;
	sram_mem[94032] = 16'b0000000000000000;
	sram_mem[94033] = 16'b0000000000000000;
	sram_mem[94034] = 16'b0000000000000000;
	sram_mem[94035] = 16'b0000000000000000;
	sram_mem[94036] = 16'b0000000000000000;
	sram_mem[94037] = 16'b0000000000000000;
	sram_mem[94038] = 16'b0000000000000000;
	sram_mem[94039] = 16'b0000000000000000;
	sram_mem[94040] = 16'b0000000000000000;
	sram_mem[94041] = 16'b0000000000000000;
	sram_mem[94042] = 16'b0000000000000000;
	sram_mem[94043] = 16'b0000000000000000;
	sram_mem[94044] = 16'b0000000000000000;
	sram_mem[94045] = 16'b0000000000000000;
	sram_mem[94046] = 16'b0000000000000000;
	sram_mem[94047] = 16'b0000000000000000;
	sram_mem[94048] = 16'b0000000000000000;
	sram_mem[94049] = 16'b0000000000000000;
	sram_mem[94050] = 16'b0000000000000000;
	sram_mem[94051] = 16'b0000000000000000;
	sram_mem[94052] = 16'b0000000000000000;
	sram_mem[94053] = 16'b0000000000000000;
	sram_mem[94054] = 16'b0000000000000000;
	sram_mem[94055] = 16'b0000000000000000;
	sram_mem[94056] = 16'b0000000000000000;
	sram_mem[94057] = 16'b0000000000000000;
	sram_mem[94058] = 16'b0000000000000000;
	sram_mem[94059] = 16'b0000000000000000;
	sram_mem[94060] = 16'b0000000000000000;
	sram_mem[94061] = 16'b0000000000000000;
	sram_mem[94062] = 16'b0000000000000000;
	sram_mem[94063] = 16'b0000000000000000;
	sram_mem[94064] = 16'b0000000000000000;
	sram_mem[94065] = 16'b0000000000000000;
	sram_mem[94066] = 16'b0000000000000000;
	sram_mem[94067] = 16'b0000000000000000;
	sram_mem[94068] = 16'b0000000000000000;
	sram_mem[94069] = 16'b0000000000000000;
	sram_mem[94070] = 16'b0000000000000000;
	sram_mem[94071] = 16'b0000000000000000;
	sram_mem[94072] = 16'b0000000000000000;
	sram_mem[94073] = 16'b0000000000000000;
	sram_mem[94074] = 16'b0000000000000000;
	sram_mem[94075] = 16'b0000000000000000;
	sram_mem[94076] = 16'b0000000000000000;
	sram_mem[94077] = 16'b0000000000000000;
	sram_mem[94078] = 16'b0000000000000000;
	sram_mem[94079] = 16'b0000000000000000;
	sram_mem[94080] = 16'b0000000000000000;
	sram_mem[94081] = 16'b0000000000000000;
	sram_mem[94082] = 16'b0000000000000000;
	sram_mem[94083] = 16'b0000000000000000;
	sram_mem[94084] = 16'b0000000000000000;
	sram_mem[94085] = 16'b0000000000000000;
	sram_mem[94086] = 16'b0000000000000000;
	sram_mem[94087] = 16'b0000000000000000;
	sram_mem[94088] = 16'b0000000000000000;
	sram_mem[94089] = 16'b0000000000000000;
	sram_mem[94090] = 16'b0000000000000000;
	sram_mem[94091] = 16'b0000000000000000;
	sram_mem[94092] = 16'b0000000000000000;
	sram_mem[94093] = 16'b0000000000000000;
	sram_mem[94094] = 16'b0000000000000000;
	sram_mem[94095] = 16'b0000000000000000;
	sram_mem[94096] = 16'b0000000000000000;
	sram_mem[94097] = 16'b0000000000000000;
	sram_mem[94098] = 16'b0000000000000000;
	sram_mem[94099] = 16'b0000000000000000;
	sram_mem[94100] = 16'b0000000000000000;
	sram_mem[94101] = 16'b0000000000000000;
	sram_mem[94102] = 16'b0000000000000000;
	sram_mem[94103] = 16'b0000000000000000;
	sram_mem[94104] = 16'b0000000000000000;
	sram_mem[94105] = 16'b0000000000000000;
	sram_mem[94106] = 16'b0000000000000000;
	sram_mem[94107] = 16'b0000000000000000;
	sram_mem[94108] = 16'b0000000000000000;
	sram_mem[94109] = 16'b0000000000000000;
	sram_mem[94110] = 16'b0000000000000000;
	sram_mem[94111] = 16'b0000000000000000;
	sram_mem[94112] = 16'b0000000000000000;
	sram_mem[94113] = 16'b0000000000000000;
	sram_mem[94114] = 16'b0000000000000000;
	sram_mem[94115] = 16'b0000000000000000;
	sram_mem[94116] = 16'b0000000000000000;
	sram_mem[94117] = 16'b0000000000000000;
	sram_mem[94118] = 16'b0000000000000000;
	sram_mem[94119] = 16'b0000000000000000;
	sram_mem[94120] = 16'b0000000000000000;
	sram_mem[94121] = 16'b0000000000000000;
	sram_mem[94122] = 16'b0000000000000000;
	sram_mem[94123] = 16'b0000000000000000;
	sram_mem[94124] = 16'b0000000000000000;
	sram_mem[94125] = 16'b0000000000000000;
	sram_mem[94126] = 16'b0000000000000000;
	sram_mem[94127] = 16'b0000000000000000;
	sram_mem[94128] = 16'b0000000000000000;
	sram_mem[94129] = 16'b0000000000000000;
	sram_mem[94130] = 16'b0000000000000000;
	sram_mem[94131] = 16'b0000000000000000;
	sram_mem[94132] = 16'b0000000000000000;
	sram_mem[94133] = 16'b0000000000000000;
	sram_mem[94134] = 16'b0000000000000000;
	sram_mem[94135] = 16'b0000000000000000;
	sram_mem[94136] = 16'b0000000000000000;
	sram_mem[94137] = 16'b0000000000000000;
	sram_mem[94138] = 16'b0000000000000000;
	sram_mem[94139] = 16'b0000000000000000;
	sram_mem[94140] = 16'b0000000000000000;
	sram_mem[94141] = 16'b0000000000000000;
	sram_mem[94142] = 16'b0000000000000000;
	sram_mem[94143] = 16'b0000000000000000;
	sram_mem[94144] = 16'b0000000000000000;
	sram_mem[94145] = 16'b0000000000000000;
	sram_mem[94146] = 16'b0000000000000000;
	sram_mem[94147] = 16'b0000000000000000;
	sram_mem[94148] = 16'b0000000000000000;
	sram_mem[94149] = 16'b0000000000000000;
	sram_mem[94150] = 16'b0000000000000000;
	sram_mem[94151] = 16'b0000000000000000;
	sram_mem[94152] = 16'b0000000000000000;
	sram_mem[94153] = 16'b0000000000000000;
	sram_mem[94154] = 16'b0000000000000000;
	sram_mem[94155] = 16'b0000000000000000;
	sram_mem[94156] = 16'b0000000000000000;
	sram_mem[94157] = 16'b0000000000000000;
	sram_mem[94158] = 16'b0000000000000000;
	sram_mem[94159] = 16'b0000000000000000;
	sram_mem[94160] = 16'b0000000000000000;
	sram_mem[94161] = 16'b0000000000000000;
	sram_mem[94162] = 16'b0000000000000000;
	sram_mem[94163] = 16'b0000000000000000;
	sram_mem[94164] = 16'b0000000000000000;
	sram_mem[94165] = 16'b0000000000000000;
	sram_mem[94166] = 16'b0000000000000000;
	sram_mem[94167] = 16'b0000000000000000;
	sram_mem[94168] = 16'b0000000000000000;
	sram_mem[94169] = 16'b0000000000000000;
	sram_mem[94170] = 16'b0000000000000000;
	sram_mem[94171] = 16'b0000000000000000;
	sram_mem[94172] = 16'b0000000000000000;
	sram_mem[94173] = 16'b0000000000000000;
	sram_mem[94174] = 16'b0000000000000000;
	sram_mem[94175] = 16'b0000000000000000;
	sram_mem[94176] = 16'b0000000000000000;
	sram_mem[94177] = 16'b0000000000000000;
	sram_mem[94178] = 16'b0000000000000000;
	sram_mem[94179] = 16'b0000000000000000;
	sram_mem[94180] = 16'b0000000000000000;
	sram_mem[94181] = 16'b0000000000000000;
	sram_mem[94182] = 16'b0000000000000000;
	sram_mem[94183] = 16'b0000000000000000;
	sram_mem[94184] = 16'b0000000000000000;
	sram_mem[94185] = 16'b0000000000000000;
	sram_mem[94186] = 16'b0000000000000000;
	sram_mem[94187] = 16'b0000000000000000;
	sram_mem[94188] = 16'b0000000000000000;
	sram_mem[94189] = 16'b0000000000000000;
	sram_mem[94190] = 16'b0000000000000000;
	sram_mem[94191] = 16'b0000000000000000;
	sram_mem[94192] = 16'b0000000000000000;
	sram_mem[94193] = 16'b0000000000000000;
	sram_mem[94194] = 16'b0000000000000000;
	sram_mem[94195] = 16'b0000000000000000;
	sram_mem[94196] = 16'b0000000000000000;
	sram_mem[94197] = 16'b0000000000000000;
	sram_mem[94198] = 16'b0000000000000000;
	sram_mem[94199] = 16'b0000000000000000;
	sram_mem[94200] = 16'b0000000000000000;
	sram_mem[94201] = 16'b0000000000000000;
	sram_mem[94202] = 16'b0000000000000000;
	sram_mem[94203] = 16'b0000000000000000;
	sram_mem[94204] = 16'b0000000000000000;
	sram_mem[94205] = 16'b0000000000000000;
	sram_mem[94206] = 16'b0000000000000000;
	sram_mem[94207] = 16'b0000000000000000;
	sram_mem[94208] = 16'b0000000000000000;
	sram_mem[94209] = 16'b0000000000000000;
	sram_mem[94210] = 16'b0000000000000000;
	sram_mem[94211] = 16'b0000000000000000;
	sram_mem[94212] = 16'b0000000000000000;
	sram_mem[94213] = 16'b0000000000000000;
	sram_mem[94214] = 16'b0000000000000000;
	sram_mem[94215] = 16'b0000000000000000;
	sram_mem[94216] = 16'b0000000000000000;
	sram_mem[94217] = 16'b0000000000000000;
	sram_mem[94218] = 16'b0000000000000000;
	sram_mem[94219] = 16'b0000000000000000;
	sram_mem[94220] = 16'b0000000000000000;
	sram_mem[94221] = 16'b0000000000000000;
	sram_mem[94222] = 16'b0000000000000000;
	sram_mem[94223] = 16'b0000000000000000;
	sram_mem[94224] = 16'b0000000000000000;
	sram_mem[94225] = 16'b0000000000000000;
	sram_mem[94226] = 16'b0000000000000000;
	sram_mem[94227] = 16'b0000000000000000;
	sram_mem[94228] = 16'b0000000000000000;
	sram_mem[94229] = 16'b0000000000000000;
	sram_mem[94230] = 16'b0000000000000000;
	sram_mem[94231] = 16'b0000000000000000;
	sram_mem[94232] = 16'b0000000000000000;
	sram_mem[94233] = 16'b0000000000000000;
	sram_mem[94234] = 16'b0000000000000000;
	sram_mem[94235] = 16'b0000000000000000;
	sram_mem[94236] = 16'b0000000000000000;
	sram_mem[94237] = 16'b0000000000000000;
	sram_mem[94238] = 16'b0000000000000000;
	sram_mem[94239] = 16'b0000000000000000;
	sram_mem[94240] = 16'b0000000000000000;
	sram_mem[94241] = 16'b0000000000000000;
	sram_mem[94242] = 16'b0000000000000000;
	sram_mem[94243] = 16'b0000000000000000;
	sram_mem[94244] = 16'b0000000000000000;
	sram_mem[94245] = 16'b0000000000000000;
	sram_mem[94246] = 16'b0000000000000000;
	sram_mem[94247] = 16'b0000000000000000;
	sram_mem[94248] = 16'b0000000000000000;
	sram_mem[94249] = 16'b0000000000000000;
	sram_mem[94250] = 16'b0000000000000000;
	sram_mem[94251] = 16'b0000000000000000;
	sram_mem[94252] = 16'b0000000000000000;
	sram_mem[94253] = 16'b0000000000000000;
	sram_mem[94254] = 16'b0000000000000000;
	sram_mem[94255] = 16'b0000000000000000;
	sram_mem[94256] = 16'b0000000000000000;
	sram_mem[94257] = 16'b0000000000000000;
	sram_mem[94258] = 16'b0000000000000000;
	sram_mem[94259] = 16'b0000000000000000;
	sram_mem[94260] = 16'b0000000000000000;
	sram_mem[94261] = 16'b0000000000000000;
	sram_mem[94262] = 16'b0000000000000000;
	sram_mem[94263] = 16'b0000000000000000;
	sram_mem[94264] = 16'b0000000000000000;
	sram_mem[94265] = 16'b0000000000000000;
	sram_mem[94266] = 16'b0000000000000000;
	sram_mem[94267] = 16'b0000000000000000;
	sram_mem[94268] = 16'b0000000000000000;
	sram_mem[94269] = 16'b0000000000000000;
	sram_mem[94270] = 16'b0000000000000000;
	sram_mem[94271] = 16'b0000000000000000;
	sram_mem[94272] = 16'b0000000000000000;
	sram_mem[94273] = 16'b0000000000000000;
	sram_mem[94274] = 16'b0000000000000000;
	sram_mem[94275] = 16'b0000000000000000;
	sram_mem[94276] = 16'b0000000000000000;
	sram_mem[94277] = 16'b0000000000000000;
	sram_mem[94278] = 16'b0000000000000000;
	sram_mem[94279] = 16'b0000000000000000;
	sram_mem[94280] = 16'b0000000000000000;
	sram_mem[94281] = 16'b0000000000000000;
	sram_mem[94282] = 16'b0000000000000000;
	sram_mem[94283] = 16'b0000000000000000;
	sram_mem[94284] = 16'b0000000000000000;
	sram_mem[94285] = 16'b0000000000000000;
	sram_mem[94286] = 16'b0000000000000000;
	sram_mem[94287] = 16'b0000000000000000;
	sram_mem[94288] = 16'b0000000000000000;
	sram_mem[94289] = 16'b0000000000000000;
	sram_mem[94290] = 16'b0000000000000000;
	sram_mem[94291] = 16'b0000000000000000;
	sram_mem[94292] = 16'b0000000000000000;
	sram_mem[94293] = 16'b0000000000000000;
	sram_mem[94294] = 16'b0000000000000000;
	sram_mem[94295] = 16'b0000000000000000;
	sram_mem[94296] = 16'b0000000000000000;
	sram_mem[94297] = 16'b0000000000000000;
	sram_mem[94298] = 16'b0000000000000000;
	sram_mem[94299] = 16'b0000000000000000;
	sram_mem[94300] = 16'b0000000000000000;
	sram_mem[94301] = 16'b0000000000000000;
	sram_mem[94302] = 16'b0000000000000000;
	sram_mem[94303] = 16'b0000000000000000;
	sram_mem[94304] = 16'b0000000000000000;
	sram_mem[94305] = 16'b0000000000000000;
	sram_mem[94306] = 16'b0000000000000000;
	sram_mem[94307] = 16'b0000000000000000;
	sram_mem[94308] = 16'b0000000000000000;
	sram_mem[94309] = 16'b0000000000000000;
	sram_mem[94310] = 16'b0000000000000000;
	sram_mem[94311] = 16'b0000000000000000;
	sram_mem[94312] = 16'b0000000000000000;
	sram_mem[94313] = 16'b0000000000000000;
	sram_mem[94314] = 16'b0000000000000000;
	sram_mem[94315] = 16'b0000000000000000;
	sram_mem[94316] = 16'b0000000000000000;
	sram_mem[94317] = 16'b0000000000000000;
	sram_mem[94318] = 16'b0000000000000000;
	sram_mem[94319] = 16'b0000000000000000;
	sram_mem[94320] = 16'b0000000000000000;
	sram_mem[94321] = 16'b0000000000000000;
	sram_mem[94322] = 16'b0000000000000000;
	sram_mem[94323] = 16'b0000000000000000;
	sram_mem[94324] = 16'b0000000000000000;
	sram_mem[94325] = 16'b0000000000000000;
	sram_mem[94326] = 16'b0000000000000000;
	sram_mem[94327] = 16'b0000000000000000;
	sram_mem[94328] = 16'b0000000000000000;
	sram_mem[94329] = 16'b0000000000000000;
	sram_mem[94330] = 16'b0000000000000000;
	sram_mem[94331] = 16'b0000000000000000;
	sram_mem[94332] = 16'b0000000000000000;
	sram_mem[94333] = 16'b0000000000000000;
	sram_mem[94334] = 16'b0000000000000000;
	sram_mem[94335] = 16'b0000000000000000;
	sram_mem[94336] = 16'b0000000000000000;
	sram_mem[94337] = 16'b0000000000000000;
	sram_mem[94338] = 16'b0000000000000000;
	sram_mem[94339] = 16'b0000000000000000;
	sram_mem[94340] = 16'b0000000000000000;
	sram_mem[94341] = 16'b0000000000000000;
	sram_mem[94342] = 16'b0000000000000000;
	sram_mem[94343] = 16'b0000000000000000;
	sram_mem[94344] = 16'b0000000000000000;
	sram_mem[94345] = 16'b0000000000000000;
	sram_mem[94346] = 16'b0000000000000000;
	sram_mem[94347] = 16'b0000000000000000;
	sram_mem[94348] = 16'b0000000000000000;
	sram_mem[94349] = 16'b0000000000000000;
	sram_mem[94350] = 16'b0000000000000000;
	sram_mem[94351] = 16'b0000000000000000;
	sram_mem[94352] = 16'b0000000000000000;
	sram_mem[94353] = 16'b0000000000000000;
	sram_mem[94354] = 16'b0000000000000000;
	sram_mem[94355] = 16'b0000000000000000;
	sram_mem[94356] = 16'b0000000000000000;
	sram_mem[94357] = 16'b0000000000000000;
	sram_mem[94358] = 16'b0000000000000000;
	sram_mem[94359] = 16'b0000000000000000;
	sram_mem[94360] = 16'b0000000000000000;
	sram_mem[94361] = 16'b0000000000000000;
	sram_mem[94362] = 16'b0000000000000000;
	sram_mem[94363] = 16'b0000000000000000;
	sram_mem[94364] = 16'b0000000000000000;
	sram_mem[94365] = 16'b0000000000000000;
	sram_mem[94366] = 16'b0000000000000000;
	sram_mem[94367] = 16'b0000000000000000;
	sram_mem[94368] = 16'b0000000000000000;
	sram_mem[94369] = 16'b0000000000000000;
	sram_mem[94370] = 16'b0000000000000000;
	sram_mem[94371] = 16'b0000000000000000;
	sram_mem[94372] = 16'b0000000000000000;
	sram_mem[94373] = 16'b0000000000000000;
	sram_mem[94374] = 16'b0000000000000000;
	sram_mem[94375] = 16'b0000000000000000;
	sram_mem[94376] = 16'b0000000000000000;
	sram_mem[94377] = 16'b0000000000000000;
	sram_mem[94378] = 16'b0000000000000000;
	sram_mem[94379] = 16'b0000000000000000;
	sram_mem[94380] = 16'b0000000000000000;
	sram_mem[94381] = 16'b0000000000000000;
	sram_mem[94382] = 16'b0000000000000000;
	sram_mem[94383] = 16'b0000000000000000;
	sram_mem[94384] = 16'b0000000000000000;
	sram_mem[94385] = 16'b0000000000000000;
	sram_mem[94386] = 16'b0000000000000000;
	sram_mem[94387] = 16'b0000000000000000;
	sram_mem[94388] = 16'b0000000000000000;
	sram_mem[94389] = 16'b0000000000000000;
	sram_mem[94390] = 16'b0000000000000000;
	sram_mem[94391] = 16'b0000000000000000;
	sram_mem[94392] = 16'b0000000000000000;
	sram_mem[94393] = 16'b0000000000000000;
	sram_mem[94394] = 16'b0000000000000000;
	sram_mem[94395] = 16'b0000000000000000;
	sram_mem[94396] = 16'b0000000000000000;
	sram_mem[94397] = 16'b0000000000000000;
	sram_mem[94398] = 16'b0000000000000000;
	sram_mem[94399] = 16'b0000000000000000;
	sram_mem[94400] = 16'b0000000000000000;
	sram_mem[94401] = 16'b0000000000000000;
	sram_mem[94402] = 16'b0000000000000000;
	sram_mem[94403] = 16'b0000000000000000;
	sram_mem[94404] = 16'b0000000000000000;
	sram_mem[94405] = 16'b0000000000000000;
	sram_mem[94406] = 16'b0000000000000000;
	sram_mem[94407] = 16'b0000000000000000;
	sram_mem[94408] = 16'b0000000000000000;
	sram_mem[94409] = 16'b0000000000000000;
	sram_mem[94410] = 16'b0000000000000000;
	sram_mem[94411] = 16'b0000000000000000;
	sram_mem[94412] = 16'b0000000000000000;
	sram_mem[94413] = 16'b0000000000000000;
	sram_mem[94414] = 16'b0000000000000000;
	sram_mem[94415] = 16'b0000000000000000;
	sram_mem[94416] = 16'b0000000000000000;
	sram_mem[94417] = 16'b0000000000000000;
	sram_mem[94418] = 16'b0000000000000000;
	sram_mem[94419] = 16'b0000000000000000;
	sram_mem[94420] = 16'b0000000000000000;
	sram_mem[94421] = 16'b0000000000000000;
	sram_mem[94422] = 16'b0000000000000000;
	sram_mem[94423] = 16'b0000000000000000;
	sram_mem[94424] = 16'b0000000000000000;
	sram_mem[94425] = 16'b0000000000000000;
	sram_mem[94426] = 16'b0000000000000000;
	sram_mem[94427] = 16'b0000000000000000;
	sram_mem[94428] = 16'b0000000000000000;
	sram_mem[94429] = 16'b0000000000000000;
	sram_mem[94430] = 16'b0000000000000000;
	sram_mem[94431] = 16'b0000000000000000;
	sram_mem[94432] = 16'b0000000000000000;
	sram_mem[94433] = 16'b0000000000000000;
	sram_mem[94434] = 16'b0000000000000000;
	sram_mem[94435] = 16'b0000000000000000;
	sram_mem[94436] = 16'b0000000000000000;
	sram_mem[94437] = 16'b0000000000000000;
	sram_mem[94438] = 16'b0000000000000000;
	sram_mem[94439] = 16'b0000000000000000;
	sram_mem[94440] = 16'b0000000000000000;
	sram_mem[94441] = 16'b0000000000000000;
	sram_mem[94442] = 16'b0000000000000000;
	sram_mem[94443] = 16'b0000000000000000;
	sram_mem[94444] = 16'b0000000000000000;
	sram_mem[94445] = 16'b0000000000000000;
	sram_mem[94446] = 16'b0000000000000000;
	sram_mem[94447] = 16'b0000000000000000;
	sram_mem[94448] = 16'b0000000000000000;
	sram_mem[94449] = 16'b0000000000000000;
	sram_mem[94450] = 16'b0000000000000000;
	sram_mem[94451] = 16'b0000000000000000;
	sram_mem[94452] = 16'b0000000000000000;
	sram_mem[94453] = 16'b0000000000000000;
	sram_mem[94454] = 16'b0000000000000000;
	sram_mem[94455] = 16'b0000000000000000;
	sram_mem[94456] = 16'b0000000000000000;
	sram_mem[94457] = 16'b0000000000000000;
	sram_mem[94458] = 16'b0000000000000000;
	sram_mem[94459] = 16'b0000000000000000;
	sram_mem[94460] = 16'b0000000000000000;
	sram_mem[94461] = 16'b0000000000000000;
	sram_mem[94462] = 16'b0000000000000000;
	sram_mem[94463] = 16'b0000000000000000;
	sram_mem[94464] = 16'b0000000000000000;
	sram_mem[94465] = 16'b0000000000000000;
	sram_mem[94466] = 16'b0000000000000000;
	sram_mem[94467] = 16'b0000000000000000;
	sram_mem[94468] = 16'b0000000000000000;
	sram_mem[94469] = 16'b0000000000000000;
	sram_mem[94470] = 16'b0000000000000000;
	sram_mem[94471] = 16'b0000000000000000;
	sram_mem[94472] = 16'b0000000000000000;
	sram_mem[94473] = 16'b0000000000000000;
	sram_mem[94474] = 16'b0000000000000000;
	sram_mem[94475] = 16'b0000000000000000;
	sram_mem[94476] = 16'b0000000000000000;
	sram_mem[94477] = 16'b0000000000000000;
	sram_mem[94478] = 16'b0000000000000000;
	sram_mem[94479] = 16'b0000000000000000;
	sram_mem[94480] = 16'b0000000000000000;
	sram_mem[94481] = 16'b0000000000000000;
	sram_mem[94482] = 16'b0000000000000000;
	sram_mem[94483] = 16'b0000000000000000;
	sram_mem[94484] = 16'b0000000000000000;
	sram_mem[94485] = 16'b0000000000000000;
	sram_mem[94486] = 16'b0000000000000000;
	sram_mem[94487] = 16'b0000000000000000;
	sram_mem[94488] = 16'b0000000000000000;
	sram_mem[94489] = 16'b0000000000000000;
	sram_mem[94490] = 16'b0000000000000000;
	sram_mem[94491] = 16'b0000000000000000;
	sram_mem[94492] = 16'b0000000000000000;
	sram_mem[94493] = 16'b0000000000000000;
	sram_mem[94494] = 16'b0000000000000000;
	sram_mem[94495] = 16'b0000000000000000;
	sram_mem[94496] = 16'b0000000000000000;
	sram_mem[94497] = 16'b0000000000000000;
	sram_mem[94498] = 16'b0000000000000000;
	sram_mem[94499] = 16'b0000000000000000;
	sram_mem[94500] = 16'b0000000000000000;
	sram_mem[94501] = 16'b0000000000000000;
	sram_mem[94502] = 16'b0000000000000000;
	sram_mem[94503] = 16'b0000000000000000;
	sram_mem[94504] = 16'b0000000000000000;
	sram_mem[94505] = 16'b0000000000000000;
	sram_mem[94506] = 16'b0000000000000000;
	sram_mem[94507] = 16'b0000000000000000;
	sram_mem[94508] = 16'b0000000000000000;
	sram_mem[94509] = 16'b0000000000000000;
	sram_mem[94510] = 16'b0000000000000000;
	sram_mem[94511] = 16'b0000000000000000;
	sram_mem[94512] = 16'b0000000000000000;
	sram_mem[94513] = 16'b0000000000000000;
	sram_mem[94514] = 16'b0000000000000000;
	sram_mem[94515] = 16'b0000000000000000;
	sram_mem[94516] = 16'b0000000000000000;
	sram_mem[94517] = 16'b0000000000000000;
	sram_mem[94518] = 16'b0000000000000000;
	sram_mem[94519] = 16'b0000000000000000;
	sram_mem[94520] = 16'b0000000000000000;
	sram_mem[94521] = 16'b0000000000000000;
	sram_mem[94522] = 16'b0000000000000000;
	sram_mem[94523] = 16'b0000000000000000;
	sram_mem[94524] = 16'b0000000000000000;
	sram_mem[94525] = 16'b0000000000000000;
	sram_mem[94526] = 16'b0000000000000000;
	sram_mem[94527] = 16'b0000000000000000;
	sram_mem[94528] = 16'b0000000000000000;
	sram_mem[94529] = 16'b0000000000000000;
	sram_mem[94530] = 16'b0000000000000000;
	sram_mem[94531] = 16'b0000000000000000;
	sram_mem[94532] = 16'b0000000000000000;
	sram_mem[94533] = 16'b0000000000000000;
	sram_mem[94534] = 16'b0000000000000000;
	sram_mem[94535] = 16'b0000000000000000;
	sram_mem[94536] = 16'b0000000000000000;
	sram_mem[94537] = 16'b0000000000000000;
	sram_mem[94538] = 16'b0000000000000000;
	sram_mem[94539] = 16'b0000000000000000;
	sram_mem[94540] = 16'b0000000000000000;
	sram_mem[94541] = 16'b0000000000000000;
	sram_mem[94542] = 16'b0000000000000000;
	sram_mem[94543] = 16'b0000000000000000;
	sram_mem[94544] = 16'b0000000000000000;
	sram_mem[94545] = 16'b0000000000000000;
	sram_mem[94546] = 16'b0000000000000000;
	sram_mem[94547] = 16'b0000000000000000;
	sram_mem[94548] = 16'b0000000000000000;
	sram_mem[94549] = 16'b0000000000000000;
	sram_mem[94550] = 16'b0000000000000000;
	sram_mem[94551] = 16'b0000000000000000;
	sram_mem[94552] = 16'b0000000000000000;
	sram_mem[94553] = 16'b0000000000000000;
	sram_mem[94554] = 16'b0000000000000000;
	sram_mem[94555] = 16'b0000000000000000;
	sram_mem[94556] = 16'b0000000000000000;
	sram_mem[94557] = 16'b0000000000000000;
	sram_mem[94558] = 16'b0000000000000000;
	sram_mem[94559] = 16'b0000000000000000;
	sram_mem[94560] = 16'b0000000000000000;
	sram_mem[94561] = 16'b0000000000000000;
	sram_mem[94562] = 16'b0000000000000000;
	sram_mem[94563] = 16'b0000000000000000;
	sram_mem[94564] = 16'b0000000000000000;
	sram_mem[94565] = 16'b0000000000000000;
	sram_mem[94566] = 16'b0000000000000000;
	sram_mem[94567] = 16'b0000000000000000;
	sram_mem[94568] = 16'b0000000000000000;
	sram_mem[94569] = 16'b0000000000000000;
	sram_mem[94570] = 16'b0000000000000000;
	sram_mem[94571] = 16'b0000000000000000;
	sram_mem[94572] = 16'b0000000000000000;
	sram_mem[94573] = 16'b0000000000000000;
	sram_mem[94574] = 16'b0000000000000000;
	sram_mem[94575] = 16'b0000000000000000;
	sram_mem[94576] = 16'b0000000000000000;
	sram_mem[94577] = 16'b0000000000000000;
	sram_mem[94578] = 16'b0000000000000000;
	sram_mem[94579] = 16'b0000000000000000;
	sram_mem[94580] = 16'b0000000000000000;
	sram_mem[94581] = 16'b0000000000000000;
	sram_mem[94582] = 16'b0000000000000000;
	sram_mem[94583] = 16'b0000000000000000;
	sram_mem[94584] = 16'b0000000000000000;
	sram_mem[94585] = 16'b0000000000000000;
	sram_mem[94586] = 16'b0000000000000000;
	sram_mem[94587] = 16'b0000000000000000;
	sram_mem[94588] = 16'b0000000000000000;
	sram_mem[94589] = 16'b0000000000000000;
	sram_mem[94590] = 16'b0000000000000000;
	sram_mem[94591] = 16'b0000000000000000;
	sram_mem[94592] = 16'b0000000000000000;
	sram_mem[94593] = 16'b0000000000000000;
	sram_mem[94594] = 16'b0000000000000000;
	sram_mem[94595] = 16'b0000000000000000;
	sram_mem[94596] = 16'b0000000000000000;
	sram_mem[94597] = 16'b0000000000000000;
	sram_mem[94598] = 16'b0000000000000000;
	sram_mem[94599] = 16'b0000000000000000;
	sram_mem[94600] = 16'b0000000000000000;
	sram_mem[94601] = 16'b0000000000000000;
	sram_mem[94602] = 16'b0000000000000000;
	sram_mem[94603] = 16'b0000000000000000;
	sram_mem[94604] = 16'b0000000000000000;
	sram_mem[94605] = 16'b0000000000000000;
	sram_mem[94606] = 16'b0000000000000000;
	sram_mem[94607] = 16'b0000000000000000;
	sram_mem[94608] = 16'b0000000000000000;
	sram_mem[94609] = 16'b0000000000000000;
	sram_mem[94610] = 16'b0000000000000000;
	sram_mem[94611] = 16'b0000000000000000;
	sram_mem[94612] = 16'b0000000000000000;
	sram_mem[94613] = 16'b0000000000000000;
	sram_mem[94614] = 16'b0000000000000000;
	sram_mem[94615] = 16'b0000000000000000;
	sram_mem[94616] = 16'b0000000000000000;
	sram_mem[94617] = 16'b0000000000000000;
	sram_mem[94618] = 16'b0000000000000000;
	sram_mem[94619] = 16'b0000000000000000;
	sram_mem[94620] = 16'b0000000000000000;
	sram_mem[94621] = 16'b0000000000000000;
	sram_mem[94622] = 16'b0000000000000000;
	sram_mem[94623] = 16'b0000000000000000;
	sram_mem[94624] = 16'b0000000000000000;
	sram_mem[94625] = 16'b0000000000000000;
	sram_mem[94626] = 16'b0000000000000000;
	sram_mem[94627] = 16'b0000000000000000;
	sram_mem[94628] = 16'b0000000000000000;
	sram_mem[94629] = 16'b0000000000000000;
	sram_mem[94630] = 16'b0000000000000000;
	sram_mem[94631] = 16'b0000000000000000;
	sram_mem[94632] = 16'b0000000000000000;
	sram_mem[94633] = 16'b0000000000000000;
	sram_mem[94634] = 16'b0000000000000000;
	sram_mem[94635] = 16'b0000000000000000;
	sram_mem[94636] = 16'b0000000000000000;
	sram_mem[94637] = 16'b0000000000000000;
	sram_mem[94638] = 16'b0000000000000000;
	sram_mem[94639] = 16'b0000000000000000;
	sram_mem[94640] = 16'b0000000000000000;
	sram_mem[94641] = 16'b0000000000000000;
	sram_mem[94642] = 16'b0000000000000000;
	sram_mem[94643] = 16'b0000000000000000;
	sram_mem[94644] = 16'b0000000000000000;
	sram_mem[94645] = 16'b0000000000000000;
	sram_mem[94646] = 16'b0000000000000000;
	sram_mem[94647] = 16'b0000000000000000;
	sram_mem[94648] = 16'b0000000000000000;
	sram_mem[94649] = 16'b0000000000000000;
	sram_mem[94650] = 16'b0000000000000000;
	sram_mem[94651] = 16'b0000000000000000;
	sram_mem[94652] = 16'b0000000000000000;
	sram_mem[94653] = 16'b0000000000000000;
	sram_mem[94654] = 16'b0000000000000000;
	sram_mem[94655] = 16'b0000000000000000;
	sram_mem[94656] = 16'b0000000000000000;
	sram_mem[94657] = 16'b0000000000000000;
	sram_mem[94658] = 16'b0000000000000000;
	sram_mem[94659] = 16'b0000000000000000;
	sram_mem[94660] = 16'b0000000000000000;
	sram_mem[94661] = 16'b0000000000000000;
	sram_mem[94662] = 16'b0000000000000000;
	sram_mem[94663] = 16'b0000000000000000;
	sram_mem[94664] = 16'b0000000000000000;
	sram_mem[94665] = 16'b0000000000000000;
	sram_mem[94666] = 16'b0000000000000000;
	sram_mem[94667] = 16'b0000000000000000;
	sram_mem[94668] = 16'b0000000000000000;
	sram_mem[94669] = 16'b0000000000000000;
	sram_mem[94670] = 16'b0000000000000000;
	sram_mem[94671] = 16'b0000000000000000;
	sram_mem[94672] = 16'b0000000000000000;
	sram_mem[94673] = 16'b0000000000000000;
	sram_mem[94674] = 16'b0000000000000000;
	sram_mem[94675] = 16'b0000000000000000;
	sram_mem[94676] = 16'b0000000000000000;
	sram_mem[94677] = 16'b0000000000000000;
	sram_mem[94678] = 16'b0000000000000000;
	sram_mem[94679] = 16'b0000000000000000;
	sram_mem[94680] = 16'b0000000000000000;
	sram_mem[94681] = 16'b0000000000000000;
	sram_mem[94682] = 16'b0000000000000000;
	sram_mem[94683] = 16'b0000000000000000;
	sram_mem[94684] = 16'b0000000000000000;
	sram_mem[94685] = 16'b0000000000000000;
	sram_mem[94686] = 16'b0000000000000000;
	sram_mem[94687] = 16'b0000000000000000;
	sram_mem[94688] = 16'b0000000000000000;
	sram_mem[94689] = 16'b0000000000000000;
	sram_mem[94690] = 16'b0000000000000000;
	sram_mem[94691] = 16'b0000000000000000;
	sram_mem[94692] = 16'b0000000000000000;
	sram_mem[94693] = 16'b0000000000000000;
	sram_mem[94694] = 16'b0000000000000000;
	sram_mem[94695] = 16'b0000000000000000;
	sram_mem[94696] = 16'b0000000000000000;
	sram_mem[94697] = 16'b0000000000000000;
	sram_mem[94698] = 16'b0000000000000000;
	sram_mem[94699] = 16'b0000000000000000;
	sram_mem[94700] = 16'b0000000000000000;
	sram_mem[94701] = 16'b0000000000000000;
	sram_mem[94702] = 16'b0000000000000000;
	sram_mem[94703] = 16'b0000000000000000;
	sram_mem[94704] = 16'b0000000000000000;
	sram_mem[94705] = 16'b0000000000000000;
	sram_mem[94706] = 16'b0000000000000000;
	sram_mem[94707] = 16'b0000000000000000;
	sram_mem[94708] = 16'b0000000000000000;
	sram_mem[94709] = 16'b0000000000000000;
	sram_mem[94710] = 16'b0000000000000000;
	sram_mem[94711] = 16'b0000000000000000;
	sram_mem[94712] = 16'b0000000000000000;
	sram_mem[94713] = 16'b0000000000000000;
	sram_mem[94714] = 16'b0000000000000000;
	sram_mem[94715] = 16'b0000000000000000;
	sram_mem[94716] = 16'b0000000000000000;
	sram_mem[94717] = 16'b0000000000000000;
	sram_mem[94718] = 16'b0000000000000000;
	sram_mem[94719] = 16'b0000000000000000;
	sram_mem[94720] = 16'b0000000000000000;
	sram_mem[94721] = 16'b0000000000000000;
	sram_mem[94722] = 16'b0000000000000000;
	sram_mem[94723] = 16'b0000000000000000;
	sram_mem[94724] = 16'b0000000000000000;
	sram_mem[94725] = 16'b0000000000000000;
	sram_mem[94726] = 16'b0000000000000000;
	sram_mem[94727] = 16'b0000000000000000;
	sram_mem[94728] = 16'b0000000000000000;
	sram_mem[94729] = 16'b0000000000000000;
	sram_mem[94730] = 16'b0000000000000000;
	sram_mem[94731] = 16'b0000000000000000;
	sram_mem[94732] = 16'b0000000000000000;
	sram_mem[94733] = 16'b0000000000000000;
	sram_mem[94734] = 16'b0000000000000000;
	sram_mem[94735] = 16'b0000000000000000;
	sram_mem[94736] = 16'b0000000000000000;
	sram_mem[94737] = 16'b0000000000000000;
	sram_mem[94738] = 16'b0000000000000000;
	sram_mem[94739] = 16'b0000000000000000;
	sram_mem[94740] = 16'b0000000000000000;
	sram_mem[94741] = 16'b0000000000000000;
	sram_mem[94742] = 16'b0000000000000000;
	sram_mem[94743] = 16'b0000000000000000;
	sram_mem[94744] = 16'b0000000000000000;
	sram_mem[94745] = 16'b0000000000000000;
	sram_mem[94746] = 16'b0000000000000000;
	sram_mem[94747] = 16'b0000000000000000;
	sram_mem[94748] = 16'b0000000000000000;
	sram_mem[94749] = 16'b0000000000000000;
	sram_mem[94750] = 16'b0000000000000000;
	sram_mem[94751] = 16'b0000000000000000;
	sram_mem[94752] = 16'b0000000000000000;
	sram_mem[94753] = 16'b0000000000000000;
	sram_mem[94754] = 16'b0000000000000000;
	sram_mem[94755] = 16'b0000000000000000;
	sram_mem[94756] = 16'b0000000000000000;
	sram_mem[94757] = 16'b0000000000000000;
	sram_mem[94758] = 16'b0000000000000000;
	sram_mem[94759] = 16'b0000000000000000;
	sram_mem[94760] = 16'b0000000000000000;
	sram_mem[94761] = 16'b0000000000000000;
	sram_mem[94762] = 16'b0000000000000000;
	sram_mem[94763] = 16'b0000000000000000;
	sram_mem[94764] = 16'b0000000000000000;
	sram_mem[94765] = 16'b0000000000000000;
	sram_mem[94766] = 16'b0000000000000000;
	sram_mem[94767] = 16'b0000000000000000;
	sram_mem[94768] = 16'b0000000000000000;
	sram_mem[94769] = 16'b0000000000000000;
	sram_mem[94770] = 16'b0000000000000000;
	sram_mem[94771] = 16'b0000000000000000;
	sram_mem[94772] = 16'b0000000000000000;
	sram_mem[94773] = 16'b0000000000000000;
	sram_mem[94774] = 16'b0000000000000000;
	sram_mem[94775] = 16'b0000000000000000;
	sram_mem[94776] = 16'b0000000000000000;
	sram_mem[94777] = 16'b0000000000000000;
	sram_mem[94778] = 16'b0000000000000000;
	sram_mem[94779] = 16'b0000000000000000;
	sram_mem[94780] = 16'b0000000000000000;
	sram_mem[94781] = 16'b0000000000000000;
	sram_mem[94782] = 16'b0000000000000000;
	sram_mem[94783] = 16'b0000000000000000;
	sram_mem[94784] = 16'b0000000000000000;
	sram_mem[94785] = 16'b0000000000000000;
	sram_mem[94786] = 16'b0000000000000000;
	sram_mem[94787] = 16'b0000000000000000;
	sram_mem[94788] = 16'b0000000000000000;
	sram_mem[94789] = 16'b0000000000000000;
	sram_mem[94790] = 16'b0000000000000000;
	sram_mem[94791] = 16'b0000000000000000;
	sram_mem[94792] = 16'b0000000000000000;
	sram_mem[94793] = 16'b0000000000000000;
	sram_mem[94794] = 16'b0000000000000000;
	sram_mem[94795] = 16'b0000000000000000;
	sram_mem[94796] = 16'b0000000000000000;
	sram_mem[94797] = 16'b0000000000000000;
	sram_mem[94798] = 16'b0000000000000000;
	sram_mem[94799] = 16'b0000000000000000;
	sram_mem[94800] = 16'b0000000000000000;
	sram_mem[94801] = 16'b0000000000000000;
	sram_mem[94802] = 16'b0000000000000000;
	sram_mem[94803] = 16'b0000000000000000;
	sram_mem[94804] = 16'b0000000000000000;
	sram_mem[94805] = 16'b0000000000000000;
	sram_mem[94806] = 16'b0000000000000000;
	sram_mem[94807] = 16'b0000000000000000;
	sram_mem[94808] = 16'b0000000000000000;
	sram_mem[94809] = 16'b0000000000000000;
	sram_mem[94810] = 16'b0000000000000000;
	sram_mem[94811] = 16'b0000000000000000;
	sram_mem[94812] = 16'b0000000000000000;
	sram_mem[94813] = 16'b0000000000000000;
	sram_mem[94814] = 16'b0000000000000000;
	sram_mem[94815] = 16'b0000000000000000;
	sram_mem[94816] = 16'b0000000000000000;
	sram_mem[94817] = 16'b0000000000000000;
	sram_mem[94818] = 16'b0000000000000000;
	sram_mem[94819] = 16'b0000000000000000;
	sram_mem[94820] = 16'b0000000000000000;
	sram_mem[94821] = 16'b0000000000000000;
	sram_mem[94822] = 16'b0000000000000000;
	sram_mem[94823] = 16'b0000000000000000;
	sram_mem[94824] = 16'b0000000000000000;
	sram_mem[94825] = 16'b0000000000000000;
	sram_mem[94826] = 16'b0000000000000000;
	sram_mem[94827] = 16'b0000000000000000;
	sram_mem[94828] = 16'b0000000000000000;
	sram_mem[94829] = 16'b0000000000000000;
	sram_mem[94830] = 16'b0000000000000000;
	sram_mem[94831] = 16'b0000000000000000;
	sram_mem[94832] = 16'b0000000000000000;
	sram_mem[94833] = 16'b0000000000000000;
	sram_mem[94834] = 16'b0000000000000000;
	sram_mem[94835] = 16'b0000000000000000;
	sram_mem[94836] = 16'b0000000000000000;
	sram_mem[94837] = 16'b0000000000000000;
	sram_mem[94838] = 16'b0000000000000000;
	sram_mem[94839] = 16'b0000000000000000;
	sram_mem[94840] = 16'b0000000000000000;
	sram_mem[94841] = 16'b0000000000000000;
	sram_mem[94842] = 16'b0000000000000000;
	sram_mem[94843] = 16'b0000000000000000;
	sram_mem[94844] = 16'b0000000000000000;
	sram_mem[94845] = 16'b0000000000000000;
	sram_mem[94846] = 16'b0000000000000000;
	sram_mem[94847] = 16'b0000000000000000;
	sram_mem[94848] = 16'b0000000000000000;
	sram_mem[94849] = 16'b0000000000000000;
	sram_mem[94850] = 16'b0000000000000000;
	sram_mem[94851] = 16'b0000000000000000;
	sram_mem[94852] = 16'b0000000000000000;
	sram_mem[94853] = 16'b0000000000000000;
	sram_mem[94854] = 16'b0000000000000000;
	sram_mem[94855] = 16'b0000000000000000;
	sram_mem[94856] = 16'b0000000000000000;
	sram_mem[94857] = 16'b0000000000000000;
	sram_mem[94858] = 16'b0000000000000000;
	sram_mem[94859] = 16'b0000000000000000;
	sram_mem[94860] = 16'b0000000000000000;
	sram_mem[94861] = 16'b0000000000000000;
	sram_mem[94862] = 16'b0000000000000000;
	sram_mem[94863] = 16'b0000000000000000;
	sram_mem[94864] = 16'b0000000000000000;
	sram_mem[94865] = 16'b0000000000000000;
	sram_mem[94866] = 16'b0000000000000000;
	sram_mem[94867] = 16'b0000000000000000;
	sram_mem[94868] = 16'b0000000000000000;
	sram_mem[94869] = 16'b0000000000000000;
	sram_mem[94870] = 16'b0000000000000000;
	sram_mem[94871] = 16'b0000000000000000;
	sram_mem[94872] = 16'b0000000000000000;
	sram_mem[94873] = 16'b0000000000000000;
	sram_mem[94874] = 16'b0000000000000000;
	sram_mem[94875] = 16'b0000000000000000;
	sram_mem[94876] = 16'b0000000000000000;
	sram_mem[94877] = 16'b0000000000000000;
	sram_mem[94878] = 16'b0000000000000000;
	sram_mem[94879] = 16'b0000000000000000;
	sram_mem[94880] = 16'b0000000000000000;
	sram_mem[94881] = 16'b0000000000000000;
	sram_mem[94882] = 16'b0000000000000000;
	sram_mem[94883] = 16'b0000000000000000;
	sram_mem[94884] = 16'b0000000000000000;
	sram_mem[94885] = 16'b0000000000000000;
	sram_mem[94886] = 16'b0000000000000000;
	sram_mem[94887] = 16'b0000000000000000;
	sram_mem[94888] = 16'b0000000000000000;
	sram_mem[94889] = 16'b0000000000000000;
	sram_mem[94890] = 16'b0000000000000000;
	sram_mem[94891] = 16'b0000000000000000;
	sram_mem[94892] = 16'b0000000000000000;
	sram_mem[94893] = 16'b0000000000000000;
	sram_mem[94894] = 16'b0000000000000000;
	sram_mem[94895] = 16'b0000000000000000;
	sram_mem[94896] = 16'b0000000000000000;
	sram_mem[94897] = 16'b0000000000000000;
	sram_mem[94898] = 16'b0000000000000000;
	sram_mem[94899] = 16'b0000000000000000;
	sram_mem[94900] = 16'b0000000000000000;
	sram_mem[94901] = 16'b0000000000000000;
	sram_mem[94902] = 16'b0000000000000000;
	sram_mem[94903] = 16'b0000000000000000;
	sram_mem[94904] = 16'b0000000000000000;
	sram_mem[94905] = 16'b0000000000000000;
	sram_mem[94906] = 16'b0000000000000000;
	sram_mem[94907] = 16'b0000000000000000;
	sram_mem[94908] = 16'b0000000000000000;
	sram_mem[94909] = 16'b0000000000000000;
	sram_mem[94910] = 16'b0000000000000000;
	sram_mem[94911] = 16'b0000000000000000;
	sram_mem[94912] = 16'b0000000000000000;
	sram_mem[94913] = 16'b0000000000000000;
	sram_mem[94914] = 16'b0000000000000000;
	sram_mem[94915] = 16'b0000000000000000;
	sram_mem[94916] = 16'b0000000000000000;
	sram_mem[94917] = 16'b0000000000000000;
	sram_mem[94918] = 16'b0000000000000000;
	sram_mem[94919] = 16'b0000000000000000;
	sram_mem[94920] = 16'b0000000000000000;
	sram_mem[94921] = 16'b0000000000000000;
	sram_mem[94922] = 16'b0000000000000000;
	sram_mem[94923] = 16'b0000000000000000;
	sram_mem[94924] = 16'b0000000000000000;
	sram_mem[94925] = 16'b0000000000000000;
	sram_mem[94926] = 16'b0000000000000000;
	sram_mem[94927] = 16'b0000000000000000;
	sram_mem[94928] = 16'b0000000000000000;
	sram_mem[94929] = 16'b0000000000000000;
	sram_mem[94930] = 16'b0000000000000000;
	sram_mem[94931] = 16'b0000000000000000;
	sram_mem[94932] = 16'b0000000000000000;
	sram_mem[94933] = 16'b0000000000000000;
	sram_mem[94934] = 16'b0000000000000000;
	sram_mem[94935] = 16'b0000000000000000;
	sram_mem[94936] = 16'b0000000000000000;
	sram_mem[94937] = 16'b0000000000000000;
	sram_mem[94938] = 16'b0000000000000000;
	sram_mem[94939] = 16'b0000000000000000;
	sram_mem[94940] = 16'b0000000000000000;
	sram_mem[94941] = 16'b0000000000000000;
	sram_mem[94942] = 16'b0000000000000000;
	sram_mem[94943] = 16'b0000000000000000;
	sram_mem[94944] = 16'b0000000000000000;
	sram_mem[94945] = 16'b0000000000000000;
	sram_mem[94946] = 16'b0000000000000000;
	sram_mem[94947] = 16'b0000000000000000;
	sram_mem[94948] = 16'b0000000000000000;
	sram_mem[94949] = 16'b0000000000000000;
	sram_mem[94950] = 16'b0000000000000000;
	sram_mem[94951] = 16'b0000000000000000;
	sram_mem[94952] = 16'b0000000000000000;
	sram_mem[94953] = 16'b0000000000000000;
	sram_mem[94954] = 16'b0000000000000000;
	sram_mem[94955] = 16'b0000000000000000;
	sram_mem[94956] = 16'b0000000000000000;
	sram_mem[94957] = 16'b0000000000000000;
	sram_mem[94958] = 16'b0000000000000000;
	sram_mem[94959] = 16'b0000000000000000;
	sram_mem[94960] = 16'b0000000000000000;
	sram_mem[94961] = 16'b0000000000000000;
	sram_mem[94962] = 16'b0000000000000000;
	sram_mem[94963] = 16'b0000000000000000;
	sram_mem[94964] = 16'b0000000000000000;
	sram_mem[94965] = 16'b0000000000000000;
	sram_mem[94966] = 16'b0000000000000000;
	sram_mem[94967] = 16'b0000000000000000;
	sram_mem[94968] = 16'b0000000000000000;
	sram_mem[94969] = 16'b0000000000000000;
	sram_mem[94970] = 16'b0000000000000000;
	sram_mem[94971] = 16'b0000000000000000;
	sram_mem[94972] = 16'b0000000000000000;
	sram_mem[94973] = 16'b0000000000000000;
	sram_mem[94974] = 16'b0000000000000000;
	sram_mem[94975] = 16'b0000000000000000;
	sram_mem[94976] = 16'b0000000000000000;
	sram_mem[94977] = 16'b0000000000000000;
	sram_mem[94978] = 16'b0000000000000000;
	sram_mem[94979] = 16'b0000000000000000;
	sram_mem[94980] = 16'b0000000000000000;
	sram_mem[94981] = 16'b0000000000000000;
	sram_mem[94982] = 16'b0000000000000000;
	sram_mem[94983] = 16'b0000000000000000;
	sram_mem[94984] = 16'b0000000000000000;
	sram_mem[94985] = 16'b0000000000000000;
	sram_mem[94986] = 16'b0000000000000000;
	sram_mem[94987] = 16'b0000000000000000;
	sram_mem[94988] = 16'b0000000000000000;
	sram_mem[94989] = 16'b0000000000000000;
	sram_mem[94990] = 16'b0000000000000000;
	sram_mem[94991] = 16'b0000000000000000;
	sram_mem[94992] = 16'b0000000000000000;
	sram_mem[94993] = 16'b0000000000000000;
	sram_mem[94994] = 16'b0000000000000000;
	sram_mem[94995] = 16'b0000000000000000;
	sram_mem[94996] = 16'b0000000000000000;
	sram_mem[94997] = 16'b0000000000000000;
	sram_mem[94998] = 16'b0000000000000000;
	sram_mem[94999] = 16'b0000000000000000;
	sram_mem[95000] = 16'b0000000000000000;
	sram_mem[95001] = 16'b0000000000000000;
	sram_mem[95002] = 16'b0000000000000000;
	sram_mem[95003] = 16'b0000000000000000;
	sram_mem[95004] = 16'b0000000000000000;
	sram_mem[95005] = 16'b0000000000000000;
	sram_mem[95006] = 16'b0000000000000000;
	sram_mem[95007] = 16'b0000000000000000;
	sram_mem[95008] = 16'b0000000000000000;
	sram_mem[95009] = 16'b0000000000000000;
	sram_mem[95010] = 16'b0000000000000000;
	sram_mem[95011] = 16'b0000000000000000;
	sram_mem[95012] = 16'b0000000000000000;
	sram_mem[95013] = 16'b0000000000000000;
	sram_mem[95014] = 16'b0000000000000000;
	sram_mem[95015] = 16'b0000000000000000;
	sram_mem[95016] = 16'b0000000000000000;
	sram_mem[95017] = 16'b0000000000000000;
	sram_mem[95018] = 16'b0000000000000000;
	sram_mem[95019] = 16'b0000000000000000;
	sram_mem[95020] = 16'b0000000000000000;
	sram_mem[95021] = 16'b0000000000000000;
	sram_mem[95022] = 16'b0000000000000000;
	sram_mem[95023] = 16'b0000000000000000;
	sram_mem[95024] = 16'b0000000000000000;
	sram_mem[95025] = 16'b0000000000000000;
	sram_mem[95026] = 16'b0000000000000000;
	sram_mem[95027] = 16'b0000000000000000;
	sram_mem[95028] = 16'b0000000000000000;
	sram_mem[95029] = 16'b0000000000000000;
	sram_mem[95030] = 16'b0000000000000000;
	sram_mem[95031] = 16'b0000000000000000;
	sram_mem[95032] = 16'b0000000000000000;
	sram_mem[95033] = 16'b0000000000000000;
	sram_mem[95034] = 16'b0000000000000000;
	sram_mem[95035] = 16'b0000000000000000;
	sram_mem[95036] = 16'b0000000000000000;
	sram_mem[95037] = 16'b0000000000000000;
	sram_mem[95038] = 16'b0000000000000000;
	sram_mem[95039] = 16'b0000000000000000;
	sram_mem[95040] = 16'b0000000000000000;
	sram_mem[95041] = 16'b0000000000000000;
	sram_mem[95042] = 16'b0000000000000000;
	sram_mem[95043] = 16'b0000000000000000;
	sram_mem[95044] = 16'b0000000000000000;
	sram_mem[95045] = 16'b0000000000000000;
	sram_mem[95046] = 16'b0000000000000000;
	sram_mem[95047] = 16'b0000000000000000;
	sram_mem[95048] = 16'b0000000000000000;
	sram_mem[95049] = 16'b0000000000000000;
	sram_mem[95050] = 16'b0000000000000000;
	sram_mem[95051] = 16'b0000000000000000;
	sram_mem[95052] = 16'b0000000000000000;
	sram_mem[95053] = 16'b0000000000000000;
	sram_mem[95054] = 16'b0000000000000000;
	sram_mem[95055] = 16'b0000000000000000;
	sram_mem[95056] = 16'b0000000000000000;
	sram_mem[95057] = 16'b0000000000000000;
	sram_mem[95058] = 16'b0000000000000000;
	sram_mem[95059] = 16'b0000000000000000;
	sram_mem[95060] = 16'b0000000000000000;
	sram_mem[95061] = 16'b0000000000000000;
	sram_mem[95062] = 16'b0000000000000000;
	sram_mem[95063] = 16'b0000000000000000;
	sram_mem[95064] = 16'b0000000000000000;
	sram_mem[95065] = 16'b0000000000000000;
	sram_mem[95066] = 16'b0000000000000000;
	sram_mem[95067] = 16'b0000000000000000;
	sram_mem[95068] = 16'b0000000000000000;
	sram_mem[95069] = 16'b0000000000000000;
	sram_mem[95070] = 16'b0000000000000000;
	sram_mem[95071] = 16'b0000000000000000;
	sram_mem[95072] = 16'b0000000000000000;
	sram_mem[95073] = 16'b0000000000000000;
	sram_mem[95074] = 16'b0000000000000000;
	sram_mem[95075] = 16'b0000000000000000;
	sram_mem[95076] = 16'b0000000000000000;
	sram_mem[95077] = 16'b0000000000000000;
	sram_mem[95078] = 16'b0000000000000000;
	sram_mem[95079] = 16'b0000000000000000;
	sram_mem[95080] = 16'b0000000000000000;
	sram_mem[95081] = 16'b0000000000000000;
	sram_mem[95082] = 16'b0000000000000000;
	sram_mem[95083] = 16'b0000000000000000;
	sram_mem[95084] = 16'b0000000000000000;
	sram_mem[95085] = 16'b0000000000000000;
	sram_mem[95086] = 16'b0000000000000000;
	sram_mem[95087] = 16'b0000000000000000;
	sram_mem[95088] = 16'b0000000000000000;
	sram_mem[95089] = 16'b0000000000000000;
	sram_mem[95090] = 16'b0000000000000000;
	sram_mem[95091] = 16'b0000000000000000;
	sram_mem[95092] = 16'b0000000000000000;
	sram_mem[95093] = 16'b0000000000000000;
	sram_mem[95094] = 16'b0000000000000000;
	sram_mem[95095] = 16'b0000000000000000;
	sram_mem[95096] = 16'b0000000000000000;
	sram_mem[95097] = 16'b0000000000000000;
	sram_mem[95098] = 16'b0000000000000000;
	sram_mem[95099] = 16'b0000000000000000;
	sram_mem[95100] = 16'b0000000000000000;
	sram_mem[95101] = 16'b0000000000000000;
	sram_mem[95102] = 16'b0000000000000000;
	sram_mem[95103] = 16'b0000000000000000;
	sram_mem[95104] = 16'b0000000000000000;
	sram_mem[95105] = 16'b0000000000000000;
	sram_mem[95106] = 16'b0000000000000000;
	sram_mem[95107] = 16'b0000000000000000;
	sram_mem[95108] = 16'b0000000000000000;
	sram_mem[95109] = 16'b0000000000000000;
	sram_mem[95110] = 16'b0000000000000000;
	sram_mem[95111] = 16'b0000000000000000;
	sram_mem[95112] = 16'b0000000000000000;
	sram_mem[95113] = 16'b0000000000000000;
	sram_mem[95114] = 16'b0000000000000000;
	sram_mem[95115] = 16'b0000000000000000;
	sram_mem[95116] = 16'b0000000000000000;
	sram_mem[95117] = 16'b0000000000000000;
	sram_mem[95118] = 16'b0000000000000000;
	sram_mem[95119] = 16'b0000000000000000;
	sram_mem[95120] = 16'b0000000000000000;
	sram_mem[95121] = 16'b0000000000000000;
	sram_mem[95122] = 16'b0000000000000000;
	sram_mem[95123] = 16'b0000000000000000;
	sram_mem[95124] = 16'b0000000000000000;
	sram_mem[95125] = 16'b0000000000000000;
	sram_mem[95126] = 16'b0000000000000000;
	sram_mem[95127] = 16'b0000000000000000;
	sram_mem[95128] = 16'b0000000000000000;
	sram_mem[95129] = 16'b0000000000000000;
	sram_mem[95130] = 16'b0000000000000000;
	sram_mem[95131] = 16'b0000000000000000;
	sram_mem[95132] = 16'b0000000000000000;
	sram_mem[95133] = 16'b0000000000000000;
	sram_mem[95134] = 16'b0000000000000000;
	sram_mem[95135] = 16'b0000000000000000;
	sram_mem[95136] = 16'b0000000000000000;
	sram_mem[95137] = 16'b0000000000000000;
	sram_mem[95138] = 16'b0000000000000000;
	sram_mem[95139] = 16'b0000000000000000;
	sram_mem[95140] = 16'b0000000000000000;
	sram_mem[95141] = 16'b0000000000000000;
	sram_mem[95142] = 16'b0000000000000000;
	sram_mem[95143] = 16'b0000000000000000;
	sram_mem[95144] = 16'b0000000000000000;
	sram_mem[95145] = 16'b0000000000000000;
	sram_mem[95146] = 16'b0000000000000000;
	sram_mem[95147] = 16'b0000000000000000;
	sram_mem[95148] = 16'b0000000000000000;
	sram_mem[95149] = 16'b0000000000000000;
	sram_mem[95150] = 16'b0000000000000000;
	sram_mem[95151] = 16'b0000000000000000;
	sram_mem[95152] = 16'b0000000000000000;
	sram_mem[95153] = 16'b0000000000000000;
	sram_mem[95154] = 16'b0000000000000000;
	sram_mem[95155] = 16'b0000000000000000;
	sram_mem[95156] = 16'b0000000000000000;
	sram_mem[95157] = 16'b0000000000000000;
	sram_mem[95158] = 16'b0000000000000000;
	sram_mem[95159] = 16'b0000000000000000;
	sram_mem[95160] = 16'b0000000000000000;
	sram_mem[95161] = 16'b0000000000000000;
	sram_mem[95162] = 16'b0000000000000000;
	sram_mem[95163] = 16'b0000000000000000;
	sram_mem[95164] = 16'b0000000000000000;
	sram_mem[95165] = 16'b0000000000000000;
	sram_mem[95166] = 16'b0000000000000000;
	sram_mem[95167] = 16'b0000000000000000;
	sram_mem[95168] = 16'b0000000000000000;
	sram_mem[95169] = 16'b0000000000000000;
	sram_mem[95170] = 16'b0000000000000000;
	sram_mem[95171] = 16'b0000000000000000;
	sram_mem[95172] = 16'b0000000000000000;
	sram_mem[95173] = 16'b0000000000000000;
	sram_mem[95174] = 16'b0000000000000000;
	sram_mem[95175] = 16'b0000000000000000;
	sram_mem[95176] = 16'b0000000000000000;
	sram_mem[95177] = 16'b0000000000000000;
	sram_mem[95178] = 16'b0000000000000000;
	sram_mem[95179] = 16'b0000000000000000;
	sram_mem[95180] = 16'b0000000000000000;
	sram_mem[95181] = 16'b0000000000000000;
	sram_mem[95182] = 16'b0000000000000000;
	sram_mem[95183] = 16'b0000000000000000;
	sram_mem[95184] = 16'b0000000000000000;
	sram_mem[95185] = 16'b0000000000000000;
	sram_mem[95186] = 16'b0000000000000000;
	sram_mem[95187] = 16'b0000000000000000;
	sram_mem[95188] = 16'b0000000000000000;
	sram_mem[95189] = 16'b0000000000000000;
	sram_mem[95190] = 16'b0000000000000000;
	sram_mem[95191] = 16'b0000000000000000;
	sram_mem[95192] = 16'b0000000000000000;
	sram_mem[95193] = 16'b0000000000000000;
	sram_mem[95194] = 16'b0000000000000000;
	sram_mem[95195] = 16'b0000000000000000;
	sram_mem[95196] = 16'b0000000000000000;
	sram_mem[95197] = 16'b0000000000000000;
	sram_mem[95198] = 16'b0000000000000000;
	sram_mem[95199] = 16'b0000000000000000;
	sram_mem[95200] = 16'b0000000000000000;
	sram_mem[95201] = 16'b0000000000000000;
	sram_mem[95202] = 16'b0000000000000000;
	sram_mem[95203] = 16'b0000000000000000;
	sram_mem[95204] = 16'b0000000000000000;
	sram_mem[95205] = 16'b0000000000000000;
	sram_mem[95206] = 16'b0000000000000000;
	sram_mem[95207] = 16'b0000000000000000;
	sram_mem[95208] = 16'b0000000000000000;
	sram_mem[95209] = 16'b0000000000000000;
	sram_mem[95210] = 16'b0000000000000000;
	sram_mem[95211] = 16'b0000000000000000;
	sram_mem[95212] = 16'b0000000000000000;
	sram_mem[95213] = 16'b0000000000000000;
	sram_mem[95214] = 16'b0000000000000000;
	sram_mem[95215] = 16'b0000000000000000;
	sram_mem[95216] = 16'b0000000000000000;
	sram_mem[95217] = 16'b0000000000000000;
	sram_mem[95218] = 16'b0000000000000000;
	sram_mem[95219] = 16'b0000000000000000;
	sram_mem[95220] = 16'b0000000000000000;
	sram_mem[95221] = 16'b0000000000000000;
	sram_mem[95222] = 16'b0000000000000000;
	sram_mem[95223] = 16'b0000000000000000;
	sram_mem[95224] = 16'b0000000000000000;
	sram_mem[95225] = 16'b0000000000000000;
	sram_mem[95226] = 16'b0000000000000000;
	sram_mem[95227] = 16'b0000000000000000;
	sram_mem[95228] = 16'b0000000000000000;
	sram_mem[95229] = 16'b0000000000000000;
	sram_mem[95230] = 16'b0000000000000000;
	sram_mem[95231] = 16'b0000000000000000;
	sram_mem[95232] = 16'b0000000000000000;
	sram_mem[95233] = 16'b0000000000000000;
	sram_mem[95234] = 16'b0000000000000000;
	sram_mem[95235] = 16'b0000000000000000;
	sram_mem[95236] = 16'b0000000000000000;
	sram_mem[95237] = 16'b0000000000000000;
	sram_mem[95238] = 16'b0000000000000000;
	sram_mem[95239] = 16'b0000000000000000;
	sram_mem[95240] = 16'b0000000000000000;
	sram_mem[95241] = 16'b0000000000000000;
	sram_mem[95242] = 16'b0000000000000000;
	sram_mem[95243] = 16'b0000000000000000;
	sram_mem[95244] = 16'b0000000000000000;
	sram_mem[95245] = 16'b0000000000000000;
	sram_mem[95246] = 16'b0000000000000000;
	sram_mem[95247] = 16'b0000000000000000;
	sram_mem[95248] = 16'b0000000000000000;
	sram_mem[95249] = 16'b0000000000000000;
	sram_mem[95250] = 16'b0000000000000000;
	sram_mem[95251] = 16'b0000000000000000;
	sram_mem[95252] = 16'b0000000000000000;
	sram_mem[95253] = 16'b0000000000000000;
	sram_mem[95254] = 16'b0000000000000000;
	sram_mem[95255] = 16'b0000000000000000;
	sram_mem[95256] = 16'b0000000000000000;
	sram_mem[95257] = 16'b0000000000000000;
	sram_mem[95258] = 16'b0000000000000000;
	sram_mem[95259] = 16'b0000000000000000;
	sram_mem[95260] = 16'b0000000000000000;
	sram_mem[95261] = 16'b0000000000000000;
	sram_mem[95262] = 16'b0000000000000000;
	sram_mem[95263] = 16'b0000000000000000;
	sram_mem[95264] = 16'b0000000000000000;
	sram_mem[95265] = 16'b0000000000000000;
	sram_mem[95266] = 16'b0000000000000000;
	sram_mem[95267] = 16'b0000000000000000;
	sram_mem[95268] = 16'b0000000000000000;
	sram_mem[95269] = 16'b0000000000000000;
	sram_mem[95270] = 16'b0000000000000000;
	sram_mem[95271] = 16'b0000000000000000;
	sram_mem[95272] = 16'b0000000000000000;
	sram_mem[95273] = 16'b0000000000000000;
	sram_mem[95274] = 16'b0000000000000000;
	sram_mem[95275] = 16'b0000000000000000;
	sram_mem[95276] = 16'b0000000000000000;
	sram_mem[95277] = 16'b0000000000000000;
	sram_mem[95278] = 16'b0000000000000000;
	sram_mem[95279] = 16'b0000000000000000;
	sram_mem[95280] = 16'b0000000000000000;
	sram_mem[95281] = 16'b0000000000000000;
	sram_mem[95282] = 16'b0000000000000000;
	sram_mem[95283] = 16'b0000000000000000;
	sram_mem[95284] = 16'b0000000000000000;
	sram_mem[95285] = 16'b0000000000000000;
	sram_mem[95286] = 16'b0000000000000000;
	sram_mem[95287] = 16'b0000000000000000;
	sram_mem[95288] = 16'b0000000000000000;
	sram_mem[95289] = 16'b0000000000000000;
	sram_mem[95290] = 16'b0000000000000000;
	sram_mem[95291] = 16'b0000000000000000;
	sram_mem[95292] = 16'b0000000000000000;
	sram_mem[95293] = 16'b0000000000000000;
	sram_mem[95294] = 16'b0000000000000000;
	sram_mem[95295] = 16'b0000000000000000;
	sram_mem[95296] = 16'b0000000000000000;
	sram_mem[95297] = 16'b0000000000000000;
	sram_mem[95298] = 16'b0000000000000000;
	sram_mem[95299] = 16'b0000000000000000;
	sram_mem[95300] = 16'b0000000000000000;
	sram_mem[95301] = 16'b0000000000000000;
	sram_mem[95302] = 16'b0000000000000000;
	sram_mem[95303] = 16'b0000000000000000;
	sram_mem[95304] = 16'b0000000000000000;
	sram_mem[95305] = 16'b0000000000000000;
	sram_mem[95306] = 16'b0000000000000000;
	sram_mem[95307] = 16'b0000000000000000;
	sram_mem[95308] = 16'b0000000000000000;
	sram_mem[95309] = 16'b0000000000000000;
	sram_mem[95310] = 16'b0000000000000000;
	sram_mem[95311] = 16'b0000000000000000;
	sram_mem[95312] = 16'b0000000000000000;
	sram_mem[95313] = 16'b0000000000000000;
	sram_mem[95314] = 16'b0000000000000000;
	sram_mem[95315] = 16'b0000000000000000;
	sram_mem[95316] = 16'b0000000000000000;
	sram_mem[95317] = 16'b0000000000000000;
	sram_mem[95318] = 16'b0000000000000000;
	sram_mem[95319] = 16'b0000000000000000;
	sram_mem[95320] = 16'b0000000000000000;
	sram_mem[95321] = 16'b0000000000000000;
	sram_mem[95322] = 16'b0000000000000000;
	sram_mem[95323] = 16'b0000000000000000;
	sram_mem[95324] = 16'b0000000000000000;
	sram_mem[95325] = 16'b0000000000000000;
	sram_mem[95326] = 16'b0000000000000000;
	sram_mem[95327] = 16'b0000000000000000;
	sram_mem[95328] = 16'b0000000000000000;
	sram_mem[95329] = 16'b0000000000000000;
	sram_mem[95330] = 16'b0000000000000000;
	sram_mem[95331] = 16'b0000000000000000;
	sram_mem[95332] = 16'b0000000000000000;
	sram_mem[95333] = 16'b0000000000000000;
	sram_mem[95334] = 16'b0000000000000000;
	sram_mem[95335] = 16'b0000000000000000;
	sram_mem[95336] = 16'b0000000000000000;
	sram_mem[95337] = 16'b0000000000000000;
	sram_mem[95338] = 16'b0000000000000000;
	sram_mem[95339] = 16'b0000000000000000;
	sram_mem[95340] = 16'b0000000000000000;
	sram_mem[95341] = 16'b0000000000000000;
	sram_mem[95342] = 16'b0000000000000000;
	sram_mem[95343] = 16'b0000000000000000;
	sram_mem[95344] = 16'b0000000000000000;
	sram_mem[95345] = 16'b0000000000000000;
	sram_mem[95346] = 16'b0000000000000000;
	sram_mem[95347] = 16'b0000000000000000;
	sram_mem[95348] = 16'b0000000000000000;
	sram_mem[95349] = 16'b0000000000000000;
	sram_mem[95350] = 16'b0000000000000000;
	sram_mem[95351] = 16'b0000000000000000;
	sram_mem[95352] = 16'b0000000000000000;
	sram_mem[95353] = 16'b0000000000000000;
	sram_mem[95354] = 16'b0000000000000000;
	sram_mem[95355] = 16'b0000000000000000;
	sram_mem[95356] = 16'b0000000000000000;
	sram_mem[95357] = 16'b0000000000000000;
	sram_mem[95358] = 16'b0000000000000000;
	sram_mem[95359] = 16'b0000000000000000;
	sram_mem[95360] = 16'b0000000000000000;
	sram_mem[95361] = 16'b0000000000000000;
	sram_mem[95362] = 16'b0000000000000000;
	sram_mem[95363] = 16'b0000000000000000;
	sram_mem[95364] = 16'b0000000000000000;
	sram_mem[95365] = 16'b0000000000000000;
	sram_mem[95366] = 16'b0000000000000000;
	sram_mem[95367] = 16'b0000000000000000;
	sram_mem[95368] = 16'b0000000000000000;
	sram_mem[95369] = 16'b0000000000000000;
	sram_mem[95370] = 16'b0000000000000000;
	sram_mem[95371] = 16'b0000000000000000;
	sram_mem[95372] = 16'b0000000000000000;
	sram_mem[95373] = 16'b0000000000000000;
	sram_mem[95374] = 16'b0000000000000000;
	sram_mem[95375] = 16'b0000000000000000;
	sram_mem[95376] = 16'b0000000000000000;
	sram_mem[95377] = 16'b0000000000000000;
	sram_mem[95378] = 16'b0000000000000000;
	sram_mem[95379] = 16'b0000000000000000;
	sram_mem[95380] = 16'b0000000000000000;
	sram_mem[95381] = 16'b0000000000000000;
	sram_mem[95382] = 16'b0000000000000000;
	sram_mem[95383] = 16'b0000000000000000;
	sram_mem[95384] = 16'b0000000000000000;
	sram_mem[95385] = 16'b0000000000000000;
	sram_mem[95386] = 16'b0000000000000000;
	sram_mem[95387] = 16'b0000000000000000;
	sram_mem[95388] = 16'b0000000000000000;
	sram_mem[95389] = 16'b0000000000000000;
	sram_mem[95390] = 16'b0000000000000000;
	sram_mem[95391] = 16'b0000000000000000;
	sram_mem[95392] = 16'b0000000000000000;
	sram_mem[95393] = 16'b0000000000000000;
	sram_mem[95394] = 16'b0000000000000000;
	sram_mem[95395] = 16'b0000000000000000;
	sram_mem[95396] = 16'b0000000000000000;
	sram_mem[95397] = 16'b0000000000000000;
	sram_mem[95398] = 16'b0000000000000000;
	sram_mem[95399] = 16'b0000000000000000;
	sram_mem[95400] = 16'b0000000000000000;
	sram_mem[95401] = 16'b0000000000000000;
	sram_mem[95402] = 16'b0000000000000000;
	sram_mem[95403] = 16'b0000000000000000;
	sram_mem[95404] = 16'b0000000000000000;
	sram_mem[95405] = 16'b0000000000000000;
	sram_mem[95406] = 16'b0000000000000000;
	sram_mem[95407] = 16'b0000000000000000;
	sram_mem[95408] = 16'b0000000000000000;
	sram_mem[95409] = 16'b0000000000000000;
	sram_mem[95410] = 16'b0000000000000000;
	sram_mem[95411] = 16'b0000000000000000;
	sram_mem[95412] = 16'b0000000000000000;
	sram_mem[95413] = 16'b0000000000000000;
	sram_mem[95414] = 16'b0000000000000000;
	sram_mem[95415] = 16'b0000000000000000;
	sram_mem[95416] = 16'b0000000000000000;
	sram_mem[95417] = 16'b0000000000000000;
	sram_mem[95418] = 16'b0000000000000000;
	sram_mem[95419] = 16'b0000000000000000;
	sram_mem[95420] = 16'b0000000000000000;
	sram_mem[95421] = 16'b0000000000000000;
	sram_mem[95422] = 16'b0000000000000000;
	sram_mem[95423] = 16'b0000000000000000;
	sram_mem[95424] = 16'b0000000000000000;
	sram_mem[95425] = 16'b0000000000000000;
	sram_mem[95426] = 16'b0000000000000000;
	sram_mem[95427] = 16'b0000000000000000;
	sram_mem[95428] = 16'b0000000000000000;
	sram_mem[95429] = 16'b0000000000000000;
	sram_mem[95430] = 16'b0000000000000000;
	sram_mem[95431] = 16'b0000000000000000;
	sram_mem[95432] = 16'b0000000000000000;
	sram_mem[95433] = 16'b0000000000000000;
	sram_mem[95434] = 16'b0000000000000000;
	sram_mem[95435] = 16'b0000000000000000;
	sram_mem[95436] = 16'b0000000000000000;
	sram_mem[95437] = 16'b0000000000000000;
	sram_mem[95438] = 16'b0000000000000000;
	sram_mem[95439] = 16'b0000000000000000;
	sram_mem[95440] = 16'b0000000000000000;
	sram_mem[95441] = 16'b0000000000000000;
	sram_mem[95442] = 16'b0000000000000000;
	sram_mem[95443] = 16'b0000000000000000;
	sram_mem[95444] = 16'b0000000000000000;
	sram_mem[95445] = 16'b0000000000000000;
	sram_mem[95446] = 16'b0000000000000000;
	sram_mem[95447] = 16'b0000000000000000;
	sram_mem[95448] = 16'b0000000000000000;
	sram_mem[95449] = 16'b0000000000000000;
	sram_mem[95450] = 16'b0000000000000000;
	sram_mem[95451] = 16'b0000000000000000;
	sram_mem[95452] = 16'b0000000000000000;
	sram_mem[95453] = 16'b0000000000000000;
	sram_mem[95454] = 16'b0000000000000000;
	sram_mem[95455] = 16'b0000000000000000;
	sram_mem[95456] = 16'b0000000000000000;
	sram_mem[95457] = 16'b0000000000000000;
	sram_mem[95458] = 16'b0000000000000000;
	sram_mem[95459] = 16'b0000000000000000;
	sram_mem[95460] = 16'b0000000000000000;
	sram_mem[95461] = 16'b0000000000000000;
	sram_mem[95462] = 16'b0000000000000000;
	sram_mem[95463] = 16'b0000000000000000;
	sram_mem[95464] = 16'b0000000000000000;
	sram_mem[95465] = 16'b0000000000000000;
	sram_mem[95466] = 16'b0000000000000000;
	sram_mem[95467] = 16'b0000000000000000;
	sram_mem[95468] = 16'b0000000000000000;
	sram_mem[95469] = 16'b0000000000000000;
	sram_mem[95470] = 16'b0000000000000000;
	sram_mem[95471] = 16'b0000000000000000;
	sram_mem[95472] = 16'b0000000000000000;
	sram_mem[95473] = 16'b0000000000000000;
	sram_mem[95474] = 16'b0000000000000000;
	sram_mem[95475] = 16'b0000000000000000;
	sram_mem[95476] = 16'b0000000000000000;
	sram_mem[95477] = 16'b0000000000000000;
	sram_mem[95478] = 16'b0000000000000000;
	sram_mem[95479] = 16'b0000000000000000;
	sram_mem[95480] = 16'b0000000000000000;
	sram_mem[95481] = 16'b0000000000000000;
	sram_mem[95482] = 16'b0000000000000000;
	sram_mem[95483] = 16'b0000000000000000;
	sram_mem[95484] = 16'b0000000000000000;
	sram_mem[95485] = 16'b0000000000000000;
	sram_mem[95486] = 16'b0000000000000000;
	sram_mem[95487] = 16'b0000000000000000;
	sram_mem[95488] = 16'b0000000000000000;
	sram_mem[95489] = 16'b0000000000000000;
	sram_mem[95490] = 16'b0000000000000000;
	sram_mem[95491] = 16'b0000000000000000;
	sram_mem[95492] = 16'b0000000000000000;
	sram_mem[95493] = 16'b0000000000000000;
	sram_mem[95494] = 16'b0000000000000000;
	sram_mem[95495] = 16'b0000000000000000;
	sram_mem[95496] = 16'b0000000000000000;
	sram_mem[95497] = 16'b0000000000000000;
	sram_mem[95498] = 16'b0000000000000000;
	sram_mem[95499] = 16'b0000000000000000;
	sram_mem[95500] = 16'b0000000000000000;
	sram_mem[95501] = 16'b0000000000000000;
	sram_mem[95502] = 16'b0000000000000000;
	sram_mem[95503] = 16'b0000000000000000;
	sram_mem[95504] = 16'b0000000000000000;
	sram_mem[95505] = 16'b0000000000000000;
	sram_mem[95506] = 16'b0000000000000000;
	sram_mem[95507] = 16'b0000000000000000;
	sram_mem[95508] = 16'b0000000000000000;
	sram_mem[95509] = 16'b0000000000000000;
	sram_mem[95510] = 16'b0000000000000000;
	sram_mem[95511] = 16'b0000000000000000;
	sram_mem[95512] = 16'b0000000000000000;
	sram_mem[95513] = 16'b0000000000000000;
	sram_mem[95514] = 16'b0000000000000000;
	sram_mem[95515] = 16'b0000000000000000;
	sram_mem[95516] = 16'b0000000000000000;
	sram_mem[95517] = 16'b0000000000000000;
	sram_mem[95518] = 16'b0000000000000000;
	sram_mem[95519] = 16'b0000000000000000;
	sram_mem[95520] = 16'b0000000000000000;
	sram_mem[95521] = 16'b0000000000000000;
	sram_mem[95522] = 16'b0000000000000000;
	sram_mem[95523] = 16'b0000000000000000;
	sram_mem[95524] = 16'b0000000000000000;
	sram_mem[95525] = 16'b0000000000000000;
	sram_mem[95526] = 16'b0000000000000000;
	sram_mem[95527] = 16'b0000000000000000;
	sram_mem[95528] = 16'b0000000000000000;
	sram_mem[95529] = 16'b0000000000000000;
	sram_mem[95530] = 16'b0000000000000000;
	sram_mem[95531] = 16'b0000000000000000;
	sram_mem[95532] = 16'b0000000000000000;
	sram_mem[95533] = 16'b0000000000000000;
	sram_mem[95534] = 16'b0000000000000000;
	sram_mem[95535] = 16'b0000000000000000;
	sram_mem[95536] = 16'b0000000000000000;
	sram_mem[95537] = 16'b0000000000000000;
	sram_mem[95538] = 16'b0000000000000000;
	sram_mem[95539] = 16'b0000000000000000;
	sram_mem[95540] = 16'b0000000000000000;
	sram_mem[95541] = 16'b0000000000000000;
	sram_mem[95542] = 16'b0000000000000000;
	sram_mem[95543] = 16'b0000000000000000;
	sram_mem[95544] = 16'b0000000000000000;
	sram_mem[95545] = 16'b0000000000000000;
	sram_mem[95546] = 16'b0000000000000000;
	sram_mem[95547] = 16'b0000000000000000;
	sram_mem[95548] = 16'b0000000000000000;
	sram_mem[95549] = 16'b0000000000000000;
	sram_mem[95550] = 16'b0000000000000000;
	sram_mem[95551] = 16'b0000000000000000;
	sram_mem[95552] = 16'b0000000000000000;
	sram_mem[95553] = 16'b0000000000000000;
	sram_mem[95554] = 16'b0000000000000000;
	sram_mem[95555] = 16'b0000000000000000;
	sram_mem[95556] = 16'b0000000000000000;
	sram_mem[95557] = 16'b0000000000000000;
	sram_mem[95558] = 16'b0000000000000000;
	sram_mem[95559] = 16'b0000000000000000;
	sram_mem[95560] = 16'b0000000000000000;
	sram_mem[95561] = 16'b0000000000000000;
	sram_mem[95562] = 16'b0000000000000000;
	sram_mem[95563] = 16'b0000000000000000;
	sram_mem[95564] = 16'b0000000000000000;
	sram_mem[95565] = 16'b0000000000000000;
	sram_mem[95566] = 16'b0000000000000000;
	sram_mem[95567] = 16'b0000000000000000;
	sram_mem[95568] = 16'b0000000000000000;
	sram_mem[95569] = 16'b0000000000000000;
	sram_mem[95570] = 16'b0000000000000000;
	sram_mem[95571] = 16'b0000000000000000;
	sram_mem[95572] = 16'b0000000000000000;
	sram_mem[95573] = 16'b0000000000000000;
	sram_mem[95574] = 16'b0000000000000000;
	sram_mem[95575] = 16'b0000000000000000;
	sram_mem[95576] = 16'b0000000000000000;
	sram_mem[95577] = 16'b0000000000000000;
	sram_mem[95578] = 16'b0000000000000000;
	sram_mem[95579] = 16'b0000000000000000;
	sram_mem[95580] = 16'b0000000000000000;
	sram_mem[95581] = 16'b0000000000000000;
	sram_mem[95582] = 16'b0000000000000000;
	sram_mem[95583] = 16'b0000000000000000;
	sram_mem[95584] = 16'b0000000000000000;
	sram_mem[95585] = 16'b0000000000000000;
	sram_mem[95586] = 16'b0000000000000000;
	sram_mem[95587] = 16'b0000000000000000;
	sram_mem[95588] = 16'b0000000000000000;
	sram_mem[95589] = 16'b0000000000000000;
	sram_mem[95590] = 16'b0000000000000000;
	sram_mem[95591] = 16'b0000000000000000;
	sram_mem[95592] = 16'b0000000000000000;
	sram_mem[95593] = 16'b0000000000000000;
	sram_mem[95594] = 16'b0000000000000000;
	sram_mem[95595] = 16'b0000000000000000;
	sram_mem[95596] = 16'b0000000000000000;
	sram_mem[95597] = 16'b0000000000000000;
	sram_mem[95598] = 16'b0000000000000000;
	sram_mem[95599] = 16'b0000000000000000;
	sram_mem[95600] = 16'b0000000000000000;
	sram_mem[95601] = 16'b0000000000000000;
	sram_mem[95602] = 16'b0000000000000000;
	sram_mem[95603] = 16'b0000000000000000;
	sram_mem[95604] = 16'b0000000000000000;
	sram_mem[95605] = 16'b0000000000000000;
	sram_mem[95606] = 16'b0000000000000000;
	sram_mem[95607] = 16'b0000000000000000;
	sram_mem[95608] = 16'b0000000000000000;
	sram_mem[95609] = 16'b0000000000000000;
	sram_mem[95610] = 16'b0000000000000000;
	sram_mem[95611] = 16'b0000000000000000;
	sram_mem[95612] = 16'b0000000000000000;
	sram_mem[95613] = 16'b0000000000000000;
	sram_mem[95614] = 16'b0000000000000000;
	sram_mem[95615] = 16'b0000000000000000;
	sram_mem[95616] = 16'b0000000000000000;
	sram_mem[95617] = 16'b0000000000000000;
	sram_mem[95618] = 16'b0000000000000000;
	sram_mem[95619] = 16'b0000000000000000;
	sram_mem[95620] = 16'b0000000000000000;
	sram_mem[95621] = 16'b0000000000000000;
	sram_mem[95622] = 16'b0000000000000000;
	sram_mem[95623] = 16'b0000000000000000;
	sram_mem[95624] = 16'b0000000000000000;
	sram_mem[95625] = 16'b0000000000000000;
	sram_mem[95626] = 16'b0000000000000000;
	sram_mem[95627] = 16'b0000000000000000;
	sram_mem[95628] = 16'b0000000000000000;
	sram_mem[95629] = 16'b0000000000000000;
	sram_mem[95630] = 16'b0000000000000000;
	sram_mem[95631] = 16'b0000000000000000;
	sram_mem[95632] = 16'b0000000000000000;
	sram_mem[95633] = 16'b0000000000000000;
	sram_mem[95634] = 16'b0000000000000000;
	sram_mem[95635] = 16'b0000000000000000;
	sram_mem[95636] = 16'b0000000000000000;
	sram_mem[95637] = 16'b0000000000000000;
	sram_mem[95638] = 16'b0000000000000000;
	sram_mem[95639] = 16'b0000000000000000;
	sram_mem[95640] = 16'b0000000000000000;
	sram_mem[95641] = 16'b0000000000000000;
	sram_mem[95642] = 16'b0000000000000000;
	sram_mem[95643] = 16'b0000000000000000;
	sram_mem[95644] = 16'b0000000000000000;
	sram_mem[95645] = 16'b0000000000000000;
	sram_mem[95646] = 16'b0000000000000000;
	sram_mem[95647] = 16'b0000000000000000;
	sram_mem[95648] = 16'b0000000000000000;
	sram_mem[95649] = 16'b0000000000000000;
	sram_mem[95650] = 16'b0000000000000000;
	sram_mem[95651] = 16'b0000000000000000;
	sram_mem[95652] = 16'b0000000000000000;
	sram_mem[95653] = 16'b0000000000000000;
	sram_mem[95654] = 16'b0000000000000000;
	sram_mem[95655] = 16'b0000000000000000;
	sram_mem[95656] = 16'b0000000000000000;
	sram_mem[95657] = 16'b0000000000000000;
	sram_mem[95658] = 16'b0000000000000000;
	sram_mem[95659] = 16'b0000000000000000;
	sram_mem[95660] = 16'b0000000000000000;
	sram_mem[95661] = 16'b0000000000000000;
	sram_mem[95662] = 16'b0000000000000000;
	sram_mem[95663] = 16'b0000000000000000;
	sram_mem[95664] = 16'b0000000000000000;
	sram_mem[95665] = 16'b0000000000000000;
	sram_mem[95666] = 16'b0000000000000000;
	sram_mem[95667] = 16'b0000000000000000;
	sram_mem[95668] = 16'b0000000000000000;
	sram_mem[95669] = 16'b0000000000000000;
	sram_mem[95670] = 16'b0000000000000000;
	sram_mem[95671] = 16'b0000000000000000;
	sram_mem[95672] = 16'b0000000000000000;
	sram_mem[95673] = 16'b0000000000000000;
	sram_mem[95674] = 16'b0000000000000000;
	sram_mem[95675] = 16'b0000000000000000;
	sram_mem[95676] = 16'b0000000000000000;
	sram_mem[95677] = 16'b0000000000000000;
	sram_mem[95678] = 16'b0000000000000000;
	sram_mem[95679] = 16'b0000000000000000;
	sram_mem[95680] = 16'b0000000000000000;
	sram_mem[95681] = 16'b0000000000000000;
	sram_mem[95682] = 16'b0000000000000000;
	sram_mem[95683] = 16'b0000000000000000;
	sram_mem[95684] = 16'b0000000000000000;
	sram_mem[95685] = 16'b0000000000000000;
	sram_mem[95686] = 16'b0000000000000000;
	sram_mem[95687] = 16'b0000000000000000;
	sram_mem[95688] = 16'b0000000000000000;
	sram_mem[95689] = 16'b0000000000000000;
	sram_mem[95690] = 16'b0000000000000000;
	sram_mem[95691] = 16'b0000000000000000;
	sram_mem[95692] = 16'b0000000000000000;
	sram_mem[95693] = 16'b0000000000000000;
	sram_mem[95694] = 16'b0000000000000000;
	sram_mem[95695] = 16'b0000000000000000;
	sram_mem[95696] = 16'b0000000000000000;
	sram_mem[95697] = 16'b0000000000000000;
	sram_mem[95698] = 16'b0000000000000000;
	sram_mem[95699] = 16'b0000000000000000;
	sram_mem[95700] = 16'b0000000000000000;
	sram_mem[95701] = 16'b0000000000000000;
	sram_mem[95702] = 16'b0000000000000000;
	sram_mem[95703] = 16'b0000000000000000;
	sram_mem[95704] = 16'b0000000000000000;
	sram_mem[95705] = 16'b0000000000000000;
	sram_mem[95706] = 16'b0000000000000000;
	sram_mem[95707] = 16'b0000000000000000;
	sram_mem[95708] = 16'b0000000000000000;
	sram_mem[95709] = 16'b0000000000000000;
	sram_mem[95710] = 16'b0000000000000000;
	sram_mem[95711] = 16'b0000000000000000;
	sram_mem[95712] = 16'b0000000000000000;
	sram_mem[95713] = 16'b0000000000000000;
	sram_mem[95714] = 16'b0000000000000000;
	sram_mem[95715] = 16'b0000000000000000;
	sram_mem[95716] = 16'b0000000000000000;
	sram_mem[95717] = 16'b0000000000000000;
	sram_mem[95718] = 16'b0000000000000000;
	sram_mem[95719] = 16'b0000000000000000;
	sram_mem[95720] = 16'b0000000000000000;
	sram_mem[95721] = 16'b0000000000000000;
	sram_mem[95722] = 16'b0000000000000000;
	sram_mem[95723] = 16'b0000000000000000;
	sram_mem[95724] = 16'b0000000000000000;
	sram_mem[95725] = 16'b0000000000000000;
	sram_mem[95726] = 16'b0000000000000000;
	sram_mem[95727] = 16'b0000000000000000;
	sram_mem[95728] = 16'b0000000000000000;
	sram_mem[95729] = 16'b0000000000000000;
	sram_mem[95730] = 16'b0000000000000000;
	sram_mem[95731] = 16'b0000000000000000;
	sram_mem[95732] = 16'b0000000000000000;
	sram_mem[95733] = 16'b0000000000000000;
	sram_mem[95734] = 16'b0000000000000000;
	sram_mem[95735] = 16'b0000000000000000;
	sram_mem[95736] = 16'b0000000000000000;
	sram_mem[95737] = 16'b0000000000000000;
	sram_mem[95738] = 16'b0000000000000000;
	sram_mem[95739] = 16'b0000000000000000;
	sram_mem[95740] = 16'b0000000000000000;
	sram_mem[95741] = 16'b0000000000000000;
	sram_mem[95742] = 16'b0000000000000000;
	sram_mem[95743] = 16'b0000000000000000;
	sram_mem[95744] = 16'b0000000000000000;
	sram_mem[95745] = 16'b0000000000000000;
	sram_mem[95746] = 16'b0000000000000000;
	sram_mem[95747] = 16'b0000000000000000;
	sram_mem[95748] = 16'b0000000000000000;
	sram_mem[95749] = 16'b0000000000000000;
	sram_mem[95750] = 16'b0000000000000000;
	sram_mem[95751] = 16'b0000000000000000;
	sram_mem[95752] = 16'b0000000000000000;
	sram_mem[95753] = 16'b0000000000000000;
	sram_mem[95754] = 16'b0000000000000000;
	sram_mem[95755] = 16'b0000000000000000;
	sram_mem[95756] = 16'b0000000000000000;
	sram_mem[95757] = 16'b0000000000000000;
	sram_mem[95758] = 16'b0000000000000000;
	sram_mem[95759] = 16'b0000000000000000;
	sram_mem[95760] = 16'b0000000000000000;
	sram_mem[95761] = 16'b0000000000000000;
	sram_mem[95762] = 16'b0000000000000000;
	sram_mem[95763] = 16'b0000000000000000;
	sram_mem[95764] = 16'b0000000000000000;
	sram_mem[95765] = 16'b0000000000000000;
	sram_mem[95766] = 16'b0000000000000000;
	sram_mem[95767] = 16'b0000000000000000;
	sram_mem[95768] = 16'b0000000000000000;
	sram_mem[95769] = 16'b0000000000000000;
	sram_mem[95770] = 16'b0000000000000000;
	sram_mem[95771] = 16'b0000000000000000;
	sram_mem[95772] = 16'b0000000000000000;
	sram_mem[95773] = 16'b0000000000000000;
	sram_mem[95774] = 16'b0000000000000000;
	sram_mem[95775] = 16'b0000000000000000;
	sram_mem[95776] = 16'b0000000000000000;
	sram_mem[95777] = 16'b0000000000000000;
	sram_mem[95778] = 16'b0000000000000000;
	sram_mem[95779] = 16'b0000000000000000;
	sram_mem[95780] = 16'b0000000000000000;
	sram_mem[95781] = 16'b0000000000000000;
	sram_mem[95782] = 16'b0000000000000000;
	sram_mem[95783] = 16'b0000000000000000;
	sram_mem[95784] = 16'b0000000000000000;
	sram_mem[95785] = 16'b0000000000000000;
	sram_mem[95786] = 16'b0000000000000000;
	sram_mem[95787] = 16'b0000000000000000;
	sram_mem[95788] = 16'b0000000000000000;
	sram_mem[95789] = 16'b0000000000000000;
	sram_mem[95790] = 16'b0000000000000000;
	sram_mem[95791] = 16'b0000000000000000;
	sram_mem[95792] = 16'b0000000000000000;
	sram_mem[95793] = 16'b0000000000000000;
	sram_mem[95794] = 16'b0000000000000000;
	sram_mem[95795] = 16'b0000000000000000;
	sram_mem[95796] = 16'b0000000000000000;
	sram_mem[95797] = 16'b0000000000000000;
	sram_mem[95798] = 16'b0000000000000000;
	sram_mem[95799] = 16'b0000000000000000;
	sram_mem[95800] = 16'b0000000000000000;
	sram_mem[95801] = 16'b0000000000000000;
	sram_mem[95802] = 16'b0000000000000000;
	sram_mem[95803] = 16'b0000000000000000;
	sram_mem[95804] = 16'b0000000000000000;
	sram_mem[95805] = 16'b0000000000000000;
	sram_mem[95806] = 16'b0000000000000000;
	sram_mem[95807] = 16'b0000000000000000;
	sram_mem[95808] = 16'b0000000000000000;
	sram_mem[95809] = 16'b0000000000000000;
	sram_mem[95810] = 16'b0000000000000000;
	sram_mem[95811] = 16'b0000000000000000;
	sram_mem[95812] = 16'b0000000000000000;
	sram_mem[95813] = 16'b0000000000000000;
	sram_mem[95814] = 16'b0000000000000000;
	sram_mem[95815] = 16'b0000000000000000;
	sram_mem[95816] = 16'b0000000000000000;
	sram_mem[95817] = 16'b0000000000000000;
	sram_mem[95818] = 16'b0000000000000000;
	sram_mem[95819] = 16'b0000000000000000;
	sram_mem[95820] = 16'b0000000000000000;
	sram_mem[95821] = 16'b0000000000000000;
	sram_mem[95822] = 16'b0000000000000000;
	sram_mem[95823] = 16'b0000000000000000;
	sram_mem[95824] = 16'b0000000000000000;
	sram_mem[95825] = 16'b0000000000000000;
	sram_mem[95826] = 16'b0000000000000000;
	sram_mem[95827] = 16'b0000000000000000;
	sram_mem[95828] = 16'b0000000000000000;
	sram_mem[95829] = 16'b0000000000000000;
	sram_mem[95830] = 16'b0000000000000000;
	sram_mem[95831] = 16'b0000000000000000;
	sram_mem[95832] = 16'b0000000000000000;
	sram_mem[95833] = 16'b0000000000000000;
	sram_mem[95834] = 16'b0000000000000000;
	sram_mem[95835] = 16'b0000000000000000;
	sram_mem[95836] = 16'b0000000000000000;
	sram_mem[95837] = 16'b0000000000000000;
	sram_mem[95838] = 16'b0000000000000000;
	sram_mem[95839] = 16'b0000000000000000;
	sram_mem[95840] = 16'b0000000000000000;
	sram_mem[95841] = 16'b0000000000000000;
	sram_mem[95842] = 16'b0000000000000000;
	sram_mem[95843] = 16'b0000000000000000;
	sram_mem[95844] = 16'b0000000000000000;
	sram_mem[95845] = 16'b0000000000000000;
	sram_mem[95846] = 16'b0000000000000000;
	sram_mem[95847] = 16'b0000000000000000;
	sram_mem[95848] = 16'b0000000000000000;
	sram_mem[95849] = 16'b0000000000000000;
	sram_mem[95850] = 16'b0000000000000000;
	sram_mem[95851] = 16'b0000000000000000;
	sram_mem[95852] = 16'b0000000000000000;
	sram_mem[95853] = 16'b0000000000000000;
	sram_mem[95854] = 16'b0000000000000000;
	sram_mem[95855] = 16'b0000000000000000;
	sram_mem[95856] = 16'b0000000000000000;
	sram_mem[95857] = 16'b0000000000000000;
	sram_mem[95858] = 16'b0000000000000000;
	sram_mem[95859] = 16'b0000000000000000;
	sram_mem[95860] = 16'b0000000000000000;
	sram_mem[95861] = 16'b0000000000000000;
	sram_mem[95862] = 16'b0000000000000000;
	sram_mem[95863] = 16'b0000000000000000;
	sram_mem[95864] = 16'b0000000000000000;
	sram_mem[95865] = 16'b0000000000000000;
	sram_mem[95866] = 16'b0000000000000000;
	sram_mem[95867] = 16'b0000000000000000;
	sram_mem[95868] = 16'b0000000000000000;
	sram_mem[95869] = 16'b0000000000000000;
	sram_mem[95870] = 16'b0000000000000000;
	sram_mem[95871] = 16'b0000000000000000;
	sram_mem[95872] = 16'b0000000000000000;
	sram_mem[95873] = 16'b0000000000000000;
	sram_mem[95874] = 16'b0000000000000000;
	sram_mem[95875] = 16'b0000000000000000;
	sram_mem[95876] = 16'b0000000000000000;
	sram_mem[95877] = 16'b0000000000000000;
	sram_mem[95878] = 16'b0000000000000000;
	sram_mem[95879] = 16'b0000000000000000;
	sram_mem[95880] = 16'b0000000000000000;
	sram_mem[95881] = 16'b0000000000000000;
	sram_mem[95882] = 16'b0000000000000000;
	sram_mem[95883] = 16'b0000000000000000;
	sram_mem[95884] = 16'b0000000000000000;
	sram_mem[95885] = 16'b0000000000000000;
	sram_mem[95886] = 16'b0000000000000000;
	sram_mem[95887] = 16'b0000000000000000;
	sram_mem[95888] = 16'b0000000000000000;
	sram_mem[95889] = 16'b0000000000000000;
	sram_mem[95890] = 16'b0000000000000000;
	sram_mem[95891] = 16'b0000000000000000;
	sram_mem[95892] = 16'b0000000000000000;
	sram_mem[95893] = 16'b0000000000000000;
	sram_mem[95894] = 16'b0000000000000000;
	sram_mem[95895] = 16'b0000000000000000;
	sram_mem[95896] = 16'b0000000000000000;
	sram_mem[95897] = 16'b0000000000000000;
	sram_mem[95898] = 16'b0000000000000000;
	sram_mem[95899] = 16'b0000000000000000;
	sram_mem[95900] = 16'b0000000000000000;
	sram_mem[95901] = 16'b0000000000000000;
	sram_mem[95902] = 16'b0000000000000000;
	sram_mem[95903] = 16'b0000000000000000;
	sram_mem[95904] = 16'b0000000000000000;
	sram_mem[95905] = 16'b0000000000000000;
	sram_mem[95906] = 16'b0000000000000000;
	sram_mem[95907] = 16'b0000000000000000;
	sram_mem[95908] = 16'b0000000000000000;
	sram_mem[95909] = 16'b0000000000000000;
	sram_mem[95910] = 16'b0000000000000000;
	sram_mem[95911] = 16'b0000000000000000;
	sram_mem[95912] = 16'b0000000000000000;
	sram_mem[95913] = 16'b0000000000000000;
	sram_mem[95914] = 16'b0000000000000000;
	sram_mem[95915] = 16'b0000000000000000;
	sram_mem[95916] = 16'b0000000000000000;
	sram_mem[95917] = 16'b0000000000000000;
	sram_mem[95918] = 16'b0000000000000000;
	sram_mem[95919] = 16'b0000000000000000;
	sram_mem[95920] = 16'b0000000000000000;
	sram_mem[95921] = 16'b0000000000000000;
	sram_mem[95922] = 16'b0000000000000000;
	sram_mem[95923] = 16'b0000000000000000;
	sram_mem[95924] = 16'b0000000000000000;
	sram_mem[95925] = 16'b0000000000000000;
	sram_mem[95926] = 16'b0000000000000000;
	sram_mem[95927] = 16'b0000000000000000;
	sram_mem[95928] = 16'b0000000000000000;
	sram_mem[95929] = 16'b0000000000000000;
	sram_mem[95930] = 16'b0000000000000000;
	sram_mem[95931] = 16'b0000000000000000;
	sram_mem[95932] = 16'b0000000000000000;
	sram_mem[95933] = 16'b0000000000000000;
	sram_mem[95934] = 16'b0000000000000000;
	sram_mem[95935] = 16'b0000000000000000;
	sram_mem[95936] = 16'b0000000000000000;
	sram_mem[95937] = 16'b0000000000000000;
	sram_mem[95938] = 16'b0000000000000000;
	sram_mem[95939] = 16'b0000000000000000;
	sram_mem[95940] = 16'b0000000000000000;
	sram_mem[95941] = 16'b0000000000000000;
	sram_mem[95942] = 16'b0000000000000000;
	sram_mem[95943] = 16'b0000000000000000;
	sram_mem[95944] = 16'b0000000000000000;
	sram_mem[95945] = 16'b0000000000000000;
	sram_mem[95946] = 16'b0000000000000000;
	sram_mem[95947] = 16'b0000000000000000;
	sram_mem[95948] = 16'b0000000000000000;
	sram_mem[95949] = 16'b0000000000000000;
	sram_mem[95950] = 16'b0000000000000000;
	sram_mem[95951] = 16'b0000000000000000;
	sram_mem[95952] = 16'b0000000000000000;
	sram_mem[95953] = 16'b0000000000000000;
	sram_mem[95954] = 16'b0000000000000000;
	sram_mem[95955] = 16'b0000000000000000;
	sram_mem[95956] = 16'b0000000000000000;
	sram_mem[95957] = 16'b0000000000000000;
	sram_mem[95958] = 16'b0000000000000000;
	sram_mem[95959] = 16'b0000000000000000;
	sram_mem[95960] = 16'b0000000000000000;
	sram_mem[95961] = 16'b0000000000000000;
	sram_mem[95962] = 16'b0000000000000000;
	sram_mem[95963] = 16'b0000000000000000;
	sram_mem[95964] = 16'b0000000000000000;
	sram_mem[95965] = 16'b0000000000000000;
	sram_mem[95966] = 16'b0000000000000000;
	sram_mem[95967] = 16'b0000000000000000;
	sram_mem[95968] = 16'b0000000000000000;
	sram_mem[95969] = 16'b0000000000000000;
	sram_mem[95970] = 16'b0000000000000000;
	sram_mem[95971] = 16'b0000000000000000;
	sram_mem[95972] = 16'b0000000000000000;
	sram_mem[95973] = 16'b0000000000000000;
	sram_mem[95974] = 16'b0000000000000000;
	sram_mem[95975] = 16'b0000000000000000;
	sram_mem[95976] = 16'b0000000000000000;
	sram_mem[95977] = 16'b0000000000000000;
	sram_mem[95978] = 16'b0000000000000000;
	sram_mem[95979] = 16'b0000000000000000;
	sram_mem[95980] = 16'b0000000000000000;
	sram_mem[95981] = 16'b0000000000000000;
	sram_mem[95982] = 16'b0000000000000000;
	sram_mem[95983] = 16'b0000000000000000;
	sram_mem[95984] = 16'b0000000000000000;
	sram_mem[95985] = 16'b0000000000000000;
	sram_mem[95986] = 16'b0000000000000000;
	sram_mem[95987] = 16'b0000000000000000;
	sram_mem[95988] = 16'b0000000000000000;
	sram_mem[95989] = 16'b0000000000000000;
	sram_mem[95990] = 16'b0000000000000000;
	sram_mem[95991] = 16'b0000000000000000;
	sram_mem[95992] = 16'b0000000000000000;
	sram_mem[95993] = 16'b0000000000000000;
	sram_mem[95994] = 16'b0000000000000000;
	sram_mem[95995] = 16'b0000000000000000;
	sram_mem[95996] = 16'b0000000000000000;
	sram_mem[95997] = 16'b0000000000000000;
	sram_mem[95998] = 16'b0000000000000000;
	sram_mem[95999] = 16'b0000000000000000;
	sram_mem[96000] = 16'b0000000000000000;
	sram_mem[96001] = 16'b0000000000000000;
	sram_mem[96002] = 16'b0000000000000000;
	sram_mem[96003] = 16'b0000000000000000;
	sram_mem[96004] = 16'b0000000000000000;
	sram_mem[96005] = 16'b0000000000000000;
	sram_mem[96006] = 16'b0000000000000000;
	sram_mem[96007] = 16'b0000000000000000;
	sram_mem[96008] = 16'b0000000000000000;
	sram_mem[96009] = 16'b0000000000000000;
	sram_mem[96010] = 16'b0000000000000000;
	sram_mem[96011] = 16'b0000000000000000;
	sram_mem[96012] = 16'b0000000000000000;
	sram_mem[96013] = 16'b0000000000000000;
	sram_mem[96014] = 16'b0000000000000000;
	sram_mem[96015] = 16'b0000000000000000;
	sram_mem[96016] = 16'b0000000000000000;
	sram_mem[96017] = 16'b0000000000000000;
	sram_mem[96018] = 16'b0000000000000000;
	sram_mem[96019] = 16'b0000000000000000;
	sram_mem[96020] = 16'b0000000000000000;
	sram_mem[96021] = 16'b0000000000000000;
	sram_mem[96022] = 16'b0000000000000000;
	sram_mem[96023] = 16'b0000000000000000;
	sram_mem[96024] = 16'b0000000000000000;
	sram_mem[96025] = 16'b0000000000000000;
	sram_mem[96026] = 16'b0000000000000000;
	sram_mem[96027] = 16'b0000000000000000;
	sram_mem[96028] = 16'b0000000000000000;
	sram_mem[96029] = 16'b0000000000000000;
	sram_mem[96030] = 16'b0000000000000000;
	sram_mem[96031] = 16'b0000000000000000;
	sram_mem[96032] = 16'b0000000000000000;
	sram_mem[96033] = 16'b0000000000000000;
	sram_mem[96034] = 16'b0000000000000000;
	sram_mem[96035] = 16'b0000000000000000;
	sram_mem[96036] = 16'b0000000000000000;
	sram_mem[96037] = 16'b0000000000000000;
	sram_mem[96038] = 16'b0000000000000000;
	sram_mem[96039] = 16'b0000000000000000;
	sram_mem[96040] = 16'b0000000000000000;
	sram_mem[96041] = 16'b0000000000000000;
	sram_mem[96042] = 16'b0000000000000000;
	sram_mem[96043] = 16'b0000000000000000;
	sram_mem[96044] = 16'b0000000000000000;
	sram_mem[96045] = 16'b0000000000000000;
	sram_mem[96046] = 16'b0000000000000000;
	sram_mem[96047] = 16'b0000000000000000;
	sram_mem[96048] = 16'b0000000000000000;
	sram_mem[96049] = 16'b0000000000000000;
	sram_mem[96050] = 16'b0000000000000000;
	sram_mem[96051] = 16'b0000000000000000;
	sram_mem[96052] = 16'b0000000000000000;
	sram_mem[96053] = 16'b0000000000000000;
	sram_mem[96054] = 16'b0000000000000000;
	sram_mem[96055] = 16'b0000000000000000;
	sram_mem[96056] = 16'b0000000000000000;
	sram_mem[96057] = 16'b0000000000000000;
	sram_mem[96058] = 16'b0000000000000000;
	sram_mem[96059] = 16'b0000000000000000;
	sram_mem[96060] = 16'b0000000000000000;
	sram_mem[96061] = 16'b0000000000000000;
	sram_mem[96062] = 16'b0000000000000000;
	sram_mem[96063] = 16'b0000000000000000;
	sram_mem[96064] = 16'b0000000000000000;
	sram_mem[96065] = 16'b0000000000000000;
	sram_mem[96066] = 16'b0000000000000000;
	sram_mem[96067] = 16'b0000000000000000;
	sram_mem[96068] = 16'b0000000000000000;
	sram_mem[96069] = 16'b0000000000000000;
	sram_mem[96070] = 16'b0000000000000000;
	sram_mem[96071] = 16'b0000000000000000;
	sram_mem[96072] = 16'b0000000000000000;
	sram_mem[96073] = 16'b0000000000000000;
	sram_mem[96074] = 16'b0000000000000000;
	sram_mem[96075] = 16'b0000000000000000;
	sram_mem[96076] = 16'b0000000000000000;
	sram_mem[96077] = 16'b0000000000000000;
	sram_mem[96078] = 16'b0000000000000000;
	sram_mem[96079] = 16'b0000000000000000;
	sram_mem[96080] = 16'b0000000000000000;
	sram_mem[96081] = 16'b0000000000000000;
	sram_mem[96082] = 16'b0000000000000000;
	sram_mem[96083] = 16'b0000000000000000;
	sram_mem[96084] = 16'b0000000000000000;
	sram_mem[96085] = 16'b0000000000000000;
	sram_mem[96086] = 16'b0000000000000000;
	sram_mem[96087] = 16'b0000000000000000;
	sram_mem[96088] = 16'b0000000000000000;
	sram_mem[96089] = 16'b0000000000000000;
	sram_mem[96090] = 16'b0000000000000000;
	sram_mem[96091] = 16'b0000000000000000;
	sram_mem[96092] = 16'b0000000000000000;
	sram_mem[96093] = 16'b0000000000000000;
	sram_mem[96094] = 16'b0000000000000000;
	sram_mem[96095] = 16'b0000000000000000;
	sram_mem[96096] = 16'b0000000000000000;
	sram_mem[96097] = 16'b0000000000000000;
	sram_mem[96098] = 16'b0000000000000000;
	sram_mem[96099] = 16'b0000000000000000;
	sram_mem[96100] = 16'b0000000000000000;
	sram_mem[96101] = 16'b0000000000000000;
	sram_mem[96102] = 16'b0000000000000000;
	sram_mem[96103] = 16'b0000000000000000;
	sram_mem[96104] = 16'b0000000000000000;
	sram_mem[96105] = 16'b0000000000000000;
	sram_mem[96106] = 16'b0000000000000000;
	sram_mem[96107] = 16'b0000000000000000;
	sram_mem[96108] = 16'b0000000000000000;
	sram_mem[96109] = 16'b0000000000000000;
	sram_mem[96110] = 16'b0000000000000000;
	sram_mem[96111] = 16'b0000000000000000;
	sram_mem[96112] = 16'b0000000000000000;
	sram_mem[96113] = 16'b0000000000000000;
	sram_mem[96114] = 16'b0000000000000000;
	sram_mem[96115] = 16'b0000000000000000;
	sram_mem[96116] = 16'b0000000000000000;
	sram_mem[96117] = 16'b0000000000000000;
	sram_mem[96118] = 16'b0000000000000000;
	sram_mem[96119] = 16'b0000000000000000;
	sram_mem[96120] = 16'b0000000000000000;
	sram_mem[96121] = 16'b0000000000000000;
	sram_mem[96122] = 16'b0000000000000000;
	sram_mem[96123] = 16'b0000000000000000;
	sram_mem[96124] = 16'b0000000000000000;
	sram_mem[96125] = 16'b0000000000000000;
	sram_mem[96126] = 16'b0000000000000000;
	sram_mem[96127] = 16'b0000000000000000;
	sram_mem[96128] = 16'b0000000000000000;
	sram_mem[96129] = 16'b0000000000000000;
	sram_mem[96130] = 16'b0000000000000000;
	sram_mem[96131] = 16'b0000000000000000;
	sram_mem[96132] = 16'b0000000000000000;
	sram_mem[96133] = 16'b0000000000000000;
	sram_mem[96134] = 16'b0000000000000000;
	sram_mem[96135] = 16'b0000000000000000;
	sram_mem[96136] = 16'b0000000000000000;
	sram_mem[96137] = 16'b0000000000000000;
	sram_mem[96138] = 16'b0000000000000000;
	sram_mem[96139] = 16'b0000000000000000;
	sram_mem[96140] = 16'b0000000000000000;
	sram_mem[96141] = 16'b0000000000000000;
	sram_mem[96142] = 16'b0000000000000000;
	sram_mem[96143] = 16'b0000000000000000;
	sram_mem[96144] = 16'b0000000000000000;
	sram_mem[96145] = 16'b0000000000000000;
	sram_mem[96146] = 16'b0000000000000000;
	sram_mem[96147] = 16'b0000000000000000;
	sram_mem[96148] = 16'b0000000000000000;
	sram_mem[96149] = 16'b0000000000000000;
	sram_mem[96150] = 16'b0000000000000000;
	sram_mem[96151] = 16'b0000000000000000;
	sram_mem[96152] = 16'b0000000000000000;
	sram_mem[96153] = 16'b0000000000000000;
	sram_mem[96154] = 16'b0000000000000000;
	sram_mem[96155] = 16'b0000000000000000;
	sram_mem[96156] = 16'b0000000000000000;
	sram_mem[96157] = 16'b0000000000000000;
	sram_mem[96158] = 16'b0000000000000000;
	sram_mem[96159] = 16'b0000000000000000;
	sram_mem[96160] = 16'b0000000000000000;
	sram_mem[96161] = 16'b0000000000000000;
	sram_mem[96162] = 16'b0000000000000000;
	sram_mem[96163] = 16'b0000000000000000;
	sram_mem[96164] = 16'b0000000000000000;
	sram_mem[96165] = 16'b0000000000000000;
	sram_mem[96166] = 16'b0000000000000000;
	sram_mem[96167] = 16'b0000000000000000;
	sram_mem[96168] = 16'b0000000000000000;
	sram_mem[96169] = 16'b0000000000000000;
	sram_mem[96170] = 16'b0000000000000000;
	sram_mem[96171] = 16'b0000000000000000;
	sram_mem[96172] = 16'b0000000000000000;
	sram_mem[96173] = 16'b0000000000000000;
	sram_mem[96174] = 16'b0000000000000000;
	sram_mem[96175] = 16'b0000000000000000;
	sram_mem[96176] = 16'b0000000000000000;
	sram_mem[96177] = 16'b0000000000000000;
	sram_mem[96178] = 16'b0000000000000000;
	sram_mem[96179] = 16'b0000000000000000;
	sram_mem[96180] = 16'b0000000000000000;
	sram_mem[96181] = 16'b0000000000000000;
	sram_mem[96182] = 16'b0000000000000000;
	sram_mem[96183] = 16'b0000000000000000;
	sram_mem[96184] = 16'b0000000000000000;
	sram_mem[96185] = 16'b0000000000000000;
	sram_mem[96186] = 16'b0000000000000000;
	sram_mem[96187] = 16'b0000000000000000;
	sram_mem[96188] = 16'b0000000000000000;
	sram_mem[96189] = 16'b0000000000000000;
	sram_mem[96190] = 16'b0000000000000000;
	sram_mem[96191] = 16'b0000000000000000;
	sram_mem[96192] = 16'b0000000000000000;
	sram_mem[96193] = 16'b0000000000000000;
	sram_mem[96194] = 16'b0000000000000000;
	sram_mem[96195] = 16'b0000000000000000;
	sram_mem[96196] = 16'b0000000000000000;
	sram_mem[96197] = 16'b0000000000000000;
	sram_mem[96198] = 16'b0000000000000000;
	sram_mem[96199] = 16'b0000000000000000;
	sram_mem[96200] = 16'b0000000000000000;
	sram_mem[96201] = 16'b0000000000000000;
	sram_mem[96202] = 16'b0000000000000000;
	sram_mem[96203] = 16'b0000000000000000;
	sram_mem[96204] = 16'b0000000000000000;
	sram_mem[96205] = 16'b0000000000000000;
	sram_mem[96206] = 16'b0000000000000000;
	sram_mem[96207] = 16'b0000000000000000;
	sram_mem[96208] = 16'b0000000000000000;
	sram_mem[96209] = 16'b0000000000000000;
	sram_mem[96210] = 16'b0000000000000000;
	sram_mem[96211] = 16'b0000000000000000;
	sram_mem[96212] = 16'b0000000000000000;
	sram_mem[96213] = 16'b0000000000000000;
	sram_mem[96214] = 16'b0000000000000000;
	sram_mem[96215] = 16'b0000000000000000;
	sram_mem[96216] = 16'b0000000000000000;
	sram_mem[96217] = 16'b0000000000000000;
	sram_mem[96218] = 16'b0000000000000000;
	sram_mem[96219] = 16'b0000000000000000;
	sram_mem[96220] = 16'b0000000000000000;
	sram_mem[96221] = 16'b0000000000000000;
	sram_mem[96222] = 16'b0000000000000000;
	sram_mem[96223] = 16'b0000000000000000;
	sram_mem[96224] = 16'b0000000000000000;
	sram_mem[96225] = 16'b0000000000000000;
	sram_mem[96226] = 16'b0000000000000000;
	sram_mem[96227] = 16'b0000000000000000;
	sram_mem[96228] = 16'b0000000000000000;
	sram_mem[96229] = 16'b0000000000000000;
	sram_mem[96230] = 16'b0000000000000000;
	sram_mem[96231] = 16'b0000000000000000;
	sram_mem[96232] = 16'b0000000000000000;
	sram_mem[96233] = 16'b0000000000000000;
	sram_mem[96234] = 16'b0000000000000000;
	sram_mem[96235] = 16'b0000000000000000;
	sram_mem[96236] = 16'b0000000000000000;
	sram_mem[96237] = 16'b0000000000000000;
	sram_mem[96238] = 16'b0000000000000000;
	sram_mem[96239] = 16'b0000000000000000;
	sram_mem[96240] = 16'b0000000000000000;
	sram_mem[96241] = 16'b0000000000000000;
	sram_mem[96242] = 16'b0000000000000000;
	sram_mem[96243] = 16'b0000000000000000;
	sram_mem[96244] = 16'b0000000000000000;
	sram_mem[96245] = 16'b0000000000000000;
	sram_mem[96246] = 16'b0000000000000000;
	sram_mem[96247] = 16'b0000000000000000;
	sram_mem[96248] = 16'b0000000000000000;
	sram_mem[96249] = 16'b0000000000000000;
	sram_mem[96250] = 16'b0000000000000000;
	sram_mem[96251] = 16'b0000000000000000;
	sram_mem[96252] = 16'b0000000000000000;
	sram_mem[96253] = 16'b0000000000000000;
	sram_mem[96254] = 16'b0000000000000000;
	sram_mem[96255] = 16'b0000000000000000;
	sram_mem[96256] = 16'b0000000000000000;
	sram_mem[96257] = 16'b0000000000000000;
	sram_mem[96258] = 16'b0000000000000000;
	sram_mem[96259] = 16'b0000000000000000;
	sram_mem[96260] = 16'b0000000000000000;
	sram_mem[96261] = 16'b0000000000000000;
	sram_mem[96262] = 16'b0000000000000000;
	sram_mem[96263] = 16'b0000000000000000;
	sram_mem[96264] = 16'b0000000000000000;
	sram_mem[96265] = 16'b0000000000000000;
	sram_mem[96266] = 16'b0000000000000000;
	sram_mem[96267] = 16'b0000000000000000;
	sram_mem[96268] = 16'b0000000000000000;
	sram_mem[96269] = 16'b0000000000000000;
	sram_mem[96270] = 16'b0000000000000000;
	sram_mem[96271] = 16'b0000000000000000;
	sram_mem[96272] = 16'b0000000000000000;
	sram_mem[96273] = 16'b0000000000000000;
	sram_mem[96274] = 16'b0000000000000000;
	sram_mem[96275] = 16'b0000000000000000;
	sram_mem[96276] = 16'b0000000000000000;
	sram_mem[96277] = 16'b0000000000000000;
	sram_mem[96278] = 16'b0000000000000000;
	sram_mem[96279] = 16'b0000000000000000;
	sram_mem[96280] = 16'b0000000000000000;
	sram_mem[96281] = 16'b0000000000000000;
	sram_mem[96282] = 16'b0000000000000000;
	sram_mem[96283] = 16'b0000000000000000;
	sram_mem[96284] = 16'b0000000000000000;
	sram_mem[96285] = 16'b0000000000000000;
	sram_mem[96286] = 16'b0000000000000000;
	sram_mem[96287] = 16'b0000000000000000;
	sram_mem[96288] = 16'b0000000000000000;
	sram_mem[96289] = 16'b0000000000000000;
	sram_mem[96290] = 16'b0000000000000000;
	sram_mem[96291] = 16'b0000000000000000;
	sram_mem[96292] = 16'b0000000000000000;
	sram_mem[96293] = 16'b0000000000000000;
	sram_mem[96294] = 16'b0000000000000000;
	sram_mem[96295] = 16'b0000000000000000;
	sram_mem[96296] = 16'b0000000000000000;
	sram_mem[96297] = 16'b0000000000000000;
	sram_mem[96298] = 16'b0000000000000000;
	sram_mem[96299] = 16'b0000000000000000;
	sram_mem[96300] = 16'b0000000000000000;
	sram_mem[96301] = 16'b0000000000000000;
	sram_mem[96302] = 16'b0000000000000000;
	sram_mem[96303] = 16'b0000000000000000;
	sram_mem[96304] = 16'b0000000000000000;
	sram_mem[96305] = 16'b0000000000000000;
	sram_mem[96306] = 16'b0000000000000000;
	sram_mem[96307] = 16'b0000000000000000;
	sram_mem[96308] = 16'b0000000000000000;
	sram_mem[96309] = 16'b0000000000000000;
	sram_mem[96310] = 16'b0000000000000000;
	sram_mem[96311] = 16'b0000000000000000;
	sram_mem[96312] = 16'b0000000000000000;
	sram_mem[96313] = 16'b0000000000000000;
	sram_mem[96314] = 16'b0000000000000000;
	sram_mem[96315] = 16'b0000000000000000;
	sram_mem[96316] = 16'b0000000000000000;
	sram_mem[96317] = 16'b0000000000000000;
	sram_mem[96318] = 16'b0000000000000000;
	sram_mem[96319] = 16'b0000000000000000;
	sram_mem[96320] = 16'b0000000000000000;
	sram_mem[96321] = 16'b0000000000000000;
	sram_mem[96322] = 16'b0000000000000000;
	sram_mem[96323] = 16'b0000000000000000;
	sram_mem[96324] = 16'b0000000000000000;
	sram_mem[96325] = 16'b0000000000000000;
	sram_mem[96326] = 16'b0000000000000000;
	sram_mem[96327] = 16'b0000000000000000;
	sram_mem[96328] = 16'b0000000000000000;
	sram_mem[96329] = 16'b0000000000000000;
	sram_mem[96330] = 16'b0000000000000000;
	sram_mem[96331] = 16'b0000000000000000;
	sram_mem[96332] = 16'b0000000000000000;
	sram_mem[96333] = 16'b0000000000000000;
	sram_mem[96334] = 16'b0000000000000000;
	sram_mem[96335] = 16'b0000000000000000;
	sram_mem[96336] = 16'b0000000000000000;
	sram_mem[96337] = 16'b0000000000000000;
	sram_mem[96338] = 16'b0000000000000000;
	sram_mem[96339] = 16'b0000000000000000;
	sram_mem[96340] = 16'b0000000000000000;
	sram_mem[96341] = 16'b0000000000000000;
	sram_mem[96342] = 16'b0000000000000000;
	sram_mem[96343] = 16'b0000000000000000;
	sram_mem[96344] = 16'b0000000000000000;
	sram_mem[96345] = 16'b0000000000000000;
	sram_mem[96346] = 16'b0000000000000000;
	sram_mem[96347] = 16'b0000000000000000;
	sram_mem[96348] = 16'b0000000000000000;
	sram_mem[96349] = 16'b0000000000000000;
	sram_mem[96350] = 16'b0000000000000000;
	sram_mem[96351] = 16'b0000000000000000;
	sram_mem[96352] = 16'b0000000000000000;
	sram_mem[96353] = 16'b0000000000000000;
	sram_mem[96354] = 16'b0000000000000000;
	sram_mem[96355] = 16'b0000000000000000;
	sram_mem[96356] = 16'b0000000000000000;
	sram_mem[96357] = 16'b0000000000000000;
	sram_mem[96358] = 16'b0000000000000000;
	sram_mem[96359] = 16'b0000000000000000;
	sram_mem[96360] = 16'b0000000000000000;
	sram_mem[96361] = 16'b0000000000000000;
	sram_mem[96362] = 16'b0000000000000000;
	sram_mem[96363] = 16'b0000000000000000;
	sram_mem[96364] = 16'b0000000000000000;
	sram_mem[96365] = 16'b0000000000000000;
	sram_mem[96366] = 16'b0000000000000000;
	sram_mem[96367] = 16'b0000000000000000;
	sram_mem[96368] = 16'b0000000000000000;
	sram_mem[96369] = 16'b0000000000000000;
	sram_mem[96370] = 16'b0000000000000000;
	sram_mem[96371] = 16'b0000000000000000;
	sram_mem[96372] = 16'b0000000000000000;
	sram_mem[96373] = 16'b0000000000000000;
	sram_mem[96374] = 16'b0000000000000000;
	sram_mem[96375] = 16'b0000000000000000;
	sram_mem[96376] = 16'b0000000000000000;
	sram_mem[96377] = 16'b0000000000000000;
	sram_mem[96378] = 16'b0000000000000000;
	sram_mem[96379] = 16'b0000000000000000;
	sram_mem[96380] = 16'b0000000000000000;
	sram_mem[96381] = 16'b0000000000000000;
	sram_mem[96382] = 16'b0000000000000000;
	sram_mem[96383] = 16'b0000000000000000;
	sram_mem[96384] = 16'b0000000000000000;
	sram_mem[96385] = 16'b0000000000000000;
	sram_mem[96386] = 16'b0000000000000000;
	sram_mem[96387] = 16'b0000000000000000;
	sram_mem[96388] = 16'b0000000000000000;
	sram_mem[96389] = 16'b0000000000000000;
	sram_mem[96390] = 16'b0000000000000000;
	sram_mem[96391] = 16'b0000000000000000;
	sram_mem[96392] = 16'b0000000000000000;
	sram_mem[96393] = 16'b0000000000000000;
	sram_mem[96394] = 16'b0000000000000000;
	sram_mem[96395] = 16'b0000000000000000;
	sram_mem[96396] = 16'b0000000000000000;
	sram_mem[96397] = 16'b0000000000000000;
	sram_mem[96398] = 16'b0000000000000000;
	sram_mem[96399] = 16'b0000000000000000;
	sram_mem[96400] = 16'b0000000000000000;
	sram_mem[96401] = 16'b0000000000000000;
	sram_mem[96402] = 16'b0000000000000000;
	sram_mem[96403] = 16'b0000000000000000;
	sram_mem[96404] = 16'b0000000000000000;
	sram_mem[96405] = 16'b0000000000000000;
	sram_mem[96406] = 16'b0000000000000000;
	sram_mem[96407] = 16'b0000000000000000;
	sram_mem[96408] = 16'b0000000000000000;
	sram_mem[96409] = 16'b0000000000000000;
	sram_mem[96410] = 16'b0000000000000000;
	sram_mem[96411] = 16'b0000000000000000;
	sram_mem[96412] = 16'b0000000000000000;
	sram_mem[96413] = 16'b0000000000000000;
	sram_mem[96414] = 16'b0000000000000000;
	sram_mem[96415] = 16'b0000000000000000;
	sram_mem[96416] = 16'b0000000000000000;
	sram_mem[96417] = 16'b0000000000000000;
	sram_mem[96418] = 16'b0000000000000000;
	sram_mem[96419] = 16'b0000000000000000;
	sram_mem[96420] = 16'b0000000000000000;
	sram_mem[96421] = 16'b0000000000000000;
	sram_mem[96422] = 16'b0000000000000000;
	sram_mem[96423] = 16'b0000000000000000;
	sram_mem[96424] = 16'b0000000000000000;
	sram_mem[96425] = 16'b0000000000000000;
	sram_mem[96426] = 16'b0000000000000000;
	sram_mem[96427] = 16'b0000000000000000;
	sram_mem[96428] = 16'b0000000000000000;
	sram_mem[96429] = 16'b0000000000000000;
	sram_mem[96430] = 16'b0000000000000000;
	sram_mem[96431] = 16'b0000000000000000;
	sram_mem[96432] = 16'b0000000000000000;
	sram_mem[96433] = 16'b0000000000000000;
	sram_mem[96434] = 16'b0000000000000000;
	sram_mem[96435] = 16'b0000000000000000;
	sram_mem[96436] = 16'b0000000000000000;
	sram_mem[96437] = 16'b0000000000000000;
	sram_mem[96438] = 16'b0000000000000000;
	sram_mem[96439] = 16'b0000000000000000;
	sram_mem[96440] = 16'b0000000000000000;
	sram_mem[96441] = 16'b0000000000000000;
	sram_mem[96442] = 16'b0000000000000000;
	sram_mem[96443] = 16'b0000000000000000;
	sram_mem[96444] = 16'b0000000000000000;
	sram_mem[96445] = 16'b0000000000000000;
	sram_mem[96446] = 16'b0000000000000000;
	sram_mem[96447] = 16'b0000000000000000;
	sram_mem[96448] = 16'b0000000000000000;
	sram_mem[96449] = 16'b0000000000000000;
	sram_mem[96450] = 16'b0000000000000000;
	sram_mem[96451] = 16'b0000000000000000;
	sram_mem[96452] = 16'b0000000000000000;
	sram_mem[96453] = 16'b0000000000000000;
	sram_mem[96454] = 16'b0000000000000000;
	sram_mem[96455] = 16'b0000000000000000;
	sram_mem[96456] = 16'b0000000000000000;
	sram_mem[96457] = 16'b0000000000000000;
	sram_mem[96458] = 16'b0000000000000000;
	sram_mem[96459] = 16'b0000000000000000;
	sram_mem[96460] = 16'b0000000000000000;
	sram_mem[96461] = 16'b0000000000000000;
	sram_mem[96462] = 16'b0000000000000000;
	sram_mem[96463] = 16'b0000000000000000;
	sram_mem[96464] = 16'b0000000000000000;
	sram_mem[96465] = 16'b0000000000000000;
	sram_mem[96466] = 16'b0000000000000000;
	sram_mem[96467] = 16'b0000000000000000;
	sram_mem[96468] = 16'b0000000000000000;
	sram_mem[96469] = 16'b0000000000000000;
	sram_mem[96470] = 16'b0000000000000000;
	sram_mem[96471] = 16'b0000000000000000;
	sram_mem[96472] = 16'b0000000000000000;
	sram_mem[96473] = 16'b0000000000000000;
	sram_mem[96474] = 16'b0000000000000000;
	sram_mem[96475] = 16'b0000000000000000;
	sram_mem[96476] = 16'b0000000000000000;
	sram_mem[96477] = 16'b0000000000000000;
	sram_mem[96478] = 16'b0000000000000000;
	sram_mem[96479] = 16'b0000000000000000;
	sram_mem[96480] = 16'b0000000000000000;
	sram_mem[96481] = 16'b0000000000000000;
	sram_mem[96482] = 16'b0000000000000000;
	sram_mem[96483] = 16'b0000000000000000;
	sram_mem[96484] = 16'b0000000000000000;
	sram_mem[96485] = 16'b0000000000000000;
	sram_mem[96486] = 16'b0000000000000000;
	sram_mem[96487] = 16'b0000000000000000;
	sram_mem[96488] = 16'b0000000000000000;
	sram_mem[96489] = 16'b0000000000000000;
	sram_mem[96490] = 16'b0000000000000000;
	sram_mem[96491] = 16'b0000000000000000;
	sram_mem[96492] = 16'b0000000000000000;
	sram_mem[96493] = 16'b0000000000000000;
	sram_mem[96494] = 16'b0000000000000000;
	sram_mem[96495] = 16'b0000000000000000;
	sram_mem[96496] = 16'b0000000000000000;
	sram_mem[96497] = 16'b0000000000000000;
	sram_mem[96498] = 16'b0000000000000000;
	sram_mem[96499] = 16'b0000000000000000;
	sram_mem[96500] = 16'b0000000000000000;
	sram_mem[96501] = 16'b0000000000000000;
	sram_mem[96502] = 16'b0000000000000000;
	sram_mem[96503] = 16'b0000000000000000;
	sram_mem[96504] = 16'b0000000000000000;
	sram_mem[96505] = 16'b0000000000000000;
	sram_mem[96506] = 16'b0000000000000000;
	sram_mem[96507] = 16'b0000000000000000;
	sram_mem[96508] = 16'b0000000000000000;
	sram_mem[96509] = 16'b0000000000000000;
	sram_mem[96510] = 16'b0000000000000000;
	sram_mem[96511] = 16'b0000000000000000;
	sram_mem[96512] = 16'b0000000000000000;
	sram_mem[96513] = 16'b0000000000000000;
	sram_mem[96514] = 16'b0000000000000000;
	sram_mem[96515] = 16'b0000000000000000;
	sram_mem[96516] = 16'b0000000000000000;
	sram_mem[96517] = 16'b0000000000000000;
	sram_mem[96518] = 16'b0000000000000000;
	sram_mem[96519] = 16'b0000000000000000;
	sram_mem[96520] = 16'b0000000000000000;
	sram_mem[96521] = 16'b0000000000000000;
	sram_mem[96522] = 16'b0000000000000000;
	sram_mem[96523] = 16'b0000000000000000;
	sram_mem[96524] = 16'b0000000000000000;
	sram_mem[96525] = 16'b0000000000000000;
	sram_mem[96526] = 16'b0000000000000000;
	sram_mem[96527] = 16'b0000000000000000;
	sram_mem[96528] = 16'b0000000000000000;
	sram_mem[96529] = 16'b0000000000000000;
	sram_mem[96530] = 16'b0000000000000000;
	sram_mem[96531] = 16'b0000000000000000;
	sram_mem[96532] = 16'b0000000000000000;
	sram_mem[96533] = 16'b0000000000000000;
	sram_mem[96534] = 16'b0000000000000000;
	sram_mem[96535] = 16'b0000000000000000;
	sram_mem[96536] = 16'b0000000000000000;
	sram_mem[96537] = 16'b0000000000000000;
	sram_mem[96538] = 16'b0000000000000000;
	sram_mem[96539] = 16'b0000000000000000;
	sram_mem[96540] = 16'b0000000000000000;
	sram_mem[96541] = 16'b0000000000000000;
	sram_mem[96542] = 16'b0000000000000000;
	sram_mem[96543] = 16'b0000000000000000;
	sram_mem[96544] = 16'b0000000000000000;
	sram_mem[96545] = 16'b0000000000000000;
	sram_mem[96546] = 16'b0000000000000000;
	sram_mem[96547] = 16'b0000000000000000;
	sram_mem[96548] = 16'b0000000000000000;
	sram_mem[96549] = 16'b0000000000000000;
	sram_mem[96550] = 16'b0000000000000000;
	sram_mem[96551] = 16'b0000000000000000;
	sram_mem[96552] = 16'b0000000000000000;
	sram_mem[96553] = 16'b0000000000000000;
	sram_mem[96554] = 16'b0000000000000000;
	sram_mem[96555] = 16'b0000000000000000;
	sram_mem[96556] = 16'b0000000000000000;
	sram_mem[96557] = 16'b0000000000000000;
	sram_mem[96558] = 16'b0000000000000000;
	sram_mem[96559] = 16'b0000000000000000;
	sram_mem[96560] = 16'b0000000000000000;
	sram_mem[96561] = 16'b0000000000000000;
	sram_mem[96562] = 16'b0000000000000000;
	sram_mem[96563] = 16'b0000000000000000;
	sram_mem[96564] = 16'b0000000000000000;
	sram_mem[96565] = 16'b0000000000000000;
	sram_mem[96566] = 16'b0000000000000000;
	sram_mem[96567] = 16'b0000000000000000;
	sram_mem[96568] = 16'b0000000000000000;
	sram_mem[96569] = 16'b0000000000000000;
	sram_mem[96570] = 16'b0000000000000000;
	sram_mem[96571] = 16'b0000000000000000;
	sram_mem[96572] = 16'b0000000000000000;
	sram_mem[96573] = 16'b0000000000000000;
	sram_mem[96574] = 16'b0000000000000000;
	sram_mem[96575] = 16'b0000000000000000;
	sram_mem[96576] = 16'b0000000000000000;
	sram_mem[96577] = 16'b0000000000000000;
	sram_mem[96578] = 16'b0000000000000000;
	sram_mem[96579] = 16'b0000000000000000;
	sram_mem[96580] = 16'b0000000000000000;
	sram_mem[96581] = 16'b0000000000000000;
	sram_mem[96582] = 16'b0000000000000000;
	sram_mem[96583] = 16'b0000000000000000;
	sram_mem[96584] = 16'b0000000000000000;
	sram_mem[96585] = 16'b0000000000000000;
	sram_mem[96586] = 16'b0000000000000000;
	sram_mem[96587] = 16'b0000000000000000;
	sram_mem[96588] = 16'b0000000000000000;
	sram_mem[96589] = 16'b0000000000000000;
	sram_mem[96590] = 16'b0000000000000000;
	sram_mem[96591] = 16'b0000000000000000;
	sram_mem[96592] = 16'b0000000000000000;
	sram_mem[96593] = 16'b0000000000000000;
	sram_mem[96594] = 16'b0000000000000000;
	sram_mem[96595] = 16'b0000000000000000;
	sram_mem[96596] = 16'b0000000000000000;
	sram_mem[96597] = 16'b0000000000000000;
	sram_mem[96598] = 16'b0000000000000000;
	sram_mem[96599] = 16'b0000000000000000;
	sram_mem[96600] = 16'b0000000000000000;
	sram_mem[96601] = 16'b0000000000000000;
	sram_mem[96602] = 16'b0000000000000000;
	sram_mem[96603] = 16'b0000000000000000;
	sram_mem[96604] = 16'b0000000000000000;
	sram_mem[96605] = 16'b0000000000000000;
	sram_mem[96606] = 16'b0000000000000000;
	sram_mem[96607] = 16'b0000000000000000;
	sram_mem[96608] = 16'b0000000000000000;
	sram_mem[96609] = 16'b0000000000000000;
	sram_mem[96610] = 16'b0000000000000000;
	sram_mem[96611] = 16'b0000000000000000;
	sram_mem[96612] = 16'b0000000000000000;
	sram_mem[96613] = 16'b0000000000000000;
	sram_mem[96614] = 16'b0000000000000000;
	sram_mem[96615] = 16'b0000000000000000;
	sram_mem[96616] = 16'b0000000000000000;
	sram_mem[96617] = 16'b0000000000000000;
	sram_mem[96618] = 16'b0000000000000000;
	sram_mem[96619] = 16'b0000000000000000;
	sram_mem[96620] = 16'b0000000000000000;
	sram_mem[96621] = 16'b0000000000000000;
	sram_mem[96622] = 16'b0000000000000000;
	sram_mem[96623] = 16'b0000000000000000;
	sram_mem[96624] = 16'b0000000000000000;
	sram_mem[96625] = 16'b0000000000000000;
	sram_mem[96626] = 16'b0000000000000000;
	sram_mem[96627] = 16'b0000000000000000;
	sram_mem[96628] = 16'b0000000000000000;
	sram_mem[96629] = 16'b0000000000000000;
	sram_mem[96630] = 16'b0000000000000000;
	sram_mem[96631] = 16'b0000000000000000;
	sram_mem[96632] = 16'b0000000000000000;
	sram_mem[96633] = 16'b0000000000000000;
	sram_mem[96634] = 16'b0000000000000000;
	sram_mem[96635] = 16'b0000000000000000;
	sram_mem[96636] = 16'b0000000000000000;
	sram_mem[96637] = 16'b0000000000000000;
	sram_mem[96638] = 16'b0000000000000000;
	sram_mem[96639] = 16'b0000000000000000;
	sram_mem[96640] = 16'b0000000000000000;
	sram_mem[96641] = 16'b0000000000000000;
	sram_mem[96642] = 16'b0000000000000000;
	sram_mem[96643] = 16'b0000000000000000;
	sram_mem[96644] = 16'b0000000000000000;
	sram_mem[96645] = 16'b0000000000000000;
	sram_mem[96646] = 16'b0000000000000000;
	sram_mem[96647] = 16'b0000000000000000;
	sram_mem[96648] = 16'b0000000000000000;
	sram_mem[96649] = 16'b0000000000000000;
	sram_mem[96650] = 16'b0000000000000000;
	sram_mem[96651] = 16'b0000000000000000;
	sram_mem[96652] = 16'b0000000000000000;
	sram_mem[96653] = 16'b0000000000000000;
	sram_mem[96654] = 16'b0000000000000000;
	sram_mem[96655] = 16'b0000000000000000;
	sram_mem[96656] = 16'b0000000000000000;
	sram_mem[96657] = 16'b0000000000000000;
	sram_mem[96658] = 16'b0000000000000000;
	sram_mem[96659] = 16'b0000000000000000;
	sram_mem[96660] = 16'b0000000000000000;
	sram_mem[96661] = 16'b0000000000000000;
	sram_mem[96662] = 16'b0000000000000000;
	sram_mem[96663] = 16'b0000000000000000;
	sram_mem[96664] = 16'b0000000000000000;
	sram_mem[96665] = 16'b0000000000000000;
	sram_mem[96666] = 16'b0000000000000000;
	sram_mem[96667] = 16'b0000000000000000;
	sram_mem[96668] = 16'b0000000000000000;
	sram_mem[96669] = 16'b0000000000000000;
	sram_mem[96670] = 16'b0000000000000000;
	sram_mem[96671] = 16'b0000000000000000;
	sram_mem[96672] = 16'b0000000000000000;
	sram_mem[96673] = 16'b0000000000000000;
	sram_mem[96674] = 16'b0000000000000000;
	sram_mem[96675] = 16'b0000000000000000;
	sram_mem[96676] = 16'b0000000000000000;
	sram_mem[96677] = 16'b0000000000000000;
	sram_mem[96678] = 16'b0000000000000000;
	sram_mem[96679] = 16'b0000000000000000;
	sram_mem[96680] = 16'b0000000000000000;
	sram_mem[96681] = 16'b0000000000000000;
	sram_mem[96682] = 16'b0000000000000000;
	sram_mem[96683] = 16'b0000000000000000;
	sram_mem[96684] = 16'b0000000000000000;
	sram_mem[96685] = 16'b0000000000000000;
	sram_mem[96686] = 16'b0000000000000000;
	sram_mem[96687] = 16'b0000000000000000;
	sram_mem[96688] = 16'b0000000000000000;
	sram_mem[96689] = 16'b0000000000000000;
	sram_mem[96690] = 16'b0000000000000000;
	sram_mem[96691] = 16'b0000000000000000;
	sram_mem[96692] = 16'b0000000000000000;
	sram_mem[96693] = 16'b0000000000000000;
	sram_mem[96694] = 16'b0000000000000000;
	sram_mem[96695] = 16'b0000000000000000;
	sram_mem[96696] = 16'b0000000000000000;
	sram_mem[96697] = 16'b0000000000000000;
	sram_mem[96698] = 16'b0000000000000000;
	sram_mem[96699] = 16'b0000000000000000;
	sram_mem[96700] = 16'b0000000000000000;
	sram_mem[96701] = 16'b0000000000000000;
	sram_mem[96702] = 16'b0000000000000000;
	sram_mem[96703] = 16'b0000000000000000;
	sram_mem[96704] = 16'b0000000000000000;
	sram_mem[96705] = 16'b0000000000000000;
	sram_mem[96706] = 16'b0000000000000000;
	sram_mem[96707] = 16'b0000000000000000;
	sram_mem[96708] = 16'b0000000000000000;
	sram_mem[96709] = 16'b0000000000000000;
	sram_mem[96710] = 16'b0000000000000000;
	sram_mem[96711] = 16'b0000000000000000;
	sram_mem[96712] = 16'b0000000000000000;
	sram_mem[96713] = 16'b0000000000000000;
	sram_mem[96714] = 16'b0000000000000000;
	sram_mem[96715] = 16'b0000000000000000;
	sram_mem[96716] = 16'b0000000000000000;
	sram_mem[96717] = 16'b0000000000000000;
	sram_mem[96718] = 16'b0000000000000000;
	sram_mem[96719] = 16'b0000000000000000;
	sram_mem[96720] = 16'b0000000000000000;
	sram_mem[96721] = 16'b0000000000000000;
	sram_mem[96722] = 16'b0000000000000000;
	sram_mem[96723] = 16'b0000000000000000;
	sram_mem[96724] = 16'b0000000000000000;
	sram_mem[96725] = 16'b0000000000000000;
	sram_mem[96726] = 16'b0000000000000000;
	sram_mem[96727] = 16'b0000000000000000;
	sram_mem[96728] = 16'b0000000000000000;
	sram_mem[96729] = 16'b0000000000000000;
	sram_mem[96730] = 16'b0000000000000000;
	sram_mem[96731] = 16'b0000000000000000;
	sram_mem[96732] = 16'b0000000000000000;
	sram_mem[96733] = 16'b0000000000000000;
	sram_mem[96734] = 16'b0000000000000000;
	sram_mem[96735] = 16'b0000000000000000;
	sram_mem[96736] = 16'b0000000000000000;
	sram_mem[96737] = 16'b0000000000000000;
	sram_mem[96738] = 16'b0000000000000000;
	sram_mem[96739] = 16'b0000000000000000;
	sram_mem[96740] = 16'b0000000000000000;
	sram_mem[96741] = 16'b0000000000000000;
	sram_mem[96742] = 16'b0000000000000000;
	sram_mem[96743] = 16'b0000000000000000;
	sram_mem[96744] = 16'b0000000000000000;
	sram_mem[96745] = 16'b0000000000000000;
	sram_mem[96746] = 16'b0000000000000000;
	sram_mem[96747] = 16'b0000000000000000;
	sram_mem[96748] = 16'b0000000000000000;
	sram_mem[96749] = 16'b0000000000000000;
	sram_mem[96750] = 16'b0000000000000000;
	sram_mem[96751] = 16'b0000000000000000;
	sram_mem[96752] = 16'b0000000000000000;
	sram_mem[96753] = 16'b0000000000000000;
	sram_mem[96754] = 16'b0000000000000000;
	sram_mem[96755] = 16'b0000000000000000;
	sram_mem[96756] = 16'b0000000000000000;
	sram_mem[96757] = 16'b0000000000000000;
	sram_mem[96758] = 16'b0000000000000000;
	sram_mem[96759] = 16'b0000000000000000;
	sram_mem[96760] = 16'b0000000000000000;
	sram_mem[96761] = 16'b0000000000000000;
	sram_mem[96762] = 16'b0000000000000000;
	sram_mem[96763] = 16'b0000000000000000;
	sram_mem[96764] = 16'b0000000000000000;
	sram_mem[96765] = 16'b0000000000000000;
	sram_mem[96766] = 16'b0000000000000000;
	sram_mem[96767] = 16'b0000000000000000;
	sram_mem[96768] = 16'b0000000000000000;
	sram_mem[96769] = 16'b0000000000000000;
	sram_mem[96770] = 16'b0000000000000000;
	sram_mem[96771] = 16'b0000000000000000;
	sram_mem[96772] = 16'b0000000000000000;
	sram_mem[96773] = 16'b0000000000000000;
	sram_mem[96774] = 16'b0000000000000000;
	sram_mem[96775] = 16'b0000000000000000;
	sram_mem[96776] = 16'b0000000000000000;
	sram_mem[96777] = 16'b0000000000000000;
	sram_mem[96778] = 16'b0000000000000000;
	sram_mem[96779] = 16'b0000000000000000;
	sram_mem[96780] = 16'b0000000000000000;
	sram_mem[96781] = 16'b0000000000000000;
	sram_mem[96782] = 16'b0000000000000000;
	sram_mem[96783] = 16'b0000000000000000;
	sram_mem[96784] = 16'b0000000000000000;
	sram_mem[96785] = 16'b0000000000000000;
	sram_mem[96786] = 16'b0000000000000000;
	sram_mem[96787] = 16'b0000000000000000;
	sram_mem[96788] = 16'b0000000000000000;
	sram_mem[96789] = 16'b0000000000000000;
	sram_mem[96790] = 16'b0000000000000000;
	sram_mem[96791] = 16'b0000000000000000;
	sram_mem[96792] = 16'b0000000000000000;
	sram_mem[96793] = 16'b0000000000000000;
	sram_mem[96794] = 16'b0000000000000000;
	sram_mem[96795] = 16'b0000000000000000;
	sram_mem[96796] = 16'b0000000000000000;
	sram_mem[96797] = 16'b0000000000000000;
	sram_mem[96798] = 16'b0000000000000000;
	sram_mem[96799] = 16'b0000000000000000;
	sram_mem[96800] = 16'b0000000000000000;
	sram_mem[96801] = 16'b0000000000000000;
	sram_mem[96802] = 16'b0000000000000000;
	sram_mem[96803] = 16'b0000000000000000;
	sram_mem[96804] = 16'b0000000000000000;
	sram_mem[96805] = 16'b0000000000000000;
	sram_mem[96806] = 16'b0000000000000000;
	sram_mem[96807] = 16'b0000000000000000;
	sram_mem[96808] = 16'b0000000000000000;
	sram_mem[96809] = 16'b0000000000000000;
	sram_mem[96810] = 16'b0000000000000000;
	sram_mem[96811] = 16'b0000000000000000;
	sram_mem[96812] = 16'b0000000000000000;
	sram_mem[96813] = 16'b0000000000000000;
	sram_mem[96814] = 16'b0000000000000000;
	sram_mem[96815] = 16'b0000000000000000;
	sram_mem[96816] = 16'b0000000000000000;
	sram_mem[96817] = 16'b0000000000000000;
	sram_mem[96818] = 16'b0000000000000000;
	sram_mem[96819] = 16'b0000000000000000;
	sram_mem[96820] = 16'b0000000000000000;
	sram_mem[96821] = 16'b0000000000000000;
	sram_mem[96822] = 16'b0000000000000000;
	sram_mem[96823] = 16'b0000000000000000;
	sram_mem[96824] = 16'b0000000000000000;
	sram_mem[96825] = 16'b0000000000000000;
	sram_mem[96826] = 16'b0000000000000000;
	sram_mem[96827] = 16'b0000000000000000;
	sram_mem[96828] = 16'b0000000000000000;
	sram_mem[96829] = 16'b0000000000000000;
	sram_mem[96830] = 16'b0000000000000000;
	sram_mem[96831] = 16'b0000000000000000;
	sram_mem[96832] = 16'b0000000000000000;
	sram_mem[96833] = 16'b0000000000000000;
	sram_mem[96834] = 16'b0000000000000000;
	sram_mem[96835] = 16'b0000000000000000;
	sram_mem[96836] = 16'b0000000000000000;
	sram_mem[96837] = 16'b0000000000000000;
	sram_mem[96838] = 16'b0000000000000000;
	sram_mem[96839] = 16'b0000000000000000;
	sram_mem[96840] = 16'b0000000000000000;
	sram_mem[96841] = 16'b0000000000000000;
	sram_mem[96842] = 16'b0000000000000000;
	sram_mem[96843] = 16'b0000000000000000;
	sram_mem[96844] = 16'b0000000000000000;
	sram_mem[96845] = 16'b0000000000000000;
	sram_mem[96846] = 16'b0000000000000000;
	sram_mem[96847] = 16'b0000000000000000;
	sram_mem[96848] = 16'b0000000000000000;
	sram_mem[96849] = 16'b0000000000000000;
	sram_mem[96850] = 16'b0000000000000000;
	sram_mem[96851] = 16'b0000000000000000;
	sram_mem[96852] = 16'b0000000000000000;
	sram_mem[96853] = 16'b0000000000000000;
	sram_mem[96854] = 16'b0000000000000000;
	sram_mem[96855] = 16'b0000000000000000;
	sram_mem[96856] = 16'b0000000000000000;
	sram_mem[96857] = 16'b0000000000000000;
	sram_mem[96858] = 16'b0000000000000000;
	sram_mem[96859] = 16'b0000000000000000;
	sram_mem[96860] = 16'b0000000000000000;
	sram_mem[96861] = 16'b0000000000000000;
	sram_mem[96862] = 16'b0000000000000000;
	sram_mem[96863] = 16'b0000000000000000;
	sram_mem[96864] = 16'b0000000000000000;
	sram_mem[96865] = 16'b0000000000000000;
	sram_mem[96866] = 16'b0000000000000000;
	sram_mem[96867] = 16'b0000000000000000;
	sram_mem[96868] = 16'b0000000000000000;
	sram_mem[96869] = 16'b0000000000000000;
	sram_mem[96870] = 16'b0000000000000000;
	sram_mem[96871] = 16'b0000000000000000;
	sram_mem[96872] = 16'b0000000000000000;
	sram_mem[96873] = 16'b0000000000000000;
	sram_mem[96874] = 16'b0000000000000000;
	sram_mem[96875] = 16'b0000000000000000;
	sram_mem[96876] = 16'b0000000000000000;
	sram_mem[96877] = 16'b0000000000000000;
	sram_mem[96878] = 16'b0000000000000000;
	sram_mem[96879] = 16'b0000000000000000;
	sram_mem[96880] = 16'b0000000000000000;
	sram_mem[96881] = 16'b0000000000000000;
	sram_mem[96882] = 16'b0000000000000000;
	sram_mem[96883] = 16'b0000000000000000;
	sram_mem[96884] = 16'b0000000000000000;
	sram_mem[96885] = 16'b0000000000000000;
	sram_mem[96886] = 16'b0000000000000000;
	sram_mem[96887] = 16'b0000000000000000;
	sram_mem[96888] = 16'b0000000000000000;
	sram_mem[96889] = 16'b0000000000000000;
	sram_mem[96890] = 16'b0000000000000000;
	sram_mem[96891] = 16'b0000000000000000;
	sram_mem[96892] = 16'b0000000000000000;
	sram_mem[96893] = 16'b0000000000000000;
	sram_mem[96894] = 16'b0000000000000000;
	sram_mem[96895] = 16'b0000000000000000;
	sram_mem[96896] = 16'b0000000000000000;
	sram_mem[96897] = 16'b0000000000000000;
	sram_mem[96898] = 16'b0000000000000000;
	sram_mem[96899] = 16'b0000000000000000;
	sram_mem[96900] = 16'b0000000000000000;
	sram_mem[96901] = 16'b0000000000000000;
	sram_mem[96902] = 16'b0000000000000000;
	sram_mem[96903] = 16'b0000000000000000;
	sram_mem[96904] = 16'b0000000000000000;
	sram_mem[96905] = 16'b0000000000000000;
	sram_mem[96906] = 16'b0000000000000000;
	sram_mem[96907] = 16'b0000000000000000;
	sram_mem[96908] = 16'b0000000000000000;
	sram_mem[96909] = 16'b0000000000000000;
	sram_mem[96910] = 16'b0000000000000000;
	sram_mem[96911] = 16'b0000000000000000;
	sram_mem[96912] = 16'b0000000000000000;
	sram_mem[96913] = 16'b0000000000000000;
	sram_mem[96914] = 16'b0000000000000000;
	sram_mem[96915] = 16'b0000000000000000;
	sram_mem[96916] = 16'b0000000000000000;
	sram_mem[96917] = 16'b0000000000000000;
	sram_mem[96918] = 16'b0000000000000000;
	sram_mem[96919] = 16'b0000000000000000;
	sram_mem[96920] = 16'b0000000000000000;
	sram_mem[96921] = 16'b0000000000000000;
	sram_mem[96922] = 16'b0000000000000000;
	sram_mem[96923] = 16'b0000000000000000;
	sram_mem[96924] = 16'b0000000000000000;
	sram_mem[96925] = 16'b0000000000000000;
	sram_mem[96926] = 16'b0000000000000000;
	sram_mem[96927] = 16'b0000000000000000;
	sram_mem[96928] = 16'b0000000000000000;
	sram_mem[96929] = 16'b0000000000000000;
	sram_mem[96930] = 16'b0000000000000000;
	sram_mem[96931] = 16'b0000000000000000;
	sram_mem[96932] = 16'b0000000000000000;
	sram_mem[96933] = 16'b0000000000000000;
	sram_mem[96934] = 16'b0000000000000000;
	sram_mem[96935] = 16'b0000000000000000;
	sram_mem[96936] = 16'b0000000000000000;
	sram_mem[96937] = 16'b0000000000000000;
	sram_mem[96938] = 16'b0000000000000000;
	sram_mem[96939] = 16'b0000000000000000;
	sram_mem[96940] = 16'b0000000000000000;
	sram_mem[96941] = 16'b0000000000000000;
	sram_mem[96942] = 16'b0000000000000000;
	sram_mem[96943] = 16'b0000000000000000;
	sram_mem[96944] = 16'b0000000000000000;
	sram_mem[96945] = 16'b0000000000000000;
	sram_mem[96946] = 16'b0000000000000000;
	sram_mem[96947] = 16'b0000000000000000;
	sram_mem[96948] = 16'b0000000000000000;
	sram_mem[96949] = 16'b0000000000000000;
	sram_mem[96950] = 16'b0000000000000000;
	sram_mem[96951] = 16'b0000000000000000;
	sram_mem[96952] = 16'b0000000000000000;
	sram_mem[96953] = 16'b0000000000000000;
	sram_mem[96954] = 16'b0000000000000000;
	sram_mem[96955] = 16'b0000000000000000;
	sram_mem[96956] = 16'b0000000000000000;
	sram_mem[96957] = 16'b0000000000000000;
	sram_mem[96958] = 16'b0000000000000000;
	sram_mem[96959] = 16'b0000000000000000;
	sram_mem[96960] = 16'b0000000000000000;
	sram_mem[96961] = 16'b0000000000000000;
	sram_mem[96962] = 16'b0000000000000000;
	sram_mem[96963] = 16'b0000000000000000;
	sram_mem[96964] = 16'b0000000000000000;
	sram_mem[96965] = 16'b0000000000000000;
	sram_mem[96966] = 16'b0000000000000000;
	sram_mem[96967] = 16'b0000000000000000;
	sram_mem[96968] = 16'b0000000000000000;
	sram_mem[96969] = 16'b0000000000000000;
	sram_mem[96970] = 16'b0000000000000000;
	sram_mem[96971] = 16'b0000000000000000;
	sram_mem[96972] = 16'b0000000000000000;
	sram_mem[96973] = 16'b0000000000000000;
	sram_mem[96974] = 16'b0000000000000000;
	sram_mem[96975] = 16'b0000000000000000;
	sram_mem[96976] = 16'b0000000000000000;
	sram_mem[96977] = 16'b0000000000000000;
	sram_mem[96978] = 16'b0000000000000000;
	sram_mem[96979] = 16'b0000000000000000;
	sram_mem[96980] = 16'b0000000000000000;
	sram_mem[96981] = 16'b0000000000000000;
	sram_mem[96982] = 16'b0000000000000000;
	sram_mem[96983] = 16'b0000000000000000;
	sram_mem[96984] = 16'b0000000000000000;
	sram_mem[96985] = 16'b0000000000000000;
	sram_mem[96986] = 16'b0000000000000000;
	sram_mem[96987] = 16'b0000000000000000;
	sram_mem[96988] = 16'b0000000000000000;
	sram_mem[96989] = 16'b0000000000000000;
	sram_mem[96990] = 16'b0000000000000000;
	sram_mem[96991] = 16'b0000000000000000;
	sram_mem[96992] = 16'b0000000000000000;
	sram_mem[96993] = 16'b0000000000000000;
	sram_mem[96994] = 16'b0000000000000000;
	sram_mem[96995] = 16'b0000000000000000;
	sram_mem[96996] = 16'b0000000000000000;
	sram_mem[96997] = 16'b0000000000000000;
	sram_mem[96998] = 16'b0000000000000000;
	sram_mem[96999] = 16'b0000000000000000;
	sram_mem[97000] = 16'b0000000000000000;
	sram_mem[97001] = 16'b0000000000000000;
	sram_mem[97002] = 16'b0000000000000000;
	sram_mem[97003] = 16'b0000000000000000;
	sram_mem[97004] = 16'b0000000000000000;
	sram_mem[97005] = 16'b0000000000000000;
	sram_mem[97006] = 16'b0000000000000000;
	sram_mem[97007] = 16'b0000000000000000;
	sram_mem[97008] = 16'b0000000000000000;
	sram_mem[97009] = 16'b0000000000000000;
	sram_mem[97010] = 16'b0000000000000000;
	sram_mem[97011] = 16'b0000000000000000;
	sram_mem[97012] = 16'b0000000000000000;
	sram_mem[97013] = 16'b0000000000000000;
	sram_mem[97014] = 16'b0000000000000000;
	sram_mem[97015] = 16'b0000000000000000;
	sram_mem[97016] = 16'b0000000000000000;
	sram_mem[97017] = 16'b0000000000000000;
	sram_mem[97018] = 16'b0000000000000000;
	sram_mem[97019] = 16'b0000000000000000;
	sram_mem[97020] = 16'b0000000000000000;
	sram_mem[97021] = 16'b0000000000000000;
	sram_mem[97022] = 16'b0000000000000000;
	sram_mem[97023] = 16'b0000000000000000;
	sram_mem[97024] = 16'b0000000000000000;
	sram_mem[97025] = 16'b0000000000000000;
	sram_mem[97026] = 16'b0000000000000000;
	sram_mem[97027] = 16'b0000000000000000;
	sram_mem[97028] = 16'b0000000000000000;
	sram_mem[97029] = 16'b0000000000000000;
	sram_mem[97030] = 16'b0000000000000000;
	sram_mem[97031] = 16'b0000000000000000;
	sram_mem[97032] = 16'b0000000000000000;
	sram_mem[97033] = 16'b0000000000000000;
	sram_mem[97034] = 16'b0000000000000000;
	sram_mem[97035] = 16'b0000000000000000;
	sram_mem[97036] = 16'b0000000000000000;
	sram_mem[97037] = 16'b0000000000000000;
	sram_mem[97038] = 16'b0000000000000000;
	sram_mem[97039] = 16'b0000000000000000;
	sram_mem[97040] = 16'b0000000000000000;
	sram_mem[97041] = 16'b0000000000000000;
	sram_mem[97042] = 16'b0000000000000000;
	sram_mem[97043] = 16'b0000000000000000;
	sram_mem[97044] = 16'b0000000000000000;
	sram_mem[97045] = 16'b0000000000000000;
	sram_mem[97046] = 16'b0000000000000000;
	sram_mem[97047] = 16'b0000000000000000;
	sram_mem[97048] = 16'b0000000000000000;
	sram_mem[97049] = 16'b0000000000000000;
	sram_mem[97050] = 16'b0000000000000000;
	sram_mem[97051] = 16'b0000000000000000;
	sram_mem[97052] = 16'b0000000000000000;
	sram_mem[97053] = 16'b0000000000000000;
	sram_mem[97054] = 16'b0000000000000000;
	sram_mem[97055] = 16'b0000000000000000;
	sram_mem[97056] = 16'b0000000000000000;
	sram_mem[97057] = 16'b0000000000000000;
	sram_mem[97058] = 16'b0000000000000000;
	sram_mem[97059] = 16'b0000000000000000;
	sram_mem[97060] = 16'b0000000000000000;
	sram_mem[97061] = 16'b0000000000000000;
	sram_mem[97062] = 16'b0000000000000000;
	sram_mem[97063] = 16'b0000000000000000;
	sram_mem[97064] = 16'b0000000000000000;
	sram_mem[97065] = 16'b0000000000000000;
	sram_mem[97066] = 16'b0000000000000000;
	sram_mem[97067] = 16'b0000000000000000;
	sram_mem[97068] = 16'b0000000000000000;
	sram_mem[97069] = 16'b0000000000000000;
	sram_mem[97070] = 16'b0000000000000000;
	sram_mem[97071] = 16'b0000000000000000;
	sram_mem[97072] = 16'b0000000000000000;
	sram_mem[97073] = 16'b0000000000000000;
	sram_mem[97074] = 16'b0000000000000000;
	sram_mem[97075] = 16'b0000000000000000;
	sram_mem[97076] = 16'b0000000000000000;
	sram_mem[97077] = 16'b0000000000000000;
	sram_mem[97078] = 16'b0000000000000000;
	sram_mem[97079] = 16'b0000000000000000;
	sram_mem[97080] = 16'b0000000000000000;
	sram_mem[97081] = 16'b0000000000000000;
	sram_mem[97082] = 16'b0000000000000000;
	sram_mem[97083] = 16'b0000000000000000;
	sram_mem[97084] = 16'b0000000000000000;
	sram_mem[97085] = 16'b0000000000000000;
	sram_mem[97086] = 16'b0000000000000000;
	sram_mem[97087] = 16'b0000000000000000;
	sram_mem[97088] = 16'b0000000000000000;
	sram_mem[97089] = 16'b0000000000000000;
	sram_mem[97090] = 16'b0000000000000000;
	sram_mem[97091] = 16'b0000000000000000;
	sram_mem[97092] = 16'b0000000000000000;
	sram_mem[97093] = 16'b0000000000000000;
	sram_mem[97094] = 16'b0000000000000000;
	sram_mem[97095] = 16'b0000000000000000;
	sram_mem[97096] = 16'b0000000000000000;
	sram_mem[97097] = 16'b0000000000000000;
	sram_mem[97098] = 16'b0000000000000000;
	sram_mem[97099] = 16'b0000000000000000;
	sram_mem[97100] = 16'b0000000000000000;
	sram_mem[97101] = 16'b0000000000000000;
	sram_mem[97102] = 16'b0000000000000000;
	sram_mem[97103] = 16'b0000000000000000;
	sram_mem[97104] = 16'b0000000000000000;
	sram_mem[97105] = 16'b0000000000000000;
	sram_mem[97106] = 16'b0000000000000000;
	sram_mem[97107] = 16'b0000000000000000;
	sram_mem[97108] = 16'b0000000000000000;
	sram_mem[97109] = 16'b0000000000000000;
	sram_mem[97110] = 16'b0000000000000000;
	sram_mem[97111] = 16'b0000000000000000;
	sram_mem[97112] = 16'b0000000000000000;
	sram_mem[97113] = 16'b0000000000000000;
	sram_mem[97114] = 16'b0000000000000000;
	sram_mem[97115] = 16'b0000000000000000;
	sram_mem[97116] = 16'b0000000000000000;
	sram_mem[97117] = 16'b0000000000000000;
	sram_mem[97118] = 16'b0000000000000000;
	sram_mem[97119] = 16'b0000000000000000;
	sram_mem[97120] = 16'b0000000000000000;
	sram_mem[97121] = 16'b0000000000000000;
	sram_mem[97122] = 16'b0000000000000000;
	sram_mem[97123] = 16'b0000000000000000;
	sram_mem[97124] = 16'b0000000000000000;
	sram_mem[97125] = 16'b0000000000000000;
	sram_mem[97126] = 16'b0000000000000000;
	sram_mem[97127] = 16'b0000000000000000;
	sram_mem[97128] = 16'b0000000000000000;
	sram_mem[97129] = 16'b0000000000000000;
	sram_mem[97130] = 16'b0000000000000000;
	sram_mem[97131] = 16'b0000000000000000;
	sram_mem[97132] = 16'b0000000000000000;
	sram_mem[97133] = 16'b0000000000000000;
	sram_mem[97134] = 16'b0000000000000000;
	sram_mem[97135] = 16'b0000000000000000;
	sram_mem[97136] = 16'b0000000000000000;
	sram_mem[97137] = 16'b0000000000000000;
	sram_mem[97138] = 16'b0000000000000000;
	sram_mem[97139] = 16'b0000000000000000;
	sram_mem[97140] = 16'b0000000000000000;
	sram_mem[97141] = 16'b0000000000000000;
	sram_mem[97142] = 16'b0000000000000000;
	sram_mem[97143] = 16'b0000000000000000;
	sram_mem[97144] = 16'b0000000000000000;
	sram_mem[97145] = 16'b0000000000000000;
	sram_mem[97146] = 16'b0000000000000000;
	sram_mem[97147] = 16'b0000000000000000;
	sram_mem[97148] = 16'b0000000000000000;
	sram_mem[97149] = 16'b0000000000000000;
	sram_mem[97150] = 16'b0000000000000000;
	sram_mem[97151] = 16'b0000000000000000;
	sram_mem[97152] = 16'b0000000000000000;
	sram_mem[97153] = 16'b0000000000000000;
	sram_mem[97154] = 16'b0000000000000000;
	sram_mem[97155] = 16'b0000000000000000;
	sram_mem[97156] = 16'b0000000000000000;
	sram_mem[97157] = 16'b0000000000000000;
	sram_mem[97158] = 16'b0000000000000000;
	sram_mem[97159] = 16'b0000000000000000;
	sram_mem[97160] = 16'b0000000000000000;
	sram_mem[97161] = 16'b0000000000000000;
	sram_mem[97162] = 16'b0000000000000000;
	sram_mem[97163] = 16'b0000000000000000;
	sram_mem[97164] = 16'b0000000000000000;
	sram_mem[97165] = 16'b0000000000000000;
	sram_mem[97166] = 16'b0000000000000000;
	sram_mem[97167] = 16'b0000000000000000;
	sram_mem[97168] = 16'b0000000000000000;
	sram_mem[97169] = 16'b0000000000000000;
	sram_mem[97170] = 16'b0000000000000000;
	sram_mem[97171] = 16'b0000000000000000;
	sram_mem[97172] = 16'b0000000000000000;
	sram_mem[97173] = 16'b0000000000000000;
	sram_mem[97174] = 16'b0000000000000000;
	sram_mem[97175] = 16'b0000000000000000;
	sram_mem[97176] = 16'b0000000000000000;
	sram_mem[97177] = 16'b0000000000000000;
	sram_mem[97178] = 16'b0000000000000000;
	sram_mem[97179] = 16'b0000000000000000;
	sram_mem[97180] = 16'b0000000000000000;
	sram_mem[97181] = 16'b0000000000000000;
	sram_mem[97182] = 16'b0000000000000000;
	sram_mem[97183] = 16'b0000000000000000;
	sram_mem[97184] = 16'b0000000000000000;
	sram_mem[97185] = 16'b0000000000000000;
	sram_mem[97186] = 16'b0000000000000000;
	sram_mem[97187] = 16'b0000000000000000;
	sram_mem[97188] = 16'b0000000000000000;
	sram_mem[97189] = 16'b0000000000000000;
	sram_mem[97190] = 16'b0000000000000000;
	sram_mem[97191] = 16'b0000000000000000;
	sram_mem[97192] = 16'b0000000000000000;
	sram_mem[97193] = 16'b0000000000000000;
	sram_mem[97194] = 16'b0000000000000000;
	sram_mem[97195] = 16'b0000000000000000;
	sram_mem[97196] = 16'b0000000000000000;
	sram_mem[97197] = 16'b0000000000000000;
	sram_mem[97198] = 16'b0000000000000000;
	sram_mem[97199] = 16'b0000000000000000;
	sram_mem[97200] = 16'b0000000000000000;
	sram_mem[97201] = 16'b0000000000000000;
	sram_mem[97202] = 16'b0000000000000000;
	sram_mem[97203] = 16'b0000000000000000;
	sram_mem[97204] = 16'b0000000000000000;
	sram_mem[97205] = 16'b0000000000000000;
	sram_mem[97206] = 16'b0000000000000000;
	sram_mem[97207] = 16'b0000000000000000;
	sram_mem[97208] = 16'b0000000000000000;
	sram_mem[97209] = 16'b0000000000000000;
	sram_mem[97210] = 16'b0000000000000000;
	sram_mem[97211] = 16'b0000000000000000;
	sram_mem[97212] = 16'b0000000000000000;
	sram_mem[97213] = 16'b0000000000000000;
	sram_mem[97214] = 16'b0000000000000000;
	sram_mem[97215] = 16'b0000000000000000;
	sram_mem[97216] = 16'b0000000000000000;
	sram_mem[97217] = 16'b0000000000000000;
	sram_mem[97218] = 16'b0000000000000000;
	sram_mem[97219] = 16'b0000000000000000;
	sram_mem[97220] = 16'b0000000000000000;
	sram_mem[97221] = 16'b0000000000000000;
	sram_mem[97222] = 16'b0000000000000000;
	sram_mem[97223] = 16'b0000000000000000;
	sram_mem[97224] = 16'b0000000000000000;
	sram_mem[97225] = 16'b0000000000000000;
	sram_mem[97226] = 16'b0000000000000000;
	sram_mem[97227] = 16'b0000000000000000;
	sram_mem[97228] = 16'b0000000000000000;
	sram_mem[97229] = 16'b0000000000000000;
	sram_mem[97230] = 16'b0000000000000000;
	sram_mem[97231] = 16'b0000000000000000;
	sram_mem[97232] = 16'b0000000000000000;
	sram_mem[97233] = 16'b0000000000000000;
	sram_mem[97234] = 16'b0000000000000000;
	sram_mem[97235] = 16'b0000000000000000;
	sram_mem[97236] = 16'b0000000000000000;
	sram_mem[97237] = 16'b0000000000000000;
	sram_mem[97238] = 16'b0000000000000000;
	sram_mem[97239] = 16'b0000000000000000;
	sram_mem[97240] = 16'b0000000000000000;
	sram_mem[97241] = 16'b0000000000000000;
	sram_mem[97242] = 16'b0000000000000000;
	sram_mem[97243] = 16'b0000000000000000;
	sram_mem[97244] = 16'b0000000000000000;
	sram_mem[97245] = 16'b0000000000000000;
	sram_mem[97246] = 16'b0000000000000000;
	sram_mem[97247] = 16'b0000000000000000;
	sram_mem[97248] = 16'b0000000000000000;
	sram_mem[97249] = 16'b0000000000000000;
	sram_mem[97250] = 16'b0000000000000000;
	sram_mem[97251] = 16'b0000000000000000;
	sram_mem[97252] = 16'b0000000000000000;
	sram_mem[97253] = 16'b0000000000000000;
	sram_mem[97254] = 16'b0000000000000000;
	sram_mem[97255] = 16'b0000000000000000;
	sram_mem[97256] = 16'b0000000000000000;
	sram_mem[97257] = 16'b0000000000000000;
	sram_mem[97258] = 16'b0000000000000000;
	sram_mem[97259] = 16'b0000000000000000;
	sram_mem[97260] = 16'b0000000000000000;
	sram_mem[97261] = 16'b0000000000000000;
	sram_mem[97262] = 16'b0000000000000000;
	sram_mem[97263] = 16'b0000000000000000;
	sram_mem[97264] = 16'b0000000000000000;
	sram_mem[97265] = 16'b0000000000000000;
	sram_mem[97266] = 16'b0000000000000000;
	sram_mem[97267] = 16'b0000000000000000;
	sram_mem[97268] = 16'b0000000000000000;
	sram_mem[97269] = 16'b0000000000000000;
	sram_mem[97270] = 16'b0000000000000000;
	sram_mem[97271] = 16'b0000000000000000;
	sram_mem[97272] = 16'b0000000000000000;
	sram_mem[97273] = 16'b0000000000000000;
	sram_mem[97274] = 16'b0000000000000000;
	sram_mem[97275] = 16'b0000000000000000;
	sram_mem[97276] = 16'b0000000000000000;
	sram_mem[97277] = 16'b0000000000000000;
	sram_mem[97278] = 16'b0000000000000000;
	sram_mem[97279] = 16'b0000000000000000;
	sram_mem[97280] = 16'b0000000000000000;
	sram_mem[97281] = 16'b0000000000000000;
	sram_mem[97282] = 16'b0000000000000000;
	sram_mem[97283] = 16'b0000000000000000;
	sram_mem[97284] = 16'b0000000000000000;
	sram_mem[97285] = 16'b0000000000000000;
	sram_mem[97286] = 16'b0000000000000000;
	sram_mem[97287] = 16'b0000000000000000;
	sram_mem[97288] = 16'b0000000000000000;
	sram_mem[97289] = 16'b0000000000000000;
	sram_mem[97290] = 16'b0000000000000000;
	sram_mem[97291] = 16'b0000000000000000;
	sram_mem[97292] = 16'b0000000000000000;
	sram_mem[97293] = 16'b0000000000000000;
	sram_mem[97294] = 16'b0000000000000000;
	sram_mem[97295] = 16'b0000000000000000;
	sram_mem[97296] = 16'b0000000000000000;
	sram_mem[97297] = 16'b0000000000000000;
	sram_mem[97298] = 16'b0000000000000000;
	sram_mem[97299] = 16'b0000000000000000;
	sram_mem[97300] = 16'b0000000000000000;
	sram_mem[97301] = 16'b0000000000000000;
	sram_mem[97302] = 16'b0000000000000000;
	sram_mem[97303] = 16'b0000000000000000;
	sram_mem[97304] = 16'b0000000000000000;
	sram_mem[97305] = 16'b0000000000000000;
	sram_mem[97306] = 16'b0000000000000000;
	sram_mem[97307] = 16'b0000000000000000;
	sram_mem[97308] = 16'b0000000000000000;
	sram_mem[97309] = 16'b0000000000000000;
	sram_mem[97310] = 16'b0000000000000000;
	sram_mem[97311] = 16'b0000000000000000;
	sram_mem[97312] = 16'b0000000000000000;
	sram_mem[97313] = 16'b0000000000000000;
	sram_mem[97314] = 16'b0000000000000000;
	sram_mem[97315] = 16'b0000000000000000;
	sram_mem[97316] = 16'b0000000000000000;
	sram_mem[97317] = 16'b0000000000000000;
	sram_mem[97318] = 16'b0000000000000000;
	sram_mem[97319] = 16'b0000000000000000;
	sram_mem[97320] = 16'b0000000000000000;
	sram_mem[97321] = 16'b0000000000000000;
	sram_mem[97322] = 16'b0000000000000000;
	sram_mem[97323] = 16'b0000000000000000;
	sram_mem[97324] = 16'b0000000000000000;
	sram_mem[97325] = 16'b0000000000000000;
	sram_mem[97326] = 16'b0000000000000000;
	sram_mem[97327] = 16'b0000000000000000;
	sram_mem[97328] = 16'b0000000000000000;
	sram_mem[97329] = 16'b0000000000000000;
	sram_mem[97330] = 16'b0000000000000000;
	sram_mem[97331] = 16'b0000000000000000;
	sram_mem[97332] = 16'b0000000000000000;
	sram_mem[97333] = 16'b0000000000000000;
	sram_mem[97334] = 16'b0000000000000000;
	sram_mem[97335] = 16'b0000000000000000;
	sram_mem[97336] = 16'b0000000000000000;
	sram_mem[97337] = 16'b0000000000000000;
	sram_mem[97338] = 16'b0000000000000000;
	sram_mem[97339] = 16'b0000000000000000;
	sram_mem[97340] = 16'b0000000000000000;
	sram_mem[97341] = 16'b0000000000000000;
	sram_mem[97342] = 16'b0000000000000000;
	sram_mem[97343] = 16'b0000000000000000;
	sram_mem[97344] = 16'b0000000000000000;
	sram_mem[97345] = 16'b0000000000000000;
	sram_mem[97346] = 16'b0000000000000000;
	sram_mem[97347] = 16'b0000000000000000;
	sram_mem[97348] = 16'b0000000000000000;
	sram_mem[97349] = 16'b0000000000000000;
	sram_mem[97350] = 16'b0000000000000000;
	sram_mem[97351] = 16'b0000000000000000;
	sram_mem[97352] = 16'b0000000000000000;
	sram_mem[97353] = 16'b0000000000000000;
	sram_mem[97354] = 16'b0000000000000000;
	sram_mem[97355] = 16'b0000000000000000;
	sram_mem[97356] = 16'b0000000000000000;
	sram_mem[97357] = 16'b0000000000000000;
	sram_mem[97358] = 16'b0000000000000000;
	sram_mem[97359] = 16'b0000000000000000;
	sram_mem[97360] = 16'b0000000000000000;
	sram_mem[97361] = 16'b0000000000000000;
	sram_mem[97362] = 16'b0000000000000000;
	sram_mem[97363] = 16'b0000000000000000;
	sram_mem[97364] = 16'b0000000000000000;
	sram_mem[97365] = 16'b0000000000000000;
	sram_mem[97366] = 16'b0000000000000000;
	sram_mem[97367] = 16'b0000000000000000;
	sram_mem[97368] = 16'b0000000000000000;
	sram_mem[97369] = 16'b0000000000000000;
	sram_mem[97370] = 16'b0000000000000000;
	sram_mem[97371] = 16'b0000000000000000;
	sram_mem[97372] = 16'b0000000000000000;
	sram_mem[97373] = 16'b0000000000000000;
	sram_mem[97374] = 16'b0000000000000000;
	sram_mem[97375] = 16'b0000000000000000;
	sram_mem[97376] = 16'b0000000000000000;
	sram_mem[97377] = 16'b0000000000000000;
	sram_mem[97378] = 16'b0000000000000000;
	sram_mem[97379] = 16'b0000000000000000;
	sram_mem[97380] = 16'b0000000000000000;
	sram_mem[97381] = 16'b0000000000000000;
	sram_mem[97382] = 16'b0000000000000000;
	sram_mem[97383] = 16'b0000000000000000;
	sram_mem[97384] = 16'b0000000000000000;
	sram_mem[97385] = 16'b0000000000000000;
	sram_mem[97386] = 16'b0000000000000000;
	sram_mem[97387] = 16'b0000000000000000;
	sram_mem[97388] = 16'b0000000000000000;
	sram_mem[97389] = 16'b0000000000000000;
	sram_mem[97390] = 16'b0000000000000000;
	sram_mem[97391] = 16'b0000000000000000;
	sram_mem[97392] = 16'b0000000000000000;
	sram_mem[97393] = 16'b0000000000000000;
	sram_mem[97394] = 16'b0000000000000000;
	sram_mem[97395] = 16'b0000000000000000;
	sram_mem[97396] = 16'b0000000000000000;
	sram_mem[97397] = 16'b0000000000000000;
	sram_mem[97398] = 16'b0000000000000000;
	sram_mem[97399] = 16'b0000000000000000;
	sram_mem[97400] = 16'b0000000000000000;
	sram_mem[97401] = 16'b0000000000000000;
	sram_mem[97402] = 16'b0000000000000000;
	sram_mem[97403] = 16'b0000000000000000;
	sram_mem[97404] = 16'b0000000000000000;
	sram_mem[97405] = 16'b0000000000000000;
	sram_mem[97406] = 16'b0000000000000000;
	sram_mem[97407] = 16'b0000000000000000;
	sram_mem[97408] = 16'b0000000000000000;
	sram_mem[97409] = 16'b0000000000000000;
	sram_mem[97410] = 16'b0000000000000000;
	sram_mem[97411] = 16'b0000000000000000;
	sram_mem[97412] = 16'b0000000000000000;
	sram_mem[97413] = 16'b0000000000000000;
	sram_mem[97414] = 16'b0000000000000000;
	sram_mem[97415] = 16'b0000000000000000;
	sram_mem[97416] = 16'b0000000000000000;
	sram_mem[97417] = 16'b0000000000000000;
	sram_mem[97418] = 16'b0000000000000000;
	sram_mem[97419] = 16'b0000000000000000;
	sram_mem[97420] = 16'b0000000000000000;
	sram_mem[97421] = 16'b0000000000000000;
	sram_mem[97422] = 16'b0000000000000000;
	sram_mem[97423] = 16'b0000000000000000;
	sram_mem[97424] = 16'b0000000000000000;
	sram_mem[97425] = 16'b0000000000000000;
	sram_mem[97426] = 16'b0000000000000000;
	sram_mem[97427] = 16'b0000000000000000;
	sram_mem[97428] = 16'b0000000000000000;
	sram_mem[97429] = 16'b0000000000000000;
	sram_mem[97430] = 16'b0000000000000000;
	sram_mem[97431] = 16'b0000000000000000;
	sram_mem[97432] = 16'b0000000000000000;
	sram_mem[97433] = 16'b0000000000000000;
	sram_mem[97434] = 16'b0000000000000000;
	sram_mem[97435] = 16'b0000000000000000;
	sram_mem[97436] = 16'b0000000000000000;
	sram_mem[97437] = 16'b0000000000000000;
	sram_mem[97438] = 16'b0000000000000000;
	sram_mem[97439] = 16'b0000000000000000;
	sram_mem[97440] = 16'b0000000000000000;
	sram_mem[97441] = 16'b0000000000000000;
	sram_mem[97442] = 16'b0000000000000000;
	sram_mem[97443] = 16'b0000000000000000;
	sram_mem[97444] = 16'b0000000000000000;
	sram_mem[97445] = 16'b0000000000000000;
	sram_mem[97446] = 16'b0000000000000000;
	sram_mem[97447] = 16'b0000000000000000;
	sram_mem[97448] = 16'b0000000000000000;
	sram_mem[97449] = 16'b0000000000000000;
	sram_mem[97450] = 16'b0000000000000000;
	sram_mem[97451] = 16'b0000000000000000;
	sram_mem[97452] = 16'b0000000000000000;
	sram_mem[97453] = 16'b0000000000000000;
	sram_mem[97454] = 16'b0000000000000000;
	sram_mem[97455] = 16'b0000000000000000;
	sram_mem[97456] = 16'b0000000000000000;
	sram_mem[97457] = 16'b0000000000000000;
	sram_mem[97458] = 16'b0000000000000000;
	sram_mem[97459] = 16'b0000000000000000;
	sram_mem[97460] = 16'b0000000000000000;
	sram_mem[97461] = 16'b0000000000000000;
	sram_mem[97462] = 16'b0000000000000000;
	sram_mem[97463] = 16'b0000000000000000;
	sram_mem[97464] = 16'b0000000000000000;
	sram_mem[97465] = 16'b0000000000000000;
	sram_mem[97466] = 16'b0000000000000000;
	sram_mem[97467] = 16'b0000000000000000;
	sram_mem[97468] = 16'b0000000000000000;
	sram_mem[97469] = 16'b0000000000000000;
	sram_mem[97470] = 16'b0000000000000000;
	sram_mem[97471] = 16'b0000000000000000;
	sram_mem[97472] = 16'b0000000000000000;
	sram_mem[97473] = 16'b0000000000000000;
	sram_mem[97474] = 16'b0000000000000000;
	sram_mem[97475] = 16'b0000000000000000;
	sram_mem[97476] = 16'b0000000000000000;
	sram_mem[97477] = 16'b0000000000000000;
	sram_mem[97478] = 16'b0000000000000000;
	sram_mem[97479] = 16'b0000000000000000;
	sram_mem[97480] = 16'b0000000000000000;
	sram_mem[97481] = 16'b0000000000000000;
	sram_mem[97482] = 16'b0000000000000000;
	sram_mem[97483] = 16'b0000000000000000;
	sram_mem[97484] = 16'b0000000000000000;
	sram_mem[97485] = 16'b0000000000000000;
	sram_mem[97486] = 16'b0000000000000000;
	sram_mem[97487] = 16'b0000000000000000;
	sram_mem[97488] = 16'b0000000000000000;
	sram_mem[97489] = 16'b0000000000000000;
	sram_mem[97490] = 16'b0000000000000000;
	sram_mem[97491] = 16'b0000000000000000;
	sram_mem[97492] = 16'b0000000000000000;
	sram_mem[97493] = 16'b0000000000000000;
	sram_mem[97494] = 16'b0000000000000000;
	sram_mem[97495] = 16'b0000000000000000;
	sram_mem[97496] = 16'b0000000000000000;
	sram_mem[97497] = 16'b0000000000000000;
	sram_mem[97498] = 16'b0000000000000000;
	sram_mem[97499] = 16'b0000000000000000;
	sram_mem[97500] = 16'b0000000000000000;
	sram_mem[97501] = 16'b0000000000000000;
	sram_mem[97502] = 16'b0000000000000000;
	sram_mem[97503] = 16'b0000000000000000;
	sram_mem[97504] = 16'b0000000000000000;
	sram_mem[97505] = 16'b0000000000000000;
	sram_mem[97506] = 16'b0000000000000000;
	sram_mem[97507] = 16'b0000000000000000;
	sram_mem[97508] = 16'b0000000000000000;
	sram_mem[97509] = 16'b0000000000000000;
	sram_mem[97510] = 16'b0000000000000000;
	sram_mem[97511] = 16'b0000000000000000;
	sram_mem[97512] = 16'b0000000000000000;
	sram_mem[97513] = 16'b0000000000000000;
	sram_mem[97514] = 16'b0000000000000000;
	sram_mem[97515] = 16'b0000000000000000;
	sram_mem[97516] = 16'b0000000000000000;
	sram_mem[97517] = 16'b0000000000000000;
	sram_mem[97518] = 16'b0000000000000000;
	sram_mem[97519] = 16'b0000000000000000;
	sram_mem[97520] = 16'b0000000000000000;
	sram_mem[97521] = 16'b0000000000000000;
	sram_mem[97522] = 16'b0000000000000000;
	sram_mem[97523] = 16'b0000000000000000;
	sram_mem[97524] = 16'b0000000000000000;
	sram_mem[97525] = 16'b0000000000000000;
	sram_mem[97526] = 16'b0000000000000000;
	sram_mem[97527] = 16'b0000000000000000;
	sram_mem[97528] = 16'b0000000000000000;
	sram_mem[97529] = 16'b0000000000000000;
	sram_mem[97530] = 16'b0000000000000000;
	sram_mem[97531] = 16'b0000000000000000;
	sram_mem[97532] = 16'b0000000000000000;
	sram_mem[97533] = 16'b0000000000000000;
	sram_mem[97534] = 16'b0000000000000000;
	sram_mem[97535] = 16'b0000000000000000;
	sram_mem[97536] = 16'b0000000000000000;
	sram_mem[97537] = 16'b0000000000000000;
	sram_mem[97538] = 16'b0000000000000000;
	sram_mem[97539] = 16'b0000000000000000;
	sram_mem[97540] = 16'b0000000000000000;
	sram_mem[97541] = 16'b0000000000000000;
	sram_mem[97542] = 16'b0000000000000000;
	sram_mem[97543] = 16'b0000000000000000;
	sram_mem[97544] = 16'b0000000000000000;
	sram_mem[97545] = 16'b0000000000000000;
	sram_mem[97546] = 16'b0000000000000000;
	sram_mem[97547] = 16'b0000000000000000;
	sram_mem[97548] = 16'b0000000000000000;
	sram_mem[97549] = 16'b0000000000000000;
	sram_mem[97550] = 16'b0000000000000000;
	sram_mem[97551] = 16'b0000000000000000;
	sram_mem[97552] = 16'b0000000000000000;
	sram_mem[97553] = 16'b0000000000000000;
	sram_mem[97554] = 16'b0000000000000000;
	sram_mem[97555] = 16'b0000000000000000;
	sram_mem[97556] = 16'b0000000000000000;
	sram_mem[97557] = 16'b0000000000000000;
	sram_mem[97558] = 16'b0000000000000000;
	sram_mem[97559] = 16'b0000000000000000;
	sram_mem[97560] = 16'b0000000000000000;
	sram_mem[97561] = 16'b0000000000000000;
	sram_mem[97562] = 16'b0000000000000000;
	sram_mem[97563] = 16'b0000000000000000;
	sram_mem[97564] = 16'b0000000000000000;
	sram_mem[97565] = 16'b0000000000000000;
	sram_mem[97566] = 16'b0000000000000000;
	sram_mem[97567] = 16'b0000000000000000;
	sram_mem[97568] = 16'b0000000000000000;
	sram_mem[97569] = 16'b0000000000000000;
	sram_mem[97570] = 16'b0000000000000000;
	sram_mem[97571] = 16'b0000000000000000;
	sram_mem[97572] = 16'b0000000000000000;
	sram_mem[97573] = 16'b0000000000000000;
	sram_mem[97574] = 16'b0000000000000000;
	sram_mem[97575] = 16'b0000000000000000;
	sram_mem[97576] = 16'b0000000000000000;
	sram_mem[97577] = 16'b0000000000000000;
	sram_mem[97578] = 16'b0000000000000000;
	sram_mem[97579] = 16'b0000000000000000;
	sram_mem[97580] = 16'b0000000000000000;
	sram_mem[97581] = 16'b0000000000000000;
	sram_mem[97582] = 16'b0000000000000000;
	sram_mem[97583] = 16'b0000000000000000;
	sram_mem[97584] = 16'b0000000000000000;
	sram_mem[97585] = 16'b0000000000000000;
	sram_mem[97586] = 16'b0000000000000000;
	sram_mem[97587] = 16'b0000000000000000;
	sram_mem[97588] = 16'b0000000000000000;
	sram_mem[97589] = 16'b0000000000000000;
	sram_mem[97590] = 16'b0000000000000000;
	sram_mem[97591] = 16'b0000000000000000;
	sram_mem[97592] = 16'b0000000000000000;
	sram_mem[97593] = 16'b0000000000000000;
	sram_mem[97594] = 16'b0000000000000000;
	sram_mem[97595] = 16'b0000000000000000;
	sram_mem[97596] = 16'b0000000000000000;
	sram_mem[97597] = 16'b0000000000000000;
	sram_mem[97598] = 16'b0000000000000000;
	sram_mem[97599] = 16'b0000000000000000;
	sram_mem[97600] = 16'b0000000000000000;
	sram_mem[97601] = 16'b0000000000000000;
	sram_mem[97602] = 16'b0000000000000000;
	sram_mem[97603] = 16'b0000000000000000;
	sram_mem[97604] = 16'b0000000000000000;
	sram_mem[97605] = 16'b0000000000000000;
	sram_mem[97606] = 16'b0000000000000000;
	sram_mem[97607] = 16'b0000000000000000;
	sram_mem[97608] = 16'b0000000000000000;
	sram_mem[97609] = 16'b0000000000000000;
	sram_mem[97610] = 16'b0000000000000000;
	sram_mem[97611] = 16'b0000000000000000;
	sram_mem[97612] = 16'b0000000000000000;
	sram_mem[97613] = 16'b0000000000000000;
	sram_mem[97614] = 16'b0000000000000000;
	sram_mem[97615] = 16'b0000000000000000;
	sram_mem[97616] = 16'b0000000000000000;
	sram_mem[97617] = 16'b0000000000000000;
	sram_mem[97618] = 16'b0000000000000000;
	sram_mem[97619] = 16'b0000000000000000;
	sram_mem[97620] = 16'b0000000000000000;
	sram_mem[97621] = 16'b0000000000000000;
	sram_mem[97622] = 16'b0000000000000000;
	sram_mem[97623] = 16'b0000000000000000;
	sram_mem[97624] = 16'b0000000000000000;
	sram_mem[97625] = 16'b0000000000000000;
	sram_mem[97626] = 16'b0000000000000000;
	sram_mem[97627] = 16'b0000000000000000;
	sram_mem[97628] = 16'b0000000000000000;
	sram_mem[97629] = 16'b0000000000000000;
	sram_mem[97630] = 16'b0000000000000000;
	sram_mem[97631] = 16'b0000000000000000;
	sram_mem[97632] = 16'b0000000000000000;
	sram_mem[97633] = 16'b0000000000000000;
	sram_mem[97634] = 16'b0000000000000000;
	sram_mem[97635] = 16'b0000000000000000;
	sram_mem[97636] = 16'b0000000000000000;
	sram_mem[97637] = 16'b0000000000000000;
	sram_mem[97638] = 16'b0000000000000000;
	sram_mem[97639] = 16'b0000000000000000;
	sram_mem[97640] = 16'b0000000000000000;
	sram_mem[97641] = 16'b0000000000000000;
	sram_mem[97642] = 16'b0000000000000000;
	sram_mem[97643] = 16'b0000000000000000;
	sram_mem[97644] = 16'b0000000000000000;
	sram_mem[97645] = 16'b0000000000000000;
	sram_mem[97646] = 16'b0000000000000000;
	sram_mem[97647] = 16'b0000000000000000;
	sram_mem[97648] = 16'b0000000000000000;
	sram_mem[97649] = 16'b0000000000000000;
	sram_mem[97650] = 16'b0000000000000000;
	sram_mem[97651] = 16'b0000000000000000;
	sram_mem[97652] = 16'b0000000000000000;
	sram_mem[97653] = 16'b0000000000000000;
	sram_mem[97654] = 16'b0000000000000000;
	sram_mem[97655] = 16'b0000000000000000;
	sram_mem[97656] = 16'b0000000000000000;
	sram_mem[97657] = 16'b0000000000000000;
	sram_mem[97658] = 16'b0000000000000000;
	sram_mem[97659] = 16'b0000000000000000;
	sram_mem[97660] = 16'b0000000000000000;
	sram_mem[97661] = 16'b0000000000000000;
	sram_mem[97662] = 16'b0000000000000000;
	sram_mem[97663] = 16'b0000000000000000;
	sram_mem[97664] = 16'b0000000000000000;
	sram_mem[97665] = 16'b0000000000000000;
	sram_mem[97666] = 16'b0000000000000000;
	sram_mem[97667] = 16'b0000000000000000;
	sram_mem[97668] = 16'b0000000000000000;
	sram_mem[97669] = 16'b0000000000000000;
	sram_mem[97670] = 16'b0000000000000000;
	sram_mem[97671] = 16'b0000000000000000;
	sram_mem[97672] = 16'b0000000000000000;
	sram_mem[97673] = 16'b0000000000000000;
	sram_mem[97674] = 16'b0000000000000000;
	sram_mem[97675] = 16'b0000000000000000;
	sram_mem[97676] = 16'b0000000000000000;
	sram_mem[97677] = 16'b0000000000000000;
	sram_mem[97678] = 16'b0000000000000000;
	sram_mem[97679] = 16'b0000000000000000;
	sram_mem[97680] = 16'b0000000000000000;
	sram_mem[97681] = 16'b0000000000000000;
	sram_mem[97682] = 16'b0000000000000000;
	sram_mem[97683] = 16'b0000000000000000;
	sram_mem[97684] = 16'b0000000000000000;
	sram_mem[97685] = 16'b0000000000000000;
	sram_mem[97686] = 16'b0000000000000000;
	sram_mem[97687] = 16'b0000000000000000;
	sram_mem[97688] = 16'b0000000000000000;
	sram_mem[97689] = 16'b0000000000000000;
	sram_mem[97690] = 16'b0000000000000000;
	sram_mem[97691] = 16'b0000000000000000;
	sram_mem[97692] = 16'b0000000000000000;
	sram_mem[97693] = 16'b0000000000000000;
	sram_mem[97694] = 16'b0000000000000000;
	sram_mem[97695] = 16'b0000000000000000;
	sram_mem[97696] = 16'b0000000000000000;
	sram_mem[97697] = 16'b0000000000000000;
	sram_mem[97698] = 16'b0000000000000000;
	sram_mem[97699] = 16'b0000000000000000;
	sram_mem[97700] = 16'b0000000000000000;
	sram_mem[97701] = 16'b0000000000000000;
	sram_mem[97702] = 16'b0000000000000000;
	sram_mem[97703] = 16'b0000000000000000;
	sram_mem[97704] = 16'b0000000000000000;
	sram_mem[97705] = 16'b0000000000000000;
	sram_mem[97706] = 16'b0000000000000000;
	sram_mem[97707] = 16'b0000000000000000;
	sram_mem[97708] = 16'b0000000000000000;
	sram_mem[97709] = 16'b0000000000000000;
	sram_mem[97710] = 16'b0000000000000000;
	sram_mem[97711] = 16'b0000000000000000;
	sram_mem[97712] = 16'b0000000000000000;
	sram_mem[97713] = 16'b0000000000000000;
	sram_mem[97714] = 16'b0000000000000000;
	sram_mem[97715] = 16'b0000000000000000;
	sram_mem[97716] = 16'b0000000000000000;
	sram_mem[97717] = 16'b0000000000000000;
	sram_mem[97718] = 16'b0000000000000000;
	sram_mem[97719] = 16'b0000000000000000;
	sram_mem[97720] = 16'b0000000000000000;
	sram_mem[97721] = 16'b0000000000000000;
	sram_mem[97722] = 16'b0000000000000000;
	sram_mem[97723] = 16'b0000000000000000;
	sram_mem[97724] = 16'b0000000000000000;
	sram_mem[97725] = 16'b0000000000000000;
	sram_mem[97726] = 16'b0000000000000000;
	sram_mem[97727] = 16'b0000000000000000;
	sram_mem[97728] = 16'b0000000000000000;
	sram_mem[97729] = 16'b0000000000000000;
	sram_mem[97730] = 16'b0000000000000000;
	sram_mem[97731] = 16'b0000000000000000;
	sram_mem[97732] = 16'b0000000000000000;
	sram_mem[97733] = 16'b0000000000000000;
	sram_mem[97734] = 16'b0000000000000000;
	sram_mem[97735] = 16'b0000000000000000;
	sram_mem[97736] = 16'b0000000000000000;
	sram_mem[97737] = 16'b0000000000000000;
	sram_mem[97738] = 16'b0000000000000000;
	sram_mem[97739] = 16'b0000000000000000;
	sram_mem[97740] = 16'b0000000000000000;
	sram_mem[97741] = 16'b0000000000000000;
	sram_mem[97742] = 16'b0000000000000000;
	sram_mem[97743] = 16'b0000000000000000;
	sram_mem[97744] = 16'b0000000000000000;
	sram_mem[97745] = 16'b0000000000000000;
	sram_mem[97746] = 16'b0000000000000000;
	sram_mem[97747] = 16'b0000000000000000;
	sram_mem[97748] = 16'b0000000000000000;
	sram_mem[97749] = 16'b0000000000000000;
	sram_mem[97750] = 16'b0000000000000000;
	sram_mem[97751] = 16'b0000000000000000;
	sram_mem[97752] = 16'b0000000000000000;
	sram_mem[97753] = 16'b0000000000000000;
	sram_mem[97754] = 16'b0000000000000000;
	sram_mem[97755] = 16'b0000000000000000;
	sram_mem[97756] = 16'b0000000000000000;
	sram_mem[97757] = 16'b0000000000000000;
	sram_mem[97758] = 16'b0000000000000000;
	sram_mem[97759] = 16'b0000000000000000;
	sram_mem[97760] = 16'b0000000000000000;
	sram_mem[97761] = 16'b0000000000000000;
	sram_mem[97762] = 16'b0000000000000000;
	sram_mem[97763] = 16'b0000000000000000;
	sram_mem[97764] = 16'b0000000000000000;
	sram_mem[97765] = 16'b0000000000000000;
	sram_mem[97766] = 16'b0000000000000000;
	sram_mem[97767] = 16'b0000000000000000;
	sram_mem[97768] = 16'b0000000000000000;
	sram_mem[97769] = 16'b0000000000000000;
	sram_mem[97770] = 16'b0000000000000000;
	sram_mem[97771] = 16'b0000000000000000;
	sram_mem[97772] = 16'b0000000000000000;
	sram_mem[97773] = 16'b0000000000000000;
	sram_mem[97774] = 16'b0000000000000000;
	sram_mem[97775] = 16'b0000000000000000;
	sram_mem[97776] = 16'b0000000000000000;
	sram_mem[97777] = 16'b0000000000000000;
	sram_mem[97778] = 16'b0000000000000000;
	sram_mem[97779] = 16'b0000000000000000;
	sram_mem[97780] = 16'b0000000000000000;
	sram_mem[97781] = 16'b0000000000000000;
	sram_mem[97782] = 16'b0000000000000000;
	sram_mem[97783] = 16'b0000000000000000;
	sram_mem[97784] = 16'b0000000000000000;
	sram_mem[97785] = 16'b0000000000000000;
	sram_mem[97786] = 16'b0000000000000000;
	sram_mem[97787] = 16'b0000000000000000;
	sram_mem[97788] = 16'b0000000000000000;
	sram_mem[97789] = 16'b0000000000000000;
	sram_mem[97790] = 16'b0000000000000000;
	sram_mem[97791] = 16'b0000000000000000;
	sram_mem[97792] = 16'b0000000000000000;
	sram_mem[97793] = 16'b0000000000000000;
	sram_mem[97794] = 16'b0000000000000000;
	sram_mem[97795] = 16'b0000000000000000;
	sram_mem[97796] = 16'b0000000000000000;
	sram_mem[97797] = 16'b0000000000000000;
	sram_mem[97798] = 16'b0000000000000000;
	sram_mem[97799] = 16'b0000000000000000;
	sram_mem[97800] = 16'b0000000000000000;
	sram_mem[97801] = 16'b0000000000000000;
	sram_mem[97802] = 16'b0000000000000000;
	sram_mem[97803] = 16'b0000000000000000;
	sram_mem[97804] = 16'b0000000000000000;
	sram_mem[97805] = 16'b0000000000000000;
	sram_mem[97806] = 16'b0000000000000000;
	sram_mem[97807] = 16'b0000000000000000;
	sram_mem[97808] = 16'b0000000000000000;
	sram_mem[97809] = 16'b0000000000000000;
	sram_mem[97810] = 16'b0000000000000000;
	sram_mem[97811] = 16'b0000000000000000;
	sram_mem[97812] = 16'b0000000000000000;
	sram_mem[97813] = 16'b0000000000000000;
	sram_mem[97814] = 16'b0000000000000000;
	sram_mem[97815] = 16'b0000000000000000;
	sram_mem[97816] = 16'b0000000000000000;
	sram_mem[97817] = 16'b0000000000000000;
	sram_mem[97818] = 16'b0000000000000000;
	sram_mem[97819] = 16'b0000000000000000;
	sram_mem[97820] = 16'b0000000000000000;
	sram_mem[97821] = 16'b0000000000000000;
	sram_mem[97822] = 16'b0000000000000000;
	sram_mem[97823] = 16'b0000000000000000;
	sram_mem[97824] = 16'b0000000000000000;
	sram_mem[97825] = 16'b0000000000000000;
	sram_mem[97826] = 16'b0000000000000000;
	sram_mem[97827] = 16'b0000000000000000;
	sram_mem[97828] = 16'b0000000000000000;
	sram_mem[97829] = 16'b0000000000000000;
	sram_mem[97830] = 16'b0000000000000000;
	sram_mem[97831] = 16'b0000000000000000;
	sram_mem[97832] = 16'b0000000000000000;
	sram_mem[97833] = 16'b0000000000000000;
	sram_mem[97834] = 16'b0000000000000000;
	sram_mem[97835] = 16'b0000000000000000;
	sram_mem[97836] = 16'b0000000000000000;
	sram_mem[97837] = 16'b0000000000000000;
	sram_mem[97838] = 16'b0000000000000000;
	sram_mem[97839] = 16'b0000000000000000;
	sram_mem[97840] = 16'b0000000000000000;
	sram_mem[97841] = 16'b0000000000000000;
	sram_mem[97842] = 16'b0000000000000000;
	sram_mem[97843] = 16'b0000000000000000;
	sram_mem[97844] = 16'b0000000000000000;
	sram_mem[97845] = 16'b0000000000000000;
	sram_mem[97846] = 16'b0000000000000000;
	sram_mem[97847] = 16'b0000000000000000;
	sram_mem[97848] = 16'b0000000000000000;
	sram_mem[97849] = 16'b0000000000000000;
	sram_mem[97850] = 16'b0000000000000000;
	sram_mem[97851] = 16'b0000000000000000;
	sram_mem[97852] = 16'b0000000000000000;
	sram_mem[97853] = 16'b0000000000000000;
	sram_mem[97854] = 16'b0000000000000000;
	sram_mem[97855] = 16'b0000000000000000;
	sram_mem[97856] = 16'b0000000000000000;
	sram_mem[97857] = 16'b0000000000000000;
	sram_mem[97858] = 16'b0000000000000000;
	sram_mem[97859] = 16'b0000000000000000;
	sram_mem[97860] = 16'b0000000000000000;
	sram_mem[97861] = 16'b0000000000000000;
	sram_mem[97862] = 16'b0000000000000000;
	sram_mem[97863] = 16'b0000000000000000;
	sram_mem[97864] = 16'b0000000000000000;
	sram_mem[97865] = 16'b0000000000000000;
	sram_mem[97866] = 16'b0000000000000000;
	sram_mem[97867] = 16'b0000000000000000;
	sram_mem[97868] = 16'b0000000000000000;
	sram_mem[97869] = 16'b0000000000000000;
	sram_mem[97870] = 16'b0000000000000000;
	sram_mem[97871] = 16'b0000000000000000;
	sram_mem[97872] = 16'b0000000000000000;
	sram_mem[97873] = 16'b0000000000000000;
	sram_mem[97874] = 16'b0000000000000000;
	sram_mem[97875] = 16'b0000000000000000;
	sram_mem[97876] = 16'b0000000000000000;
	sram_mem[97877] = 16'b0000000000000000;
	sram_mem[97878] = 16'b0000000000000000;
	sram_mem[97879] = 16'b0000000000000000;
	sram_mem[97880] = 16'b0000000000000000;
	sram_mem[97881] = 16'b0000000000000000;
	sram_mem[97882] = 16'b0000000000000000;
	sram_mem[97883] = 16'b0000000000000000;
	sram_mem[97884] = 16'b0000000000000000;
	sram_mem[97885] = 16'b0000000000000000;
	sram_mem[97886] = 16'b0000000000000000;
	sram_mem[97887] = 16'b0000000000000000;
	sram_mem[97888] = 16'b0000000000000000;
	sram_mem[97889] = 16'b0000000000000000;
	sram_mem[97890] = 16'b0000000000000000;
	sram_mem[97891] = 16'b0000000000000000;
	sram_mem[97892] = 16'b0000000000000000;
	sram_mem[97893] = 16'b0000000000000000;
	sram_mem[97894] = 16'b0000000000000000;
	sram_mem[97895] = 16'b0000000000000000;
	sram_mem[97896] = 16'b0000000000000000;
	sram_mem[97897] = 16'b0000000000000000;
	sram_mem[97898] = 16'b0000000000000000;
	sram_mem[97899] = 16'b0000000000000000;
	sram_mem[97900] = 16'b0000000000000000;
	sram_mem[97901] = 16'b0000000000000000;
	sram_mem[97902] = 16'b0000000000000000;
	sram_mem[97903] = 16'b0000000000000000;
	sram_mem[97904] = 16'b0000000000000000;
	sram_mem[97905] = 16'b0000000000000000;
	sram_mem[97906] = 16'b0000000000000000;
	sram_mem[97907] = 16'b0000000000000000;
	sram_mem[97908] = 16'b0000000000000000;
	sram_mem[97909] = 16'b0000000000000000;
	sram_mem[97910] = 16'b0000000000000000;
	sram_mem[97911] = 16'b0000000000000000;
	sram_mem[97912] = 16'b0000000000000000;
	sram_mem[97913] = 16'b0000000000000000;
	sram_mem[97914] = 16'b0000000000000000;
	sram_mem[97915] = 16'b0000000000000000;
	sram_mem[97916] = 16'b0000000000000000;
	sram_mem[97917] = 16'b0000000000000000;
	sram_mem[97918] = 16'b0000000000000000;
	sram_mem[97919] = 16'b0000000000000000;
	sram_mem[97920] = 16'b0000000000000000;
	sram_mem[97921] = 16'b0000000000000000;
	sram_mem[97922] = 16'b0000000000000000;
	sram_mem[97923] = 16'b0000000000000000;
	sram_mem[97924] = 16'b0000000000000000;
	sram_mem[97925] = 16'b0000000000000000;
	sram_mem[97926] = 16'b0000000000000000;
	sram_mem[97927] = 16'b0000000000000000;
	sram_mem[97928] = 16'b0000000000000000;
	sram_mem[97929] = 16'b0000000000000000;
	sram_mem[97930] = 16'b0000000000000000;
	sram_mem[97931] = 16'b0000000000000000;
	sram_mem[97932] = 16'b0000000000000000;
	sram_mem[97933] = 16'b0000000000000000;
	sram_mem[97934] = 16'b0000000000000000;
	sram_mem[97935] = 16'b0000000000000000;
	sram_mem[97936] = 16'b0000000000000000;
	sram_mem[97937] = 16'b0000000000000000;
	sram_mem[97938] = 16'b0000000000000000;
	sram_mem[97939] = 16'b0000000000000000;
	sram_mem[97940] = 16'b0000000000000000;
	sram_mem[97941] = 16'b0000000000000000;
	sram_mem[97942] = 16'b0000000000000000;
	sram_mem[97943] = 16'b0000000000000000;
	sram_mem[97944] = 16'b0000000000000000;
	sram_mem[97945] = 16'b0000000000000000;
	sram_mem[97946] = 16'b0000000000000000;
	sram_mem[97947] = 16'b0000000000000000;
	sram_mem[97948] = 16'b0000000000000000;
	sram_mem[97949] = 16'b0000000000000000;
	sram_mem[97950] = 16'b0000000000000000;
	sram_mem[97951] = 16'b0000000000000000;
	sram_mem[97952] = 16'b0000000000000000;
	sram_mem[97953] = 16'b0000000000000000;
	sram_mem[97954] = 16'b0000000000000000;
	sram_mem[97955] = 16'b0000000000000000;
	sram_mem[97956] = 16'b0000000000000000;
	sram_mem[97957] = 16'b0000000000000000;
	sram_mem[97958] = 16'b0000000000000000;
	sram_mem[97959] = 16'b0000000000000000;
	sram_mem[97960] = 16'b0000000000000000;
	sram_mem[97961] = 16'b0000000000000000;
	sram_mem[97962] = 16'b0000000000000000;
	sram_mem[97963] = 16'b0000000000000000;
	sram_mem[97964] = 16'b0000000000000000;
	sram_mem[97965] = 16'b0000000000000000;
	sram_mem[97966] = 16'b0000000000000000;
	sram_mem[97967] = 16'b0000000000000000;
	sram_mem[97968] = 16'b0000000000000000;
	sram_mem[97969] = 16'b0000000000000000;
	sram_mem[97970] = 16'b0000000000000000;
	sram_mem[97971] = 16'b0000000000000000;
	sram_mem[97972] = 16'b0000000000000000;
	sram_mem[97973] = 16'b0000000000000000;
	sram_mem[97974] = 16'b0000000000000000;
	sram_mem[97975] = 16'b0000000000000000;
	sram_mem[97976] = 16'b0000000000000000;
	sram_mem[97977] = 16'b0000000000000000;
	sram_mem[97978] = 16'b0000000000000000;
	sram_mem[97979] = 16'b0000000000000000;
	sram_mem[97980] = 16'b0000000000000000;
	sram_mem[97981] = 16'b0000000000000000;
	sram_mem[97982] = 16'b0000000000000000;
	sram_mem[97983] = 16'b0000000000000000;
	sram_mem[97984] = 16'b0000000000000000;
	sram_mem[97985] = 16'b0000000000000000;
	sram_mem[97986] = 16'b0000000000000000;
	sram_mem[97987] = 16'b0000000000000000;
	sram_mem[97988] = 16'b0000000000000000;
	sram_mem[97989] = 16'b0000000000000000;
	sram_mem[97990] = 16'b0000000000000000;
	sram_mem[97991] = 16'b0000000000000000;
	sram_mem[97992] = 16'b0000000000000000;
	sram_mem[97993] = 16'b0000000000000000;
	sram_mem[97994] = 16'b0000000000000000;
	sram_mem[97995] = 16'b0000000000000000;
	sram_mem[97996] = 16'b0000000000000000;
	sram_mem[97997] = 16'b0000000000000000;
	sram_mem[97998] = 16'b0000000000000000;
	sram_mem[97999] = 16'b0000000000000000;
	sram_mem[98000] = 16'b0000000000000000;
	sram_mem[98001] = 16'b0000000000000000;
	sram_mem[98002] = 16'b0000000000000000;
	sram_mem[98003] = 16'b0000000000000000;
	sram_mem[98004] = 16'b0000000000000000;
	sram_mem[98005] = 16'b0000000000000000;
	sram_mem[98006] = 16'b0000000000000000;
	sram_mem[98007] = 16'b0000000000000000;
	sram_mem[98008] = 16'b0000000000000000;
	sram_mem[98009] = 16'b0000000000000000;
	sram_mem[98010] = 16'b0000000000000000;
	sram_mem[98011] = 16'b0000000000000000;
	sram_mem[98012] = 16'b0000000000000000;
	sram_mem[98013] = 16'b0000000000000000;
	sram_mem[98014] = 16'b0000000000000000;
	sram_mem[98015] = 16'b0000000000000000;
	sram_mem[98016] = 16'b0000000000000000;
	sram_mem[98017] = 16'b0000000000000000;
	sram_mem[98018] = 16'b0000000000000000;
	sram_mem[98019] = 16'b0000000000000000;
	sram_mem[98020] = 16'b0000000000000000;
	sram_mem[98021] = 16'b0000000000000000;
	sram_mem[98022] = 16'b0000000000000000;
	sram_mem[98023] = 16'b0000000000000000;
	sram_mem[98024] = 16'b0000000000000000;
	sram_mem[98025] = 16'b0000000000000000;
	sram_mem[98026] = 16'b0000000000000000;
	sram_mem[98027] = 16'b0000000000000000;
	sram_mem[98028] = 16'b0000000000000000;
	sram_mem[98029] = 16'b0000000000000000;
	sram_mem[98030] = 16'b0000000000000000;
	sram_mem[98031] = 16'b0000000000000000;
	sram_mem[98032] = 16'b0000000000000000;
	sram_mem[98033] = 16'b0000000000000000;
	sram_mem[98034] = 16'b0000000000000000;
	sram_mem[98035] = 16'b0000000000000000;
	sram_mem[98036] = 16'b0000000000000000;
	sram_mem[98037] = 16'b0000000000000000;
	sram_mem[98038] = 16'b0000000000000000;
	sram_mem[98039] = 16'b0000000000000000;
	sram_mem[98040] = 16'b0000000000000000;
	sram_mem[98041] = 16'b0000000000000000;
	sram_mem[98042] = 16'b0000000000000000;
	sram_mem[98043] = 16'b0000000000000000;
	sram_mem[98044] = 16'b0000000000000000;
	sram_mem[98045] = 16'b0000000000000000;
	sram_mem[98046] = 16'b0000000000000000;
	sram_mem[98047] = 16'b0000000000000000;
	sram_mem[98048] = 16'b0000000000000000;
	sram_mem[98049] = 16'b0000000000000000;
	sram_mem[98050] = 16'b0000000000000000;
	sram_mem[98051] = 16'b0000000000000000;
	sram_mem[98052] = 16'b0000000000000000;
	sram_mem[98053] = 16'b0000000000000000;
	sram_mem[98054] = 16'b0000000000000000;
	sram_mem[98055] = 16'b0000000000000000;
	sram_mem[98056] = 16'b0000000000000000;
	sram_mem[98057] = 16'b0000000000000000;
	sram_mem[98058] = 16'b0000000000000000;
	sram_mem[98059] = 16'b0000000000000000;
	sram_mem[98060] = 16'b0000000000000000;
	sram_mem[98061] = 16'b0000000000000000;
	sram_mem[98062] = 16'b0000000000000000;
	sram_mem[98063] = 16'b0000000000000000;
	sram_mem[98064] = 16'b0000000000000000;
	sram_mem[98065] = 16'b0000000000000000;
	sram_mem[98066] = 16'b0000000000000000;
	sram_mem[98067] = 16'b0000000000000000;
	sram_mem[98068] = 16'b0000000000000000;
	sram_mem[98069] = 16'b0000000000000000;
	sram_mem[98070] = 16'b0000000000000000;
	sram_mem[98071] = 16'b0000000000000000;
	sram_mem[98072] = 16'b0000000000000000;
	sram_mem[98073] = 16'b0000000000000000;
	sram_mem[98074] = 16'b0000000000000000;
	sram_mem[98075] = 16'b0000000000000000;
	sram_mem[98076] = 16'b0000000000000000;
	sram_mem[98077] = 16'b0000000000000000;
	sram_mem[98078] = 16'b0000000000000000;
	sram_mem[98079] = 16'b0000000000000000;
	sram_mem[98080] = 16'b0000000000000000;
	sram_mem[98081] = 16'b0000000000000000;
	sram_mem[98082] = 16'b0000000000000000;
	sram_mem[98083] = 16'b0000000000000000;
	sram_mem[98084] = 16'b0000000000000000;
	sram_mem[98085] = 16'b0000000000000000;
	sram_mem[98086] = 16'b0000000000000000;
	sram_mem[98087] = 16'b0000000000000000;
	sram_mem[98088] = 16'b0000000000000000;
	sram_mem[98089] = 16'b0000000000000000;
	sram_mem[98090] = 16'b0000000000000000;
	sram_mem[98091] = 16'b0000000000000000;
	sram_mem[98092] = 16'b0000000000000000;
	sram_mem[98093] = 16'b0000000000000000;
	sram_mem[98094] = 16'b0000000000000000;
	sram_mem[98095] = 16'b0000000000000000;
	sram_mem[98096] = 16'b0000000000000000;
	sram_mem[98097] = 16'b0000000000000000;
	sram_mem[98098] = 16'b0000000000000000;
	sram_mem[98099] = 16'b0000000000000000;
	sram_mem[98100] = 16'b0000000000000000;
	sram_mem[98101] = 16'b0000000000000000;
	sram_mem[98102] = 16'b0000000000000000;
	sram_mem[98103] = 16'b0000000000000000;
	sram_mem[98104] = 16'b0000000000000000;
	sram_mem[98105] = 16'b0000000000000000;
	sram_mem[98106] = 16'b0000000000000000;
	sram_mem[98107] = 16'b0000000000000000;
	sram_mem[98108] = 16'b0000000000000000;
	sram_mem[98109] = 16'b0000000000000000;
	sram_mem[98110] = 16'b0000000000000000;
	sram_mem[98111] = 16'b0000000000000000;
	sram_mem[98112] = 16'b0000000000000000;
	sram_mem[98113] = 16'b0000000000000000;
	sram_mem[98114] = 16'b0000000000000000;
	sram_mem[98115] = 16'b0000000000000000;
	sram_mem[98116] = 16'b0000000000000000;
	sram_mem[98117] = 16'b0000000000000000;
	sram_mem[98118] = 16'b0000000000000000;
	sram_mem[98119] = 16'b0000000000000000;
	sram_mem[98120] = 16'b0000000000000000;
	sram_mem[98121] = 16'b0000000000000000;
	sram_mem[98122] = 16'b0000000000000000;
	sram_mem[98123] = 16'b0000000000000000;
	sram_mem[98124] = 16'b0000000000000000;
	sram_mem[98125] = 16'b0000000000000000;
	sram_mem[98126] = 16'b0000000000000000;
	sram_mem[98127] = 16'b0000000000000000;
	sram_mem[98128] = 16'b0000000000000000;
	sram_mem[98129] = 16'b0000000000000000;
	sram_mem[98130] = 16'b0000000000000000;
	sram_mem[98131] = 16'b0000000000000000;
	sram_mem[98132] = 16'b0000000000000000;
	sram_mem[98133] = 16'b0000000000000000;
	sram_mem[98134] = 16'b0000000000000000;
	sram_mem[98135] = 16'b0000000000000000;
	sram_mem[98136] = 16'b0000000000000000;
	sram_mem[98137] = 16'b0000000000000000;
	sram_mem[98138] = 16'b0000000000000000;
	sram_mem[98139] = 16'b0000000000000000;
	sram_mem[98140] = 16'b0000000000000000;
	sram_mem[98141] = 16'b0000000000000000;
	sram_mem[98142] = 16'b0000000000000000;
	sram_mem[98143] = 16'b0000000000000000;
	sram_mem[98144] = 16'b0000000000000000;
	sram_mem[98145] = 16'b0000000000000000;
	sram_mem[98146] = 16'b0000000000000000;
	sram_mem[98147] = 16'b0000000000000000;
	sram_mem[98148] = 16'b0000000000000000;
	sram_mem[98149] = 16'b0000000000000000;
	sram_mem[98150] = 16'b0000000000000000;
	sram_mem[98151] = 16'b0000000000000000;
	sram_mem[98152] = 16'b0000000000000000;
	sram_mem[98153] = 16'b0000000000000000;
	sram_mem[98154] = 16'b0000000000000000;
	sram_mem[98155] = 16'b0000000000000000;
	sram_mem[98156] = 16'b0000000000000000;
	sram_mem[98157] = 16'b0000000000000000;
	sram_mem[98158] = 16'b0000000000000000;
	sram_mem[98159] = 16'b0000000000000000;
	sram_mem[98160] = 16'b0000000000000000;
	sram_mem[98161] = 16'b0000000000000000;
	sram_mem[98162] = 16'b0000000000000000;
	sram_mem[98163] = 16'b0000000000000000;
	sram_mem[98164] = 16'b0000000000000000;
	sram_mem[98165] = 16'b0000000000000000;
	sram_mem[98166] = 16'b0000000000000000;
	sram_mem[98167] = 16'b0000000000000000;
	sram_mem[98168] = 16'b0000000000000000;
	sram_mem[98169] = 16'b0000000000000000;
	sram_mem[98170] = 16'b0000000000000000;
	sram_mem[98171] = 16'b0000000000000000;
	sram_mem[98172] = 16'b0000000000000000;
	sram_mem[98173] = 16'b0000000000000000;
	sram_mem[98174] = 16'b0000000000000000;
	sram_mem[98175] = 16'b0000000000000000;
	sram_mem[98176] = 16'b0000000000000000;
	sram_mem[98177] = 16'b0000000000000000;
	sram_mem[98178] = 16'b0000000000000000;
	sram_mem[98179] = 16'b0000000000000000;
	sram_mem[98180] = 16'b0000000000000000;
	sram_mem[98181] = 16'b0000000000000000;
	sram_mem[98182] = 16'b0000000000000000;
	sram_mem[98183] = 16'b0000000000000000;
	sram_mem[98184] = 16'b0000000000000000;
	sram_mem[98185] = 16'b0000000000000000;
	sram_mem[98186] = 16'b0000000000000000;
	sram_mem[98187] = 16'b0000000000000000;
	sram_mem[98188] = 16'b0000000000000000;
	sram_mem[98189] = 16'b0000000000000000;
	sram_mem[98190] = 16'b0000000000000000;
	sram_mem[98191] = 16'b0000000000000000;
	sram_mem[98192] = 16'b0000000000000000;
	sram_mem[98193] = 16'b0000000000000000;
	sram_mem[98194] = 16'b0000000000000000;
	sram_mem[98195] = 16'b0000000000000000;
	sram_mem[98196] = 16'b0000000000000000;
	sram_mem[98197] = 16'b0000000000000000;
	sram_mem[98198] = 16'b0000000000000000;
	sram_mem[98199] = 16'b0000000000000000;
	sram_mem[98200] = 16'b0000000000000000;
	sram_mem[98201] = 16'b0000000000000000;
	sram_mem[98202] = 16'b0000000000000000;
	sram_mem[98203] = 16'b0000000000000000;
	sram_mem[98204] = 16'b0000000000000000;
	sram_mem[98205] = 16'b0000000000000000;
	sram_mem[98206] = 16'b0000000000000000;
	sram_mem[98207] = 16'b0000000000000000;
	sram_mem[98208] = 16'b0000000000000000;
	sram_mem[98209] = 16'b0000000000000000;
	sram_mem[98210] = 16'b0000000000000000;
	sram_mem[98211] = 16'b0000000000000000;
	sram_mem[98212] = 16'b0000000000000000;
	sram_mem[98213] = 16'b0000000000000000;
	sram_mem[98214] = 16'b0000000000000000;
	sram_mem[98215] = 16'b0000000000000000;
	sram_mem[98216] = 16'b0000000000000000;
	sram_mem[98217] = 16'b0000000000000000;
	sram_mem[98218] = 16'b0000000000000000;
	sram_mem[98219] = 16'b0000000000000000;
	sram_mem[98220] = 16'b0000000000000000;
	sram_mem[98221] = 16'b0000000000000000;
	sram_mem[98222] = 16'b0000000000000000;
	sram_mem[98223] = 16'b0000000000000000;
	sram_mem[98224] = 16'b0000000000000000;
	sram_mem[98225] = 16'b0000000000000000;
	sram_mem[98226] = 16'b0000000000000000;
	sram_mem[98227] = 16'b0000000000000000;
	sram_mem[98228] = 16'b0000000000000000;
	sram_mem[98229] = 16'b0000000000000000;
	sram_mem[98230] = 16'b0000000000000000;
	sram_mem[98231] = 16'b0000000000000000;
	sram_mem[98232] = 16'b0000000000000000;
	sram_mem[98233] = 16'b0000000000000000;
	sram_mem[98234] = 16'b0000000000000000;
	sram_mem[98235] = 16'b0000000000000000;
	sram_mem[98236] = 16'b0000000000000000;
	sram_mem[98237] = 16'b0000000000000000;
	sram_mem[98238] = 16'b0000000000000000;
	sram_mem[98239] = 16'b0000000000000000;
	sram_mem[98240] = 16'b0000000000000000;
	sram_mem[98241] = 16'b0000000000000000;
	sram_mem[98242] = 16'b0000000000000000;
	sram_mem[98243] = 16'b0000000000000000;
	sram_mem[98244] = 16'b0000000000000000;
	sram_mem[98245] = 16'b0000000000000000;
	sram_mem[98246] = 16'b0000000000000000;
	sram_mem[98247] = 16'b0000000000000000;
	sram_mem[98248] = 16'b0000000000000000;
	sram_mem[98249] = 16'b0000000000000000;
	sram_mem[98250] = 16'b0000000000000000;
	sram_mem[98251] = 16'b0000000000000000;
	sram_mem[98252] = 16'b0000000000000000;
	sram_mem[98253] = 16'b0000000000000000;
	sram_mem[98254] = 16'b0000000000000000;
	sram_mem[98255] = 16'b0000000000000000;
	sram_mem[98256] = 16'b0000000000000000;
	sram_mem[98257] = 16'b0000000000000000;
	sram_mem[98258] = 16'b0000000000000000;
	sram_mem[98259] = 16'b0000000000000000;
	sram_mem[98260] = 16'b0000000000000000;
	sram_mem[98261] = 16'b0000000000000000;
	sram_mem[98262] = 16'b0000000000000000;
	sram_mem[98263] = 16'b0000000000000000;
	sram_mem[98264] = 16'b0000000000000000;
	sram_mem[98265] = 16'b0000000000000000;
	sram_mem[98266] = 16'b0000000000000000;
	sram_mem[98267] = 16'b0000000000000000;
	sram_mem[98268] = 16'b0000000000000000;
	sram_mem[98269] = 16'b0000000000000000;
	sram_mem[98270] = 16'b0000000000000000;
	sram_mem[98271] = 16'b0000000000000000;
	sram_mem[98272] = 16'b0000000000000000;
	sram_mem[98273] = 16'b0000000000000000;
	sram_mem[98274] = 16'b0000000000000000;
	sram_mem[98275] = 16'b0000000000000000;
	sram_mem[98276] = 16'b0000000000000000;
	sram_mem[98277] = 16'b0000000000000000;
	sram_mem[98278] = 16'b0000000000000000;
	sram_mem[98279] = 16'b0000000000000000;
	sram_mem[98280] = 16'b0000000000000000;
	sram_mem[98281] = 16'b0000000000000000;
	sram_mem[98282] = 16'b0000000000000000;
	sram_mem[98283] = 16'b0000000000000000;
	sram_mem[98284] = 16'b0000000000000000;
	sram_mem[98285] = 16'b0000000000000000;
	sram_mem[98286] = 16'b0000000000000000;
	sram_mem[98287] = 16'b0000000000000000;
	sram_mem[98288] = 16'b0000000000000000;
	sram_mem[98289] = 16'b0000000000000000;
	sram_mem[98290] = 16'b0000000000000000;
	sram_mem[98291] = 16'b0000000000000000;
	sram_mem[98292] = 16'b0000000000000000;
	sram_mem[98293] = 16'b0000000000000000;
	sram_mem[98294] = 16'b0000000000000000;
	sram_mem[98295] = 16'b0000000000000000;
	sram_mem[98296] = 16'b0000000000000000;
	sram_mem[98297] = 16'b0000000000000000;
	sram_mem[98298] = 16'b0000000000000000;
	sram_mem[98299] = 16'b0000000000000000;
	sram_mem[98300] = 16'b0000000000000000;
	sram_mem[98301] = 16'b0000000000000000;
	sram_mem[98302] = 16'b0000000000000000;
	sram_mem[98303] = 16'b0000000000000000;
	sram_mem[98304] = 16'b0000000000000000;
	sram_mem[98305] = 16'b0000000000000000;
	sram_mem[98306] = 16'b0000000000000000;
	sram_mem[98307] = 16'b0000000000000000;
	sram_mem[98308] = 16'b0000000000000000;
	sram_mem[98309] = 16'b0000000000000000;
	sram_mem[98310] = 16'b0000000000000000;
	sram_mem[98311] = 16'b0000000000000000;
	sram_mem[98312] = 16'b0000000000000000;
	sram_mem[98313] = 16'b0000000000000000;
	sram_mem[98314] = 16'b0000000000000000;
	sram_mem[98315] = 16'b0000000000000000;
	sram_mem[98316] = 16'b0000000000000000;
	sram_mem[98317] = 16'b0000000000000000;
	sram_mem[98318] = 16'b0000000000000000;
	sram_mem[98319] = 16'b0000000000000000;
	sram_mem[98320] = 16'b0000000000000000;
	sram_mem[98321] = 16'b0000000000000000;
	sram_mem[98322] = 16'b0000000000000000;
	sram_mem[98323] = 16'b0000000000000000;
	sram_mem[98324] = 16'b0000000000000000;
	sram_mem[98325] = 16'b0000000000000000;
	sram_mem[98326] = 16'b0000000000000000;
	sram_mem[98327] = 16'b0000000000000000;
	sram_mem[98328] = 16'b0000000000000000;
	sram_mem[98329] = 16'b0000000000000000;
	sram_mem[98330] = 16'b0000000000000000;
	sram_mem[98331] = 16'b0000000000000000;
	sram_mem[98332] = 16'b0000000000000000;
	sram_mem[98333] = 16'b0000000000000000;
	sram_mem[98334] = 16'b0000000000000000;
	sram_mem[98335] = 16'b0000000000000000;
	sram_mem[98336] = 16'b0000000000000000;
	sram_mem[98337] = 16'b0000000000000000;
	sram_mem[98338] = 16'b0000000000000000;
	sram_mem[98339] = 16'b0000000000000000;
	sram_mem[98340] = 16'b0000000000000000;
	sram_mem[98341] = 16'b0000000000000000;
	sram_mem[98342] = 16'b0000000000000000;
	sram_mem[98343] = 16'b0000000000000000;
	sram_mem[98344] = 16'b0000000000000000;
	sram_mem[98345] = 16'b0000000000000000;
	sram_mem[98346] = 16'b0000000000000000;
	sram_mem[98347] = 16'b0000000000000000;
	sram_mem[98348] = 16'b0000000000000000;
	sram_mem[98349] = 16'b0000000000000000;
	sram_mem[98350] = 16'b0000000000000000;
	sram_mem[98351] = 16'b0000000000000000;
	sram_mem[98352] = 16'b0000000000000000;
	sram_mem[98353] = 16'b0000000000000000;
	sram_mem[98354] = 16'b0000000000000000;
	sram_mem[98355] = 16'b0000000000000000;
	sram_mem[98356] = 16'b0000000000000000;
	sram_mem[98357] = 16'b0000000000000000;
	sram_mem[98358] = 16'b0000000000000000;
	sram_mem[98359] = 16'b0000000000000000;
	sram_mem[98360] = 16'b0000000000000000;
	sram_mem[98361] = 16'b0000000000000000;
	sram_mem[98362] = 16'b0000000000000000;
	sram_mem[98363] = 16'b0000000000000000;
	sram_mem[98364] = 16'b0000000000000000;
	sram_mem[98365] = 16'b0000000000000000;
	sram_mem[98366] = 16'b0000000000000000;
	sram_mem[98367] = 16'b0000000000000000;
	sram_mem[98368] = 16'b0000000000000000;
	sram_mem[98369] = 16'b0000000000000000;
	sram_mem[98370] = 16'b0000000000000000;
	sram_mem[98371] = 16'b0000000000000000;
	sram_mem[98372] = 16'b0000000000000000;
	sram_mem[98373] = 16'b0000000000000000;
	sram_mem[98374] = 16'b0000000000000000;
	sram_mem[98375] = 16'b0000000000000000;
	sram_mem[98376] = 16'b0000000000000000;
	sram_mem[98377] = 16'b0000000000000000;
	sram_mem[98378] = 16'b0000000000000000;
	sram_mem[98379] = 16'b0000000000000000;
	sram_mem[98380] = 16'b0000000000000000;
	sram_mem[98381] = 16'b0000000000000000;
	sram_mem[98382] = 16'b0000000000000000;
	sram_mem[98383] = 16'b0000000000000000;
	sram_mem[98384] = 16'b0000000000000000;
	sram_mem[98385] = 16'b0000000000000000;
	sram_mem[98386] = 16'b0000000000000000;
	sram_mem[98387] = 16'b0000000000000000;
	sram_mem[98388] = 16'b0000000000000000;
	sram_mem[98389] = 16'b0000000000000000;
	sram_mem[98390] = 16'b0000000000000000;
	sram_mem[98391] = 16'b0000000000000000;
	sram_mem[98392] = 16'b0000000000000000;
	sram_mem[98393] = 16'b0000000000000000;
	sram_mem[98394] = 16'b0000000000000000;
	sram_mem[98395] = 16'b0000000000000000;
	sram_mem[98396] = 16'b0000000000000000;
	sram_mem[98397] = 16'b0000000000000000;
	sram_mem[98398] = 16'b0000000000000000;
	sram_mem[98399] = 16'b0000000000000000;
	sram_mem[98400] = 16'b0000000000000000;
	sram_mem[98401] = 16'b0000000000000000;
	sram_mem[98402] = 16'b0000000000000000;
	sram_mem[98403] = 16'b0000000000000000;
	sram_mem[98404] = 16'b0000000000000000;
	sram_mem[98405] = 16'b0000000000000000;
	sram_mem[98406] = 16'b0000000000000000;
	sram_mem[98407] = 16'b0000000000000000;
	sram_mem[98408] = 16'b0000000000000000;
	sram_mem[98409] = 16'b0000000000000000;
	sram_mem[98410] = 16'b0000000000000000;
	sram_mem[98411] = 16'b0000000000000000;
	sram_mem[98412] = 16'b0000000000000000;
	sram_mem[98413] = 16'b0000000000000000;
	sram_mem[98414] = 16'b0000000000000000;
	sram_mem[98415] = 16'b0000000000000000;
	sram_mem[98416] = 16'b0000000000000000;
	sram_mem[98417] = 16'b0000000000000000;
	sram_mem[98418] = 16'b0000000000000000;
	sram_mem[98419] = 16'b0000000000000000;
	sram_mem[98420] = 16'b0000000000000000;
	sram_mem[98421] = 16'b0000000000000000;
	sram_mem[98422] = 16'b0000000000000000;
	sram_mem[98423] = 16'b0000000000000000;
	sram_mem[98424] = 16'b0000000000000000;
	sram_mem[98425] = 16'b0000000000000000;
	sram_mem[98426] = 16'b0000000000000000;
	sram_mem[98427] = 16'b0000000000000000;
	sram_mem[98428] = 16'b0000000000000000;
	sram_mem[98429] = 16'b0000000000000000;
	sram_mem[98430] = 16'b0000000000000000;
	sram_mem[98431] = 16'b0000000000000000;
	sram_mem[98432] = 16'b0000000000000000;
	sram_mem[98433] = 16'b0000000000000000;
	sram_mem[98434] = 16'b0000000000000000;
	sram_mem[98435] = 16'b0000000000000000;
	sram_mem[98436] = 16'b0000000000000000;
	sram_mem[98437] = 16'b0000000000000000;
	sram_mem[98438] = 16'b0000000000000000;
	sram_mem[98439] = 16'b0000000000000000;
	sram_mem[98440] = 16'b0000000000000000;
	sram_mem[98441] = 16'b0000000000000000;
	sram_mem[98442] = 16'b0000000000000000;
	sram_mem[98443] = 16'b0000000000000000;
	sram_mem[98444] = 16'b0000000000000000;
	sram_mem[98445] = 16'b0000000000000000;
	sram_mem[98446] = 16'b0000000000000000;
	sram_mem[98447] = 16'b0000000000000000;
	sram_mem[98448] = 16'b0000000000000000;
	sram_mem[98449] = 16'b0000000000000000;
	sram_mem[98450] = 16'b0000000000000000;
	sram_mem[98451] = 16'b0000000000000000;
	sram_mem[98452] = 16'b0000000000000000;
	sram_mem[98453] = 16'b0000000000000000;
	sram_mem[98454] = 16'b0000000000000000;
	sram_mem[98455] = 16'b0000000000000000;
	sram_mem[98456] = 16'b0000000000000000;
	sram_mem[98457] = 16'b0000000000000000;
	sram_mem[98458] = 16'b0000000000000000;
	sram_mem[98459] = 16'b0000000000000000;
	sram_mem[98460] = 16'b0000000000000000;
	sram_mem[98461] = 16'b0000000000000000;
	sram_mem[98462] = 16'b0000000000000000;
	sram_mem[98463] = 16'b0000000000000000;
	sram_mem[98464] = 16'b0000000000000000;
	sram_mem[98465] = 16'b0000000000000000;
	sram_mem[98466] = 16'b0000000000000000;
	sram_mem[98467] = 16'b0000000000000000;
	sram_mem[98468] = 16'b0000000000000000;
	sram_mem[98469] = 16'b0000000000000000;
	sram_mem[98470] = 16'b0000000000000000;
	sram_mem[98471] = 16'b0000000000000000;
	sram_mem[98472] = 16'b0000000000000000;
	sram_mem[98473] = 16'b0000000000000000;
	sram_mem[98474] = 16'b0000000000000000;
	sram_mem[98475] = 16'b0000000000000000;
	sram_mem[98476] = 16'b0000000000000000;
	sram_mem[98477] = 16'b0000000000000000;
	sram_mem[98478] = 16'b0000000000000000;
	sram_mem[98479] = 16'b0000000000000000;
	sram_mem[98480] = 16'b0000000000000000;
	sram_mem[98481] = 16'b0000000000000000;
	sram_mem[98482] = 16'b0000000000000000;
	sram_mem[98483] = 16'b0000000000000000;
	sram_mem[98484] = 16'b0000000000000000;
	sram_mem[98485] = 16'b0000000000000000;
	sram_mem[98486] = 16'b0000000000000000;
	sram_mem[98487] = 16'b0000000000000000;
	sram_mem[98488] = 16'b0000000000000000;
	sram_mem[98489] = 16'b0000000000000000;
	sram_mem[98490] = 16'b0000000000000000;
	sram_mem[98491] = 16'b0000000000000000;
	sram_mem[98492] = 16'b0000000000000000;
	sram_mem[98493] = 16'b0000000000000000;
	sram_mem[98494] = 16'b0000000000000000;
	sram_mem[98495] = 16'b0000000000000000;
	sram_mem[98496] = 16'b0000000000000000;
	sram_mem[98497] = 16'b0000000000000000;
	sram_mem[98498] = 16'b0000000000000000;
	sram_mem[98499] = 16'b0000000000000000;
	sram_mem[98500] = 16'b0000000000000000;
	sram_mem[98501] = 16'b0000000000000000;
	sram_mem[98502] = 16'b0000000000000000;
	sram_mem[98503] = 16'b0000000000000000;
	sram_mem[98504] = 16'b0000000000000000;
	sram_mem[98505] = 16'b0000000000000000;
	sram_mem[98506] = 16'b0000000000000000;
	sram_mem[98507] = 16'b0000000000000000;
	sram_mem[98508] = 16'b0000000000000000;
	sram_mem[98509] = 16'b0000000000000000;
	sram_mem[98510] = 16'b0000000000000000;
	sram_mem[98511] = 16'b0000000000000000;
	sram_mem[98512] = 16'b0000000000000000;
	sram_mem[98513] = 16'b0000000000000000;
	sram_mem[98514] = 16'b0000000000000000;
	sram_mem[98515] = 16'b0000000000000000;
	sram_mem[98516] = 16'b0000000000000000;
	sram_mem[98517] = 16'b0000000000000000;
	sram_mem[98518] = 16'b0000000000000000;
	sram_mem[98519] = 16'b0000000000000000;
	sram_mem[98520] = 16'b0000000000000000;
	sram_mem[98521] = 16'b0000000000000000;
	sram_mem[98522] = 16'b0000000000000000;
	sram_mem[98523] = 16'b0000000000000000;
	sram_mem[98524] = 16'b0000000000000000;
	sram_mem[98525] = 16'b0000000000000000;
	sram_mem[98526] = 16'b0000000000000000;
	sram_mem[98527] = 16'b0000000000000000;
	sram_mem[98528] = 16'b0000000000000000;
	sram_mem[98529] = 16'b0000000000000000;
	sram_mem[98530] = 16'b0000000000000000;
	sram_mem[98531] = 16'b0000000000000000;
	sram_mem[98532] = 16'b0000000000000000;
	sram_mem[98533] = 16'b0000000000000000;
	sram_mem[98534] = 16'b0000000000000000;
	sram_mem[98535] = 16'b0000000000000000;
	sram_mem[98536] = 16'b0000000000000000;
	sram_mem[98537] = 16'b0000000000000000;
	sram_mem[98538] = 16'b0000000000000000;
	sram_mem[98539] = 16'b0000000000000000;
	sram_mem[98540] = 16'b0000000000000000;
	sram_mem[98541] = 16'b0000000000000000;
	sram_mem[98542] = 16'b0000000000000000;
	sram_mem[98543] = 16'b0000000000000000;
	sram_mem[98544] = 16'b0000000000000000;
	sram_mem[98545] = 16'b0000000000000000;
	sram_mem[98546] = 16'b0000000000000000;
	sram_mem[98547] = 16'b0000000000000000;
	sram_mem[98548] = 16'b0000000000000000;
	sram_mem[98549] = 16'b0000000000000000;
	sram_mem[98550] = 16'b0000000000000000;
	sram_mem[98551] = 16'b0000000000000000;
	sram_mem[98552] = 16'b0000000000000000;
	sram_mem[98553] = 16'b0000000000000000;
	sram_mem[98554] = 16'b0000000000000000;
	sram_mem[98555] = 16'b0000000000000000;
	sram_mem[98556] = 16'b0000000000000000;
	sram_mem[98557] = 16'b0000000000000000;
	sram_mem[98558] = 16'b0000000000000000;
	sram_mem[98559] = 16'b0000000000000000;
	sram_mem[98560] = 16'b0000000000000000;
	sram_mem[98561] = 16'b0000000000000000;
	sram_mem[98562] = 16'b0000000000000000;
	sram_mem[98563] = 16'b0000000000000000;
	sram_mem[98564] = 16'b0000000000000000;
	sram_mem[98565] = 16'b0000000000000000;
	sram_mem[98566] = 16'b0000000000000000;
	sram_mem[98567] = 16'b0000000000000000;
	sram_mem[98568] = 16'b0000000000000000;
	sram_mem[98569] = 16'b0000000000000000;
	sram_mem[98570] = 16'b0000000000000000;
	sram_mem[98571] = 16'b0000000000000000;
	sram_mem[98572] = 16'b0000000000000000;
	sram_mem[98573] = 16'b0000000000000000;
	sram_mem[98574] = 16'b0000000000000000;
	sram_mem[98575] = 16'b0000000000000000;
	sram_mem[98576] = 16'b0000000000000000;
	sram_mem[98577] = 16'b0000000000000000;
	sram_mem[98578] = 16'b0000000000000000;
	sram_mem[98579] = 16'b0000000000000000;
	sram_mem[98580] = 16'b0000000000000000;
	sram_mem[98581] = 16'b0000000000000000;
	sram_mem[98582] = 16'b0000000000000000;
	sram_mem[98583] = 16'b0000000000000000;
	sram_mem[98584] = 16'b0000000000000000;
	sram_mem[98585] = 16'b0000000000000000;
	sram_mem[98586] = 16'b0000000000000000;
	sram_mem[98587] = 16'b0000000000000000;
	sram_mem[98588] = 16'b0000000000000000;
	sram_mem[98589] = 16'b0000000000000000;
	sram_mem[98590] = 16'b0000000000000000;
	sram_mem[98591] = 16'b0000000000000000;
	sram_mem[98592] = 16'b0000000000000000;
	sram_mem[98593] = 16'b0000000000000000;
	sram_mem[98594] = 16'b0000000000000000;
	sram_mem[98595] = 16'b0000000000000000;
	sram_mem[98596] = 16'b0000000000000000;
	sram_mem[98597] = 16'b0000000000000000;
	sram_mem[98598] = 16'b0000000000000000;
	sram_mem[98599] = 16'b0000000000000000;
	sram_mem[98600] = 16'b0000000000000000;
	sram_mem[98601] = 16'b0000000000000000;
	sram_mem[98602] = 16'b0000000000000000;
	sram_mem[98603] = 16'b0000000000000000;
	sram_mem[98604] = 16'b0000000000000000;
	sram_mem[98605] = 16'b0000000000000000;
	sram_mem[98606] = 16'b0000000000000000;
	sram_mem[98607] = 16'b0000000000000000;
	sram_mem[98608] = 16'b0000000000000000;
	sram_mem[98609] = 16'b0000000000000000;
	sram_mem[98610] = 16'b0000000000000000;
	sram_mem[98611] = 16'b0000000000000000;
	sram_mem[98612] = 16'b0000000000000000;
	sram_mem[98613] = 16'b0000000000000000;
	sram_mem[98614] = 16'b0000000000000000;
	sram_mem[98615] = 16'b0000000000000000;
	sram_mem[98616] = 16'b0000000000000000;
	sram_mem[98617] = 16'b0000000000000000;
	sram_mem[98618] = 16'b0000000000000000;
	sram_mem[98619] = 16'b0000000000000000;
	sram_mem[98620] = 16'b0000000000000000;
	sram_mem[98621] = 16'b0000000000000000;
	sram_mem[98622] = 16'b0000000000000000;
	sram_mem[98623] = 16'b0000000000000000;
	sram_mem[98624] = 16'b0000000000000000;
	sram_mem[98625] = 16'b0000000000000000;
	sram_mem[98626] = 16'b0000000000000000;
	sram_mem[98627] = 16'b0000000000000000;
	sram_mem[98628] = 16'b0000000000000000;
	sram_mem[98629] = 16'b0000000000000000;
	sram_mem[98630] = 16'b0000000000000000;
	sram_mem[98631] = 16'b0000000000000000;
	sram_mem[98632] = 16'b0000000000000000;
	sram_mem[98633] = 16'b0000000000000000;
	sram_mem[98634] = 16'b0000000000000000;
	sram_mem[98635] = 16'b0000000000000000;
	sram_mem[98636] = 16'b0000000000000000;
	sram_mem[98637] = 16'b0000000000000000;
	sram_mem[98638] = 16'b0000000000000000;
	sram_mem[98639] = 16'b0000000000000000;
	sram_mem[98640] = 16'b0000000000000000;
	sram_mem[98641] = 16'b0000000000000000;
	sram_mem[98642] = 16'b0000000000000000;
	sram_mem[98643] = 16'b0000000000000000;
	sram_mem[98644] = 16'b0000000000000000;
	sram_mem[98645] = 16'b0000000000000000;
	sram_mem[98646] = 16'b0000000000000000;
	sram_mem[98647] = 16'b0000000000000000;
	sram_mem[98648] = 16'b0000000000000000;
	sram_mem[98649] = 16'b0000000000000000;
	sram_mem[98650] = 16'b0000000000000000;
	sram_mem[98651] = 16'b0000000000000000;
	sram_mem[98652] = 16'b0000000000000000;
	sram_mem[98653] = 16'b0000000000000000;
	sram_mem[98654] = 16'b0000000000000000;
	sram_mem[98655] = 16'b0000000000000000;
	sram_mem[98656] = 16'b0000000000000000;
	sram_mem[98657] = 16'b0000000000000000;
	sram_mem[98658] = 16'b0000000000000000;
	sram_mem[98659] = 16'b0000000000000000;
	sram_mem[98660] = 16'b0000000000000000;
	sram_mem[98661] = 16'b0000000000000000;
	sram_mem[98662] = 16'b0000000000000000;
	sram_mem[98663] = 16'b0000000000000000;
	sram_mem[98664] = 16'b0000000000000000;
	sram_mem[98665] = 16'b0000000000000000;
	sram_mem[98666] = 16'b0000000000000000;
	sram_mem[98667] = 16'b0000000000000000;
	sram_mem[98668] = 16'b0000000000000000;
	sram_mem[98669] = 16'b0000000000000000;
	sram_mem[98670] = 16'b0000000000000000;
	sram_mem[98671] = 16'b0000000000000000;
	sram_mem[98672] = 16'b0000000000000000;
	sram_mem[98673] = 16'b0000000000000000;
	sram_mem[98674] = 16'b0000000000000000;
	sram_mem[98675] = 16'b0000000000000000;
	sram_mem[98676] = 16'b0000000000000000;
	sram_mem[98677] = 16'b0000000000000000;
	sram_mem[98678] = 16'b0000000000000000;
	sram_mem[98679] = 16'b0000000000000000;
	sram_mem[98680] = 16'b0000000000000000;
	sram_mem[98681] = 16'b0000000000000000;
	sram_mem[98682] = 16'b0000000000000000;
	sram_mem[98683] = 16'b0000000000000000;
	sram_mem[98684] = 16'b0000000000000000;
	sram_mem[98685] = 16'b0000000000000000;
	sram_mem[98686] = 16'b0000000000000000;
	sram_mem[98687] = 16'b0000000000000000;
	sram_mem[98688] = 16'b0000000000000000;
	sram_mem[98689] = 16'b0000000000000000;
	sram_mem[98690] = 16'b0000000000000000;
	sram_mem[98691] = 16'b0000000000000000;
	sram_mem[98692] = 16'b0000000000000000;
	sram_mem[98693] = 16'b0000000000000000;
	sram_mem[98694] = 16'b0000000000000000;
	sram_mem[98695] = 16'b0000000000000000;
	sram_mem[98696] = 16'b0000000000000000;
	sram_mem[98697] = 16'b0000000000000000;
	sram_mem[98698] = 16'b0000000000000000;
	sram_mem[98699] = 16'b0000000000000000;
	sram_mem[98700] = 16'b0000000000000000;
	sram_mem[98701] = 16'b0000000000000000;
	sram_mem[98702] = 16'b0000000000000000;
	sram_mem[98703] = 16'b0000000000000000;
	sram_mem[98704] = 16'b0000000000000000;
	sram_mem[98705] = 16'b0000000000000000;
	sram_mem[98706] = 16'b0000000000000000;
	sram_mem[98707] = 16'b0000000000000000;
	sram_mem[98708] = 16'b0000000000000000;
	sram_mem[98709] = 16'b0000000000000000;
	sram_mem[98710] = 16'b0000000000000000;
	sram_mem[98711] = 16'b0000000000000000;
	sram_mem[98712] = 16'b0000000000000000;
	sram_mem[98713] = 16'b0000000000000000;
	sram_mem[98714] = 16'b0000000000000000;
	sram_mem[98715] = 16'b0000000000000000;
	sram_mem[98716] = 16'b0000000000000000;
	sram_mem[98717] = 16'b0000000000000000;
	sram_mem[98718] = 16'b0000000000000000;
	sram_mem[98719] = 16'b0000000000000000;
	sram_mem[98720] = 16'b0000000000000000;
	sram_mem[98721] = 16'b0000000000000000;
	sram_mem[98722] = 16'b0000000000000000;
	sram_mem[98723] = 16'b0000000000000000;
	sram_mem[98724] = 16'b0000000000000000;
	sram_mem[98725] = 16'b0000000000000000;
	sram_mem[98726] = 16'b0000000000000000;
	sram_mem[98727] = 16'b0000000000000000;
	sram_mem[98728] = 16'b0000000000000000;
	sram_mem[98729] = 16'b0000000000000000;
	sram_mem[98730] = 16'b0000000000000000;
	sram_mem[98731] = 16'b0000000000000000;
	sram_mem[98732] = 16'b0000000000000000;
	sram_mem[98733] = 16'b0000000000000000;
	sram_mem[98734] = 16'b0000000000000000;
	sram_mem[98735] = 16'b0000000000000000;
	sram_mem[98736] = 16'b0000000000000000;
	sram_mem[98737] = 16'b0000000000000000;
	sram_mem[98738] = 16'b0000000000000000;
	sram_mem[98739] = 16'b0000000000000000;
	sram_mem[98740] = 16'b0000000000000000;
	sram_mem[98741] = 16'b0000000000000000;
	sram_mem[98742] = 16'b0000000000000000;
	sram_mem[98743] = 16'b0000000000000000;
	sram_mem[98744] = 16'b0000000000000000;
	sram_mem[98745] = 16'b0000000000000000;
	sram_mem[98746] = 16'b0000000000000000;
	sram_mem[98747] = 16'b0000000000000000;
	sram_mem[98748] = 16'b0000000000000000;
	sram_mem[98749] = 16'b0000000000000000;
	sram_mem[98750] = 16'b0000000000000000;
	sram_mem[98751] = 16'b0000000000000000;
	sram_mem[98752] = 16'b0000000000000000;
	sram_mem[98753] = 16'b0000000000000000;
	sram_mem[98754] = 16'b0000000000000000;
	sram_mem[98755] = 16'b0000000000000000;
	sram_mem[98756] = 16'b0000000000000000;
	sram_mem[98757] = 16'b0000000000000000;
	sram_mem[98758] = 16'b0000000000000000;
	sram_mem[98759] = 16'b0000000000000000;
	sram_mem[98760] = 16'b0000000000000000;
	sram_mem[98761] = 16'b0000000000000000;
	sram_mem[98762] = 16'b0000000000000000;
	sram_mem[98763] = 16'b0000000000000000;
	sram_mem[98764] = 16'b0000000000000000;
	sram_mem[98765] = 16'b0000000000000000;
	sram_mem[98766] = 16'b0000000000000000;
	sram_mem[98767] = 16'b0000000000000000;
	sram_mem[98768] = 16'b0000000000000000;
	sram_mem[98769] = 16'b0000000000000000;
	sram_mem[98770] = 16'b0000000000000000;
	sram_mem[98771] = 16'b0000000000000000;
	sram_mem[98772] = 16'b0000000000000000;
	sram_mem[98773] = 16'b0000000000000000;
	sram_mem[98774] = 16'b0000000000000000;
	sram_mem[98775] = 16'b0000000000000000;
	sram_mem[98776] = 16'b0000000000000000;
	sram_mem[98777] = 16'b0000000000000000;
	sram_mem[98778] = 16'b0000000000000000;
	sram_mem[98779] = 16'b0000000000000000;
	sram_mem[98780] = 16'b0000000000000000;
	sram_mem[98781] = 16'b0000000000000000;
	sram_mem[98782] = 16'b0000000000000000;
	sram_mem[98783] = 16'b0000000000000000;
	sram_mem[98784] = 16'b0000000000000000;
	sram_mem[98785] = 16'b0000000000000000;
	sram_mem[98786] = 16'b0000000000000000;
	sram_mem[98787] = 16'b0000000000000000;
	sram_mem[98788] = 16'b0000000000000000;
	sram_mem[98789] = 16'b0000000000000000;
	sram_mem[98790] = 16'b0000000000000000;
	sram_mem[98791] = 16'b0000000000000000;
	sram_mem[98792] = 16'b0000000000000000;
	sram_mem[98793] = 16'b0000000000000000;
	sram_mem[98794] = 16'b0000000000000000;
	sram_mem[98795] = 16'b0000000000000000;
	sram_mem[98796] = 16'b0000000000000000;
	sram_mem[98797] = 16'b0000000000000000;
	sram_mem[98798] = 16'b0000000000000000;
	sram_mem[98799] = 16'b0000000000000000;
	sram_mem[98800] = 16'b0000000000000000;
	sram_mem[98801] = 16'b0000000000000000;
	sram_mem[98802] = 16'b0000000000000000;
	sram_mem[98803] = 16'b0000000000000000;
	sram_mem[98804] = 16'b0000000000000000;
	sram_mem[98805] = 16'b0000000000000000;
	sram_mem[98806] = 16'b0000000000000000;
	sram_mem[98807] = 16'b0000000000000000;
	sram_mem[98808] = 16'b0000000000000000;
	sram_mem[98809] = 16'b0000000000000000;
	sram_mem[98810] = 16'b0000000000000000;
	sram_mem[98811] = 16'b0000000000000000;
	sram_mem[98812] = 16'b0000000000000000;
	sram_mem[98813] = 16'b0000000000000000;
	sram_mem[98814] = 16'b0000000000000000;
	sram_mem[98815] = 16'b0000000000000000;
	sram_mem[98816] = 16'b0000000000000000;
	sram_mem[98817] = 16'b0000000000000000;
	sram_mem[98818] = 16'b0000000000000000;
	sram_mem[98819] = 16'b0000000000000000;
	sram_mem[98820] = 16'b0000000000000000;
	sram_mem[98821] = 16'b0000000000000000;
	sram_mem[98822] = 16'b0000000000000000;
	sram_mem[98823] = 16'b0000000000000000;
	sram_mem[98824] = 16'b0000000000000000;
	sram_mem[98825] = 16'b0000000000000000;
	sram_mem[98826] = 16'b0000000000000000;
	sram_mem[98827] = 16'b0000000000000000;
	sram_mem[98828] = 16'b0000000000000000;
	sram_mem[98829] = 16'b0000000000000000;
	sram_mem[98830] = 16'b0000000000000000;
	sram_mem[98831] = 16'b0000000000000000;
	sram_mem[98832] = 16'b0000000000000000;
	sram_mem[98833] = 16'b0000000000000000;
	sram_mem[98834] = 16'b0000000000000000;
	sram_mem[98835] = 16'b0000000000000000;
	sram_mem[98836] = 16'b0000000000000000;
	sram_mem[98837] = 16'b0000000000000000;
	sram_mem[98838] = 16'b0000000000000000;
	sram_mem[98839] = 16'b0000000000000000;
	sram_mem[98840] = 16'b0000000000000000;
	sram_mem[98841] = 16'b0000000000000000;
	sram_mem[98842] = 16'b0000000000000000;
	sram_mem[98843] = 16'b0000000000000000;
	sram_mem[98844] = 16'b0000000000000000;
	sram_mem[98845] = 16'b0000000000000000;
	sram_mem[98846] = 16'b0000000000000000;
	sram_mem[98847] = 16'b0000000000000000;
	sram_mem[98848] = 16'b0000000000000000;
	sram_mem[98849] = 16'b0000000000000000;
	sram_mem[98850] = 16'b0000000000000000;
	sram_mem[98851] = 16'b0000000000000000;
	sram_mem[98852] = 16'b0000000000000000;
	sram_mem[98853] = 16'b0000000000000000;
	sram_mem[98854] = 16'b0000000000000000;
	sram_mem[98855] = 16'b0000000000000000;
	sram_mem[98856] = 16'b0000000000000000;
	sram_mem[98857] = 16'b0000000000000000;
	sram_mem[98858] = 16'b0000000000000000;
	sram_mem[98859] = 16'b0000000000000000;
	sram_mem[98860] = 16'b0000000000000000;
	sram_mem[98861] = 16'b0000000000000000;
	sram_mem[98862] = 16'b0000000000000000;
	sram_mem[98863] = 16'b0000000000000000;
	sram_mem[98864] = 16'b0000000000000000;
	sram_mem[98865] = 16'b0000000000000000;
	sram_mem[98866] = 16'b0000000000000000;
	sram_mem[98867] = 16'b0000000000000000;
	sram_mem[98868] = 16'b0000000000000000;
	sram_mem[98869] = 16'b0000000000000000;
	sram_mem[98870] = 16'b0000000000000000;
	sram_mem[98871] = 16'b0000000000000000;
	sram_mem[98872] = 16'b0000000000000000;
	sram_mem[98873] = 16'b0000000000000000;
	sram_mem[98874] = 16'b0000000000000000;
	sram_mem[98875] = 16'b0000000000000000;
	sram_mem[98876] = 16'b0000000000000000;
	sram_mem[98877] = 16'b0000000000000000;
	sram_mem[98878] = 16'b0000000000000000;
	sram_mem[98879] = 16'b0000000000000000;
	sram_mem[98880] = 16'b0000000000000000;
	sram_mem[98881] = 16'b0000000000000000;
	sram_mem[98882] = 16'b0000000000000000;
	sram_mem[98883] = 16'b0000000000000000;
	sram_mem[98884] = 16'b0000000000000000;
	sram_mem[98885] = 16'b0000000000000000;
	sram_mem[98886] = 16'b0000000000000000;
	sram_mem[98887] = 16'b0000000000000000;
	sram_mem[98888] = 16'b0000000000000000;
	sram_mem[98889] = 16'b0000000000000000;
	sram_mem[98890] = 16'b0000000000000000;
	sram_mem[98891] = 16'b0000000000000000;
	sram_mem[98892] = 16'b0000000000000000;
	sram_mem[98893] = 16'b0000000000000000;
	sram_mem[98894] = 16'b0000000000000000;
	sram_mem[98895] = 16'b0000000000000000;
	sram_mem[98896] = 16'b0000000000000000;
	sram_mem[98897] = 16'b0000000000000000;
	sram_mem[98898] = 16'b0000000000000000;
	sram_mem[98899] = 16'b0000000000000000;
	sram_mem[98900] = 16'b0000000000000000;
	sram_mem[98901] = 16'b0000000000000000;
	sram_mem[98902] = 16'b0000000000000000;
	sram_mem[98903] = 16'b0000000000000000;
	sram_mem[98904] = 16'b0000000000000000;
	sram_mem[98905] = 16'b0000000000000000;
	sram_mem[98906] = 16'b0000000000000000;
	sram_mem[98907] = 16'b0000000000000000;
	sram_mem[98908] = 16'b0000000000000000;
	sram_mem[98909] = 16'b0000000000000000;
	sram_mem[98910] = 16'b0000000000000000;
	sram_mem[98911] = 16'b0000000000000000;
	sram_mem[98912] = 16'b0000000000000000;
	sram_mem[98913] = 16'b0000000000000000;
	sram_mem[98914] = 16'b0000000000000000;
	sram_mem[98915] = 16'b0000000000000000;
	sram_mem[98916] = 16'b0000000000000000;
	sram_mem[98917] = 16'b0000000000000000;
	sram_mem[98918] = 16'b0000000000000000;
	sram_mem[98919] = 16'b0000000000000000;
	sram_mem[98920] = 16'b0000000000000000;
	sram_mem[98921] = 16'b0000000000000000;
	sram_mem[98922] = 16'b0000000000000000;
	sram_mem[98923] = 16'b0000000000000000;
	sram_mem[98924] = 16'b0000000000000000;
	sram_mem[98925] = 16'b0000000000000000;
	sram_mem[98926] = 16'b0000000000000000;
	sram_mem[98927] = 16'b0000000000000000;
	sram_mem[98928] = 16'b0000000000000000;
	sram_mem[98929] = 16'b0000000000000000;
	sram_mem[98930] = 16'b0000000000000000;
	sram_mem[98931] = 16'b0000000000000000;
	sram_mem[98932] = 16'b0000000000000000;
	sram_mem[98933] = 16'b0000000000000000;
	sram_mem[98934] = 16'b0000000000000000;
	sram_mem[98935] = 16'b0000000000000000;
	sram_mem[98936] = 16'b0000000000000000;
	sram_mem[98937] = 16'b0000000000000000;
	sram_mem[98938] = 16'b0000000000000000;
	sram_mem[98939] = 16'b0000000000000000;
	sram_mem[98940] = 16'b0000000000000000;
	sram_mem[98941] = 16'b0000000000000000;
	sram_mem[98942] = 16'b0000000000000000;
	sram_mem[98943] = 16'b0000000000000000;
	sram_mem[98944] = 16'b0000000000000000;
	sram_mem[98945] = 16'b0000000000000000;
	sram_mem[98946] = 16'b0000000000000000;
	sram_mem[98947] = 16'b0000000000000000;
	sram_mem[98948] = 16'b0000000000000000;
	sram_mem[98949] = 16'b0000000000000000;
	sram_mem[98950] = 16'b0000000000000000;
	sram_mem[98951] = 16'b0000000000000000;
	sram_mem[98952] = 16'b0000000000000000;
	sram_mem[98953] = 16'b0000000000000000;
	sram_mem[98954] = 16'b0000000000000000;
	sram_mem[98955] = 16'b0000000000000000;
	sram_mem[98956] = 16'b0000000000000000;
	sram_mem[98957] = 16'b0000000000000000;
	sram_mem[98958] = 16'b0000000000000000;
	sram_mem[98959] = 16'b0000000000000000;
	sram_mem[98960] = 16'b0000000000000000;
	sram_mem[98961] = 16'b0000000000000000;
	sram_mem[98962] = 16'b0000000000000000;
	sram_mem[98963] = 16'b0000000000000000;
	sram_mem[98964] = 16'b0000000000000000;
	sram_mem[98965] = 16'b0000000000000000;
	sram_mem[98966] = 16'b0000000000000000;
	sram_mem[98967] = 16'b0000000000000000;
	sram_mem[98968] = 16'b0000000000000000;
	sram_mem[98969] = 16'b0000000000000000;
	sram_mem[98970] = 16'b0000000000000000;
	sram_mem[98971] = 16'b0000000000000000;
	sram_mem[98972] = 16'b0000000000000000;
	sram_mem[98973] = 16'b0000000000000000;
	sram_mem[98974] = 16'b0000000000000000;
	sram_mem[98975] = 16'b0000000000000000;
	sram_mem[98976] = 16'b0000000000000000;
	sram_mem[98977] = 16'b0000000000000000;
	sram_mem[98978] = 16'b0000000000000000;
	sram_mem[98979] = 16'b0000000000000000;
	sram_mem[98980] = 16'b0000000000000000;
	sram_mem[98981] = 16'b0000000000000000;
	sram_mem[98982] = 16'b0000000000000000;
	sram_mem[98983] = 16'b0000000000000000;
	sram_mem[98984] = 16'b0000000000000000;
	sram_mem[98985] = 16'b0000000000000000;
	sram_mem[98986] = 16'b0000000000000000;
	sram_mem[98987] = 16'b0000000000000000;
	sram_mem[98988] = 16'b0000000000000000;
	sram_mem[98989] = 16'b0000000000000000;
	sram_mem[98990] = 16'b0000000000000000;
	sram_mem[98991] = 16'b0000000000000000;
	sram_mem[98992] = 16'b0000000000000000;
	sram_mem[98993] = 16'b0000000000000000;
	sram_mem[98994] = 16'b0000000000000000;
	sram_mem[98995] = 16'b0000000000000000;
	sram_mem[98996] = 16'b0000000000000000;
	sram_mem[98997] = 16'b0000000000000000;
	sram_mem[98998] = 16'b0000000000000000;
	sram_mem[98999] = 16'b0000000000000000;
	sram_mem[99000] = 16'b0000000000000000;
	sram_mem[99001] = 16'b0000000000000000;
	sram_mem[99002] = 16'b0000000000000000;
	sram_mem[99003] = 16'b0000000000000000;
	sram_mem[99004] = 16'b0000000000000000;
	sram_mem[99005] = 16'b0000000000000000;
	sram_mem[99006] = 16'b0000000000000000;
	sram_mem[99007] = 16'b0000000000000000;
	sram_mem[99008] = 16'b0000000000000000;
	sram_mem[99009] = 16'b0000000000000000;
	sram_mem[99010] = 16'b0000000000000000;
	sram_mem[99011] = 16'b0000000000000000;
	sram_mem[99012] = 16'b0000000000000000;
	sram_mem[99013] = 16'b0000000000000000;
	sram_mem[99014] = 16'b0000000000000000;
	sram_mem[99015] = 16'b0000000000000000;
	sram_mem[99016] = 16'b0000000000000000;
	sram_mem[99017] = 16'b0000000000000000;
	sram_mem[99018] = 16'b0000000000000000;
	sram_mem[99019] = 16'b0000000000000000;
	sram_mem[99020] = 16'b0000000000000000;
	sram_mem[99021] = 16'b0000000000000000;
	sram_mem[99022] = 16'b0000000000000000;
	sram_mem[99023] = 16'b0000000000000000;
	sram_mem[99024] = 16'b0000000000000000;
	sram_mem[99025] = 16'b0000000000000000;
	sram_mem[99026] = 16'b0000000000000000;
	sram_mem[99027] = 16'b0000000000000000;
	sram_mem[99028] = 16'b0000000000000000;
	sram_mem[99029] = 16'b0000000000000000;
	sram_mem[99030] = 16'b0000000000000000;
	sram_mem[99031] = 16'b0000000000000000;
	sram_mem[99032] = 16'b0000000000000000;
	sram_mem[99033] = 16'b0000000000000000;
	sram_mem[99034] = 16'b0000000000000000;
	sram_mem[99035] = 16'b0000000000000000;
	sram_mem[99036] = 16'b0000000000000000;
	sram_mem[99037] = 16'b0000000000000000;
	sram_mem[99038] = 16'b0000000000000000;
	sram_mem[99039] = 16'b0000000000000000;
	sram_mem[99040] = 16'b0000000000000000;
	sram_mem[99041] = 16'b0000000000000000;
	sram_mem[99042] = 16'b0000000000000000;
	sram_mem[99043] = 16'b0000000000000000;
	sram_mem[99044] = 16'b0000000000000000;
	sram_mem[99045] = 16'b0000000000000000;
	sram_mem[99046] = 16'b0000000000000000;
	sram_mem[99047] = 16'b0000000000000000;
	sram_mem[99048] = 16'b0000000000000000;
	sram_mem[99049] = 16'b0000000000000000;
	sram_mem[99050] = 16'b0000000000000000;
	sram_mem[99051] = 16'b0000000000000000;
	sram_mem[99052] = 16'b0000000000000000;
	sram_mem[99053] = 16'b0000000000000000;
	sram_mem[99054] = 16'b0000000000000000;
	sram_mem[99055] = 16'b0000000000000000;
	sram_mem[99056] = 16'b0000000000000000;
	sram_mem[99057] = 16'b0000000000000000;
	sram_mem[99058] = 16'b0000000000000000;
	sram_mem[99059] = 16'b0000000000000000;
	sram_mem[99060] = 16'b0000000000000000;
	sram_mem[99061] = 16'b0000000000000000;
	sram_mem[99062] = 16'b0000000000000000;
	sram_mem[99063] = 16'b0000000000000000;
	sram_mem[99064] = 16'b0000000000000000;
	sram_mem[99065] = 16'b0000000000000000;
	sram_mem[99066] = 16'b0000000000000000;
	sram_mem[99067] = 16'b0000000000000000;
	sram_mem[99068] = 16'b0000000000000000;
	sram_mem[99069] = 16'b0000000000000000;
	sram_mem[99070] = 16'b0000000000000000;
	sram_mem[99071] = 16'b0000000000000000;
	sram_mem[99072] = 16'b0000000000000000;
	sram_mem[99073] = 16'b0000000000000000;
	sram_mem[99074] = 16'b0000000000000000;
	sram_mem[99075] = 16'b0000000000000000;
	sram_mem[99076] = 16'b0000000000000000;
	sram_mem[99077] = 16'b0000000000000000;
	sram_mem[99078] = 16'b0000000000000000;
	sram_mem[99079] = 16'b0000000000000000;
	sram_mem[99080] = 16'b0000000000000000;
	sram_mem[99081] = 16'b0000000000000000;
	sram_mem[99082] = 16'b0000000000000000;
	sram_mem[99083] = 16'b0000000000000000;
	sram_mem[99084] = 16'b0000000000000000;
	sram_mem[99085] = 16'b0000000000000000;
	sram_mem[99086] = 16'b0000000000000000;
	sram_mem[99087] = 16'b0000000000000000;
	sram_mem[99088] = 16'b0000000000000000;
	sram_mem[99089] = 16'b0000000000000000;
	sram_mem[99090] = 16'b0000000000000000;
	sram_mem[99091] = 16'b0000000000000000;
	sram_mem[99092] = 16'b0000000000000000;
	sram_mem[99093] = 16'b0000000000000000;
	sram_mem[99094] = 16'b0000000000000000;
	sram_mem[99095] = 16'b0000000000000000;
	sram_mem[99096] = 16'b0000000000000000;
	sram_mem[99097] = 16'b0000000000000000;
	sram_mem[99098] = 16'b0000000000000000;
	sram_mem[99099] = 16'b0000000000000000;
	sram_mem[99100] = 16'b0000000000000000;
	sram_mem[99101] = 16'b0000000000000000;
	sram_mem[99102] = 16'b0000000000000000;
	sram_mem[99103] = 16'b0000000000000000;
	sram_mem[99104] = 16'b0000000000000000;
	sram_mem[99105] = 16'b0000000000000000;
	sram_mem[99106] = 16'b0000000000000000;
	sram_mem[99107] = 16'b0000000000000000;
	sram_mem[99108] = 16'b0000000000000000;
	sram_mem[99109] = 16'b0000000000000000;
	sram_mem[99110] = 16'b0000000000000000;
	sram_mem[99111] = 16'b0000000000000000;
	sram_mem[99112] = 16'b0000000000000000;
	sram_mem[99113] = 16'b0000000000000000;
	sram_mem[99114] = 16'b0000000000000000;
	sram_mem[99115] = 16'b0000000000000000;
	sram_mem[99116] = 16'b0000000000000000;
	sram_mem[99117] = 16'b0000000000000000;
	sram_mem[99118] = 16'b0000000000000000;
	sram_mem[99119] = 16'b0000000000000000;
	sram_mem[99120] = 16'b0000000000000000;
	sram_mem[99121] = 16'b0000000000000000;
	sram_mem[99122] = 16'b0000000000000000;
	sram_mem[99123] = 16'b0000000000000000;
	sram_mem[99124] = 16'b0000000000000000;
	sram_mem[99125] = 16'b0000000000000000;
	sram_mem[99126] = 16'b0000000000000000;
	sram_mem[99127] = 16'b0000000000000000;
	sram_mem[99128] = 16'b0000000000000000;
	sram_mem[99129] = 16'b0000000000000000;
	sram_mem[99130] = 16'b0000000000000000;
	sram_mem[99131] = 16'b0000000000000000;
	sram_mem[99132] = 16'b0000000000000000;
	sram_mem[99133] = 16'b0000000000000000;
	sram_mem[99134] = 16'b0000000000000000;
	sram_mem[99135] = 16'b0000000000000000;
	sram_mem[99136] = 16'b0000000000000000;
	sram_mem[99137] = 16'b0000000000000000;
	sram_mem[99138] = 16'b0000000000000000;
	sram_mem[99139] = 16'b0000000000000000;
	sram_mem[99140] = 16'b0000000000000000;
	sram_mem[99141] = 16'b0000000000000000;
	sram_mem[99142] = 16'b0000000000000000;
	sram_mem[99143] = 16'b0000000000000000;
	sram_mem[99144] = 16'b0000000000000000;
	sram_mem[99145] = 16'b0000000000000000;
	sram_mem[99146] = 16'b0000000000000000;
	sram_mem[99147] = 16'b0000000000000000;
	sram_mem[99148] = 16'b0000000000000000;
	sram_mem[99149] = 16'b0000000000000000;
	sram_mem[99150] = 16'b0000000000000000;
	sram_mem[99151] = 16'b0000000000000000;
	sram_mem[99152] = 16'b0000000000000000;
	sram_mem[99153] = 16'b0000000000000000;
	sram_mem[99154] = 16'b0000000000000000;
	sram_mem[99155] = 16'b0000000000000000;
	sram_mem[99156] = 16'b0000000000000000;
	sram_mem[99157] = 16'b0000000000000000;
	sram_mem[99158] = 16'b0000000000000000;
	sram_mem[99159] = 16'b0000000000000000;
	sram_mem[99160] = 16'b0000000000000000;
	sram_mem[99161] = 16'b0000000000000000;
	sram_mem[99162] = 16'b0000000000000000;
	sram_mem[99163] = 16'b0000000000000000;
	sram_mem[99164] = 16'b0000000000000000;
	sram_mem[99165] = 16'b0000000000000000;
	sram_mem[99166] = 16'b0000000000000000;
	sram_mem[99167] = 16'b0000000000000000;
	sram_mem[99168] = 16'b0000000000000000;
	sram_mem[99169] = 16'b0000000000000000;
	sram_mem[99170] = 16'b0000000000000000;
	sram_mem[99171] = 16'b0000000000000000;
	sram_mem[99172] = 16'b0000000000000000;
	sram_mem[99173] = 16'b0000000000000000;
	sram_mem[99174] = 16'b0000000000000000;
	sram_mem[99175] = 16'b0000000000000000;
	sram_mem[99176] = 16'b0000000000000000;
	sram_mem[99177] = 16'b0000000000000000;
	sram_mem[99178] = 16'b0000000000000000;
	sram_mem[99179] = 16'b0000000000000000;
	sram_mem[99180] = 16'b0000000000000000;
	sram_mem[99181] = 16'b0000000000000000;
	sram_mem[99182] = 16'b0000000000000000;
	sram_mem[99183] = 16'b0000000000000000;
	sram_mem[99184] = 16'b0000000000000000;
	sram_mem[99185] = 16'b0000000000000000;
	sram_mem[99186] = 16'b0000000000000000;
	sram_mem[99187] = 16'b0000000000000000;
	sram_mem[99188] = 16'b0000000000000000;
	sram_mem[99189] = 16'b0000000000000000;
	sram_mem[99190] = 16'b0000000000000000;
	sram_mem[99191] = 16'b0000000000000000;
	sram_mem[99192] = 16'b0000000000000000;
	sram_mem[99193] = 16'b0000000000000000;
	sram_mem[99194] = 16'b0000000000000000;
	sram_mem[99195] = 16'b0000000000000000;
	sram_mem[99196] = 16'b0000000000000000;
	sram_mem[99197] = 16'b0000000000000000;
	sram_mem[99198] = 16'b0000000000000000;
	sram_mem[99199] = 16'b0000000000000000;
	sram_mem[99200] = 16'b0000000000000000;
	sram_mem[99201] = 16'b0000000000000000;
	sram_mem[99202] = 16'b0000000000000000;
	sram_mem[99203] = 16'b0000000000000000;
	sram_mem[99204] = 16'b0000000000000000;
	sram_mem[99205] = 16'b0000000000000000;
	sram_mem[99206] = 16'b0000000000000000;
	sram_mem[99207] = 16'b0000000000000000;
	sram_mem[99208] = 16'b0000000000000000;
	sram_mem[99209] = 16'b0000000000000000;
	sram_mem[99210] = 16'b0000000000000000;
	sram_mem[99211] = 16'b0000000000000000;
	sram_mem[99212] = 16'b0000000000000000;
	sram_mem[99213] = 16'b0000000000000000;
	sram_mem[99214] = 16'b0000000000000000;
	sram_mem[99215] = 16'b0000000000000000;
	sram_mem[99216] = 16'b0000000000000000;
	sram_mem[99217] = 16'b0000000000000000;
	sram_mem[99218] = 16'b0000000000000000;
	sram_mem[99219] = 16'b0000000000000000;
	sram_mem[99220] = 16'b0000000000000000;
	sram_mem[99221] = 16'b0000000000000000;
	sram_mem[99222] = 16'b0000000000000000;
	sram_mem[99223] = 16'b0000000000000000;
	sram_mem[99224] = 16'b0000000000000000;
	sram_mem[99225] = 16'b0000000000000000;
	sram_mem[99226] = 16'b0000000000000000;
	sram_mem[99227] = 16'b0000000000000000;
	sram_mem[99228] = 16'b0000000000000000;
	sram_mem[99229] = 16'b0000000000000000;
	sram_mem[99230] = 16'b0000000000000000;
	sram_mem[99231] = 16'b0000000000000000;
	sram_mem[99232] = 16'b0000000000000000;
	sram_mem[99233] = 16'b0000000000000000;
	sram_mem[99234] = 16'b0000000000000000;
	sram_mem[99235] = 16'b0000000000000000;
	sram_mem[99236] = 16'b0000000000000000;
	sram_mem[99237] = 16'b0000000000000000;
	sram_mem[99238] = 16'b0000000000000000;
	sram_mem[99239] = 16'b0000000000000000;
	sram_mem[99240] = 16'b0000000000000000;
	sram_mem[99241] = 16'b0000000000000000;
	sram_mem[99242] = 16'b0000000000000000;
	sram_mem[99243] = 16'b0000000000000000;
	sram_mem[99244] = 16'b0000000000000000;
	sram_mem[99245] = 16'b0000000000000000;
	sram_mem[99246] = 16'b0000000000000000;
	sram_mem[99247] = 16'b0000000000000000;
	sram_mem[99248] = 16'b0000000000000000;
	sram_mem[99249] = 16'b0000000000000000;
	sram_mem[99250] = 16'b0000000000000000;
	sram_mem[99251] = 16'b0000000000000000;
	sram_mem[99252] = 16'b0000000000000000;
	sram_mem[99253] = 16'b0000000000000000;
	sram_mem[99254] = 16'b0000000000000000;
	sram_mem[99255] = 16'b0000000000000000;
	sram_mem[99256] = 16'b0000000000000000;
	sram_mem[99257] = 16'b0000000000000000;
	sram_mem[99258] = 16'b0000000000000000;
	sram_mem[99259] = 16'b0000000000000000;
	sram_mem[99260] = 16'b0000000000000000;
	sram_mem[99261] = 16'b0000000000000000;
	sram_mem[99262] = 16'b0000000000000000;
	sram_mem[99263] = 16'b0000000000000000;
	sram_mem[99264] = 16'b0000000000000000;
	sram_mem[99265] = 16'b0000000000000000;
	sram_mem[99266] = 16'b0000000000000000;
	sram_mem[99267] = 16'b0000000000000000;
	sram_mem[99268] = 16'b0000000000000000;
	sram_mem[99269] = 16'b0000000000000000;
	sram_mem[99270] = 16'b0000000000000000;
	sram_mem[99271] = 16'b0000000000000000;
	sram_mem[99272] = 16'b0000000000000000;
	sram_mem[99273] = 16'b0000000000000000;
	sram_mem[99274] = 16'b0000000000000000;
	sram_mem[99275] = 16'b0000000000000000;
	sram_mem[99276] = 16'b0000000000000000;
	sram_mem[99277] = 16'b0000000000000000;
	sram_mem[99278] = 16'b0000000000000000;
	sram_mem[99279] = 16'b0000000000000000;
	sram_mem[99280] = 16'b0000000000000000;
	sram_mem[99281] = 16'b0000000000000000;
	sram_mem[99282] = 16'b0000000000000000;
	sram_mem[99283] = 16'b0000000000000000;
	sram_mem[99284] = 16'b0000000000000000;
	sram_mem[99285] = 16'b0000000000000000;
	sram_mem[99286] = 16'b0000000000000000;
	sram_mem[99287] = 16'b0000000000000000;
	sram_mem[99288] = 16'b0000000000000000;
	sram_mem[99289] = 16'b0000000000000000;
	sram_mem[99290] = 16'b0000000000000000;
	sram_mem[99291] = 16'b0000000000000000;
	sram_mem[99292] = 16'b0000000000000000;
	sram_mem[99293] = 16'b0000000000000000;
	sram_mem[99294] = 16'b0000000000000000;
	sram_mem[99295] = 16'b0000000000000000;
	sram_mem[99296] = 16'b0000000000000000;
	sram_mem[99297] = 16'b0000000000000000;
	sram_mem[99298] = 16'b0000000000000000;
	sram_mem[99299] = 16'b0000000000000000;
	sram_mem[99300] = 16'b0000000000000000;
	sram_mem[99301] = 16'b0000000000000000;
	sram_mem[99302] = 16'b0000000000000000;
	sram_mem[99303] = 16'b0000000000000000;
	sram_mem[99304] = 16'b0000000000000000;
	sram_mem[99305] = 16'b0000000000000000;
	sram_mem[99306] = 16'b0000000000000000;
	sram_mem[99307] = 16'b0000000000000000;
	sram_mem[99308] = 16'b0000000000000000;
	sram_mem[99309] = 16'b0000000000000000;
	sram_mem[99310] = 16'b0000000000000000;
	sram_mem[99311] = 16'b0000000000000000;
	sram_mem[99312] = 16'b0000000000000000;
	sram_mem[99313] = 16'b0000000000000000;
	sram_mem[99314] = 16'b0000000000000000;
	sram_mem[99315] = 16'b0000000000000000;
	sram_mem[99316] = 16'b0000000000000000;
	sram_mem[99317] = 16'b0000000000000000;
	sram_mem[99318] = 16'b0000000000000000;
	sram_mem[99319] = 16'b0000000000000000;
	sram_mem[99320] = 16'b0000000000000000;
	sram_mem[99321] = 16'b0000000000000000;
	sram_mem[99322] = 16'b0000000000000000;
	sram_mem[99323] = 16'b0000000000000000;
	sram_mem[99324] = 16'b0000000000000000;
	sram_mem[99325] = 16'b0000000000000000;
	sram_mem[99326] = 16'b0000000000000000;
	sram_mem[99327] = 16'b0000000000000000;
	sram_mem[99328] = 16'b0000000000000000;
	sram_mem[99329] = 16'b0000000000000000;
	sram_mem[99330] = 16'b0000000000000000;
	sram_mem[99331] = 16'b0000000000000000;
	sram_mem[99332] = 16'b0000000000000000;
	sram_mem[99333] = 16'b0000000000000000;
	sram_mem[99334] = 16'b0000000000000000;
	sram_mem[99335] = 16'b0000000000000000;
	sram_mem[99336] = 16'b0000000000000000;
	sram_mem[99337] = 16'b0000000000000000;
	sram_mem[99338] = 16'b0000000000000000;
	sram_mem[99339] = 16'b0000000000000000;
	sram_mem[99340] = 16'b0000000000000000;
	sram_mem[99341] = 16'b0000000000000000;
	sram_mem[99342] = 16'b0000000000000000;
	sram_mem[99343] = 16'b0000000000000000;
	sram_mem[99344] = 16'b0000000000000000;
	sram_mem[99345] = 16'b0000000000000000;
	sram_mem[99346] = 16'b0000000000000000;
	sram_mem[99347] = 16'b0000000000000000;
	sram_mem[99348] = 16'b0000000000000000;
	sram_mem[99349] = 16'b0000000000000000;
	sram_mem[99350] = 16'b0000000000000000;
	sram_mem[99351] = 16'b0000000000000000;
	sram_mem[99352] = 16'b0000000000000000;
	sram_mem[99353] = 16'b0000000000000000;
	sram_mem[99354] = 16'b0000000000000000;
	sram_mem[99355] = 16'b0000000000000000;
	sram_mem[99356] = 16'b0000000000000000;
	sram_mem[99357] = 16'b0000000000000000;
	sram_mem[99358] = 16'b0000000000000000;
	sram_mem[99359] = 16'b0000000000000000;
	sram_mem[99360] = 16'b0000000000000000;
	sram_mem[99361] = 16'b0000000000000000;
	sram_mem[99362] = 16'b0000000000000000;
	sram_mem[99363] = 16'b0000000000000000;
	sram_mem[99364] = 16'b0000000000000000;
	sram_mem[99365] = 16'b0000000000000000;
	sram_mem[99366] = 16'b0000000000000000;
	sram_mem[99367] = 16'b0000000000000000;
	sram_mem[99368] = 16'b0000000000000000;
	sram_mem[99369] = 16'b0000000000000000;
	sram_mem[99370] = 16'b0000000000000000;
	sram_mem[99371] = 16'b0000000000000000;
	sram_mem[99372] = 16'b0000000000000000;
	sram_mem[99373] = 16'b0000000000000000;
	sram_mem[99374] = 16'b0000000000000000;
	sram_mem[99375] = 16'b0000000000000000;
	sram_mem[99376] = 16'b0000000000000000;
	sram_mem[99377] = 16'b0000000000000000;
	sram_mem[99378] = 16'b0000000000000000;
	sram_mem[99379] = 16'b0000000000000000;
	sram_mem[99380] = 16'b0000000000000000;
	sram_mem[99381] = 16'b0000000000000000;
	sram_mem[99382] = 16'b0000000000000000;
	sram_mem[99383] = 16'b0000000000000000;
	sram_mem[99384] = 16'b0000000000000000;
	sram_mem[99385] = 16'b0000000000000000;
	sram_mem[99386] = 16'b0000000000000000;
	sram_mem[99387] = 16'b0000000000000000;
	sram_mem[99388] = 16'b0000000000000000;
	sram_mem[99389] = 16'b0000000000000000;
	sram_mem[99390] = 16'b0000000000000000;
	sram_mem[99391] = 16'b0000000000000000;
	sram_mem[99392] = 16'b0000000000000000;
	sram_mem[99393] = 16'b0000000000000000;
	sram_mem[99394] = 16'b0000000000000000;
	sram_mem[99395] = 16'b0000000000000000;
	sram_mem[99396] = 16'b0000000000000000;
	sram_mem[99397] = 16'b0000000000000000;
	sram_mem[99398] = 16'b0000000000000000;
	sram_mem[99399] = 16'b0000000000000000;
	sram_mem[99400] = 16'b0000000000000000;
	sram_mem[99401] = 16'b0000000000000000;
	sram_mem[99402] = 16'b0000000000000000;
	sram_mem[99403] = 16'b0000000000000000;
	sram_mem[99404] = 16'b0000000000000000;
	sram_mem[99405] = 16'b0000000000000000;
	sram_mem[99406] = 16'b0000000000000000;
	sram_mem[99407] = 16'b0000000000000000;
	sram_mem[99408] = 16'b0000000000000000;
	sram_mem[99409] = 16'b0000000000000000;
	sram_mem[99410] = 16'b0000000000000000;
	sram_mem[99411] = 16'b0000000000000000;
	sram_mem[99412] = 16'b0000000000000000;
	sram_mem[99413] = 16'b0000000000000000;
	sram_mem[99414] = 16'b0000000000000000;
	sram_mem[99415] = 16'b0000000000000000;
	sram_mem[99416] = 16'b0000000000000000;
	sram_mem[99417] = 16'b0000000000000000;
	sram_mem[99418] = 16'b0000000000000000;
	sram_mem[99419] = 16'b0000000000000000;
	sram_mem[99420] = 16'b0000000000000000;
	sram_mem[99421] = 16'b0000000000000000;
	sram_mem[99422] = 16'b0000000000000000;
	sram_mem[99423] = 16'b0000000000000000;
	sram_mem[99424] = 16'b0000000000000000;
	sram_mem[99425] = 16'b0000000000000000;
	sram_mem[99426] = 16'b0000000000000000;
	sram_mem[99427] = 16'b0000000000000000;
	sram_mem[99428] = 16'b0000000000000000;
	sram_mem[99429] = 16'b0000000000000000;
	sram_mem[99430] = 16'b0000000000000000;
	sram_mem[99431] = 16'b0000000000000000;
	sram_mem[99432] = 16'b0000000000000000;
	sram_mem[99433] = 16'b0000000000000000;
	sram_mem[99434] = 16'b0000000000000000;
	sram_mem[99435] = 16'b0000000000000000;
	sram_mem[99436] = 16'b0000000000000000;
	sram_mem[99437] = 16'b0000000000000000;
	sram_mem[99438] = 16'b0000000000000000;
	sram_mem[99439] = 16'b0000000000000000;
	sram_mem[99440] = 16'b0000000000000000;
	sram_mem[99441] = 16'b0000000000000000;
	sram_mem[99442] = 16'b0000000000000000;
	sram_mem[99443] = 16'b0000000000000000;
	sram_mem[99444] = 16'b0000000000000000;
	sram_mem[99445] = 16'b0000000000000000;
	sram_mem[99446] = 16'b0000000000000000;
	sram_mem[99447] = 16'b0000000000000000;
	sram_mem[99448] = 16'b0000000000000000;
	sram_mem[99449] = 16'b0000000000000000;
	sram_mem[99450] = 16'b0000000000000000;
	sram_mem[99451] = 16'b0000000000000000;
	sram_mem[99452] = 16'b0000000000000000;
	sram_mem[99453] = 16'b0000000000000000;
	sram_mem[99454] = 16'b0000000000000000;
	sram_mem[99455] = 16'b0000000000000000;
	sram_mem[99456] = 16'b0000000000000000;
	sram_mem[99457] = 16'b0000000000000000;
	sram_mem[99458] = 16'b0000000000000000;
	sram_mem[99459] = 16'b0000000000000000;
	sram_mem[99460] = 16'b0000000000000000;
	sram_mem[99461] = 16'b0000000000000000;
	sram_mem[99462] = 16'b0000000000000000;
	sram_mem[99463] = 16'b0000000000000000;
	sram_mem[99464] = 16'b0000000000000000;
	sram_mem[99465] = 16'b0000000000000000;
	sram_mem[99466] = 16'b0000000000000000;
	sram_mem[99467] = 16'b0000000000000000;
	sram_mem[99468] = 16'b0000000000000000;
	sram_mem[99469] = 16'b0000000000000000;
	sram_mem[99470] = 16'b0000000000000000;
	sram_mem[99471] = 16'b0000000000000000;
	sram_mem[99472] = 16'b0000000000000000;
	sram_mem[99473] = 16'b0000000000000000;
	sram_mem[99474] = 16'b0000000000000000;
	sram_mem[99475] = 16'b0000000000000000;
	sram_mem[99476] = 16'b0000000000000000;
	sram_mem[99477] = 16'b0000000000000000;
	sram_mem[99478] = 16'b0000000000000000;
	sram_mem[99479] = 16'b0000000000000000;
	sram_mem[99480] = 16'b0000000000000000;
	sram_mem[99481] = 16'b0000000000000000;
	sram_mem[99482] = 16'b0000000000000000;
	sram_mem[99483] = 16'b0000000000000000;
	sram_mem[99484] = 16'b0000000000000000;
	sram_mem[99485] = 16'b0000000000000000;
	sram_mem[99486] = 16'b0000000000000000;
	sram_mem[99487] = 16'b0000000000000000;
	sram_mem[99488] = 16'b0000000000000000;
	sram_mem[99489] = 16'b0000000000000000;
	sram_mem[99490] = 16'b0000000000000000;
	sram_mem[99491] = 16'b0000000000000000;
	sram_mem[99492] = 16'b0000000000000000;
	sram_mem[99493] = 16'b0000000000000000;
	sram_mem[99494] = 16'b0000000000000000;
	sram_mem[99495] = 16'b0000000000000000;
	sram_mem[99496] = 16'b0000000000000000;
	sram_mem[99497] = 16'b0000000000000000;
	sram_mem[99498] = 16'b0000000000000000;
	sram_mem[99499] = 16'b0000000000000000;
	sram_mem[99500] = 16'b0000000000000000;
	sram_mem[99501] = 16'b0000000000000000;
	sram_mem[99502] = 16'b0000000000000000;
	sram_mem[99503] = 16'b0000000000000000;
	sram_mem[99504] = 16'b0000000000000000;
	sram_mem[99505] = 16'b0000000000000000;
	sram_mem[99506] = 16'b0000000000000000;
	sram_mem[99507] = 16'b0000000000000000;
	sram_mem[99508] = 16'b0000000000000000;
	sram_mem[99509] = 16'b0000000000000000;
	sram_mem[99510] = 16'b0000000000000000;
	sram_mem[99511] = 16'b0000000000000000;
	sram_mem[99512] = 16'b0000000000000000;
	sram_mem[99513] = 16'b0000000000000000;
	sram_mem[99514] = 16'b0000000000000000;
	sram_mem[99515] = 16'b0000000000000000;
	sram_mem[99516] = 16'b0000000000000000;
	sram_mem[99517] = 16'b0000000000000000;
	sram_mem[99518] = 16'b0000000000000000;
	sram_mem[99519] = 16'b0000000000000000;
	sram_mem[99520] = 16'b0000000000000000;
	sram_mem[99521] = 16'b0000000000000000;
	sram_mem[99522] = 16'b0000000000000000;
	sram_mem[99523] = 16'b0000000000000000;
	sram_mem[99524] = 16'b0000000000000000;
	sram_mem[99525] = 16'b0000000000000000;
	sram_mem[99526] = 16'b0000000000000000;
	sram_mem[99527] = 16'b0000000000000000;
	sram_mem[99528] = 16'b0000000000000000;
	sram_mem[99529] = 16'b0000000000000000;
	sram_mem[99530] = 16'b0000000000000000;
	sram_mem[99531] = 16'b0000000000000000;
	sram_mem[99532] = 16'b0000000000000000;
	sram_mem[99533] = 16'b0000000000000000;
	sram_mem[99534] = 16'b0000000000000000;
	sram_mem[99535] = 16'b0000000000000000;
	sram_mem[99536] = 16'b0000000000000000;
	sram_mem[99537] = 16'b0000000000000000;
	sram_mem[99538] = 16'b0000000000000000;
	sram_mem[99539] = 16'b0000000000000000;
	sram_mem[99540] = 16'b0000000000000000;
	sram_mem[99541] = 16'b0000000000000000;
	sram_mem[99542] = 16'b0000000000000000;
	sram_mem[99543] = 16'b0000000000000000;
	sram_mem[99544] = 16'b0000000000000000;
	sram_mem[99545] = 16'b0000000000000000;
	sram_mem[99546] = 16'b0000000000000000;
	sram_mem[99547] = 16'b0000000000000000;
	sram_mem[99548] = 16'b0000000000000000;
	sram_mem[99549] = 16'b0000000000000000;
	sram_mem[99550] = 16'b0000000000000000;
	sram_mem[99551] = 16'b0000000000000000;
	sram_mem[99552] = 16'b0000000000000000;
	sram_mem[99553] = 16'b0000000000000000;
	sram_mem[99554] = 16'b0000000000000000;
	sram_mem[99555] = 16'b0000000000000000;
	sram_mem[99556] = 16'b0000000000000000;
	sram_mem[99557] = 16'b0000000000000000;
	sram_mem[99558] = 16'b0000000000000000;
	sram_mem[99559] = 16'b0000000000000000;
	sram_mem[99560] = 16'b0000000000000000;
	sram_mem[99561] = 16'b0000000000000000;
	sram_mem[99562] = 16'b0000000000000000;
	sram_mem[99563] = 16'b0000000000000000;
	sram_mem[99564] = 16'b0000000000000000;
	sram_mem[99565] = 16'b0000000000000000;
	sram_mem[99566] = 16'b0000000000000000;
	sram_mem[99567] = 16'b0000000000000000;
	sram_mem[99568] = 16'b0000000000000000;
	sram_mem[99569] = 16'b0000000000000000;
	sram_mem[99570] = 16'b0000000000000000;
	sram_mem[99571] = 16'b0000000000000000;
	sram_mem[99572] = 16'b0000000000000000;
	sram_mem[99573] = 16'b0000000000000000;
	sram_mem[99574] = 16'b0000000000000000;
	sram_mem[99575] = 16'b0000000000000000;
	sram_mem[99576] = 16'b0000000000000000;
	sram_mem[99577] = 16'b0000000000000000;
	sram_mem[99578] = 16'b0000000000000000;
	sram_mem[99579] = 16'b0000000000000000;
	sram_mem[99580] = 16'b0000000000000000;
	sram_mem[99581] = 16'b0000000000000000;
	sram_mem[99582] = 16'b0000000000000000;
	sram_mem[99583] = 16'b0000000000000000;
	sram_mem[99584] = 16'b0000000000000000;
	sram_mem[99585] = 16'b0000000000000000;
	sram_mem[99586] = 16'b0000000000000000;
	sram_mem[99587] = 16'b0000000000000000;
	sram_mem[99588] = 16'b0000000000000000;
	sram_mem[99589] = 16'b0000000000000000;
	sram_mem[99590] = 16'b0000000000000000;
	sram_mem[99591] = 16'b0000000000000000;
	sram_mem[99592] = 16'b0000000000000000;
	sram_mem[99593] = 16'b0000000000000000;
	sram_mem[99594] = 16'b0000000000000000;
	sram_mem[99595] = 16'b0000000000000000;
	sram_mem[99596] = 16'b0000000000000000;
	sram_mem[99597] = 16'b0000000000000000;
	sram_mem[99598] = 16'b0000000000000000;
	sram_mem[99599] = 16'b0000000000000000;
	sram_mem[99600] = 16'b0000000000000000;
	sram_mem[99601] = 16'b0000000000000000;
	sram_mem[99602] = 16'b0000000000000000;
	sram_mem[99603] = 16'b0000000000000000;
	sram_mem[99604] = 16'b0000000000000000;
	sram_mem[99605] = 16'b0000000000000000;
	sram_mem[99606] = 16'b0000000000000000;
	sram_mem[99607] = 16'b0000000000000000;
	sram_mem[99608] = 16'b0000000000000000;
	sram_mem[99609] = 16'b0000000000000000;
	sram_mem[99610] = 16'b0000000000000000;
	sram_mem[99611] = 16'b0000000000000000;
	sram_mem[99612] = 16'b0000000000000000;
	sram_mem[99613] = 16'b0000000000000000;
	sram_mem[99614] = 16'b0000000000000000;
	sram_mem[99615] = 16'b0000000000000000;
	sram_mem[99616] = 16'b0000000000000000;
	sram_mem[99617] = 16'b0000000000000000;
	sram_mem[99618] = 16'b0000000000000000;
	sram_mem[99619] = 16'b0000000000000000;
	sram_mem[99620] = 16'b0000000000000000;
	sram_mem[99621] = 16'b0000000000000000;
	sram_mem[99622] = 16'b0000000000000000;
	sram_mem[99623] = 16'b0000000000000000;
	sram_mem[99624] = 16'b0000000000000000;
	sram_mem[99625] = 16'b0000000000000000;
	sram_mem[99626] = 16'b0000000000000000;
	sram_mem[99627] = 16'b0000000000000000;
	sram_mem[99628] = 16'b0000000000000000;
	sram_mem[99629] = 16'b0000000000000000;
	sram_mem[99630] = 16'b0000000000000000;
	sram_mem[99631] = 16'b0000000000000000;
	sram_mem[99632] = 16'b0000000000000000;
	sram_mem[99633] = 16'b0000000000000000;
	sram_mem[99634] = 16'b0000000000000000;
	sram_mem[99635] = 16'b0000000000000000;
	sram_mem[99636] = 16'b0000000000000000;
	sram_mem[99637] = 16'b0000000000000000;
	sram_mem[99638] = 16'b0000000000000000;
	sram_mem[99639] = 16'b0000000000000000;
	sram_mem[99640] = 16'b0000000000000000;
	sram_mem[99641] = 16'b0000000000000000;
	sram_mem[99642] = 16'b0000000000000000;
	sram_mem[99643] = 16'b0000000000000000;
	sram_mem[99644] = 16'b0000000000000000;
	sram_mem[99645] = 16'b0000000000000000;
	sram_mem[99646] = 16'b0000000000000000;
	sram_mem[99647] = 16'b0000000000000000;
	sram_mem[99648] = 16'b0000000000000000;
	sram_mem[99649] = 16'b0000000000000000;
	sram_mem[99650] = 16'b0000000000000000;
	sram_mem[99651] = 16'b0000000000000000;
	sram_mem[99652] = 16'b0000000000000000;
	sram_mem[99653] = 16'b0000000000000000;
	sram_mem[99654] = 16'b0000000000000000;
	sram_mem[99655] = 16'b0000000000000000;
	sram_mem[99656] = 16'b0000000000000000;
	sram_mem[99657] = 16'b0000000000000000;
	sram_mem[99658] = 16'b0000000000000000;
	sram_mem[99659] = 16'b0000000000000000;
	sram_mem[99660] = 16'b0000000000000000;
	sram_mem[99661] = 16'b0000000000000000;
	sram_mem[99662] = 16'b0000000000000000;
	sram_mem[99663] = 16'b0000000000000000;
	sram_mem[99664] = 16'b0000000000000000;
	sram_mem[99665] = 16'b0000000000000000;
	sram_mem[99666] = 16'b0000000000000000;
	sram_mem[99667] = 16'b0000000000000000;
	sram_mem[99668] = 16'b0000000000000000;
	sram_mem[99669] = 16'b0000000000000000;
	sram_mem[99670] = 16'b0000000000000000;
	sram_mem[99671] = 16'b0000000000000000;
	sram_mem[99672] = 16'b0000000000000000;
	sram_mem[99673] = 16'b0000000000000000;
	sram_mem[99674] = 16'b0000000000000000;
	sram_mem[99675] = 16'b0000000000000000;
	sram_mem[99676] = 16'b0000000000000000;
	sram_mem[99677] = 16'b0000000000000000;
	sram_mem[99678] = 16'b0000000000000000;
	sram_mem[99679] = 16'b0000000000000000;
	sram_mem[99680] = 16'b0000000000000000;
	sram_mem[99681] = 16'b0000000000000000;
	sram_mem[99682] = 16'b0000000000000000;
	sram_mem[99683] = 16'b0000000000000000;
	sram_mem[99684] = 16'b0000000000000000;
	sram_mem[99685] = 16'b0000000000000000;
	sram_mem[99686] = 16'b0000000000000000;
	sram_mem[99687] = 16'b0000000000000000;
	sram_mem[99688] = 16'b0000000000000000;
	sram_mem[99689] = 16'b0000000000000000;
	sram_mem[99690] = 16'b0000000000000000;
	sram_mem[99691] = 16'b0000000000000000;
	sram_mem[99692] = 16'b0000000000000000;
	sram_mem[99693] = 16'b0000000000000000;
	sram_mem[99694] = 16'b0000000000000000;
	sram_mem[99695] = 16'b0000000000000000;
	sram_mem[99696] = 16'b0000000000000000;
	sram_mem[99697] = 16'b0000000000000000;
	sram_mem[99698] = 16'b0000000000000000;
	sram_mem[99699] = 16'b0000000000000000;
	sram_mem[99700] = 16'b0000000000000000;
	sram_mem[99701] = 16'b0000000000000000;
	sram_mem[99702] = 16'b0000000000000000;
	sram_mem[99703] = 16'b0000000000000000;
	sram_mem[99704] = 16'b0000000000000000;
	sram_mem[99705] = 16'b0000000000000000;
	sram_mem[99706] = 16'b0000000000000000;
	sram_mem[99707] = 16'b0000000000000000;
	sram_mem[99708] = 16'b0000000000000000;
	sram_mem[99709] = 16'b0000000000000000;
	sram_mem[99710] = 16'b0000000000000000;
	sram_mem[99711] = 16'b0000000000000000;
	sram_mem[99712] = 16'b0000000000000000;
	sram_mem[99713] = 16'b0000000000000000;
	sram_mem[99714] = 16'b0000000000000000;
	sram_mem[99715] = 16'b0000000000000000;
	sram_mem[99716] = 16'b0000000000000000;
	sram_mem[99717] = 16'b0000000000000000;
	sram_mem[99718] = 16'b0000000000000000;
	sram_mem[99719] = 16'b0000000000000000;
	sram_mem[99720] = 16'b0000000000000000;
	sram_mem[99721] = 16'b0000000000000000;
	sram_mem[99722] = 16'b0000000000000000;
	sram_mem[99723] = 16'b0000000000000000;
	sram_mem[99724] = 16'b0000000000000000;
	sram_mem[99725] = 16'b0000000000000000;
	sram_mem[99726] = 16'b0000000000000000;
	sram_mem[99727] = 16'b0000000000000000;
	sram_mem[99728] = 16'b0000000000000000;
	sram_mem[99729] = 16'b0000000000000000;
	sram_mem[99730] = 16'b0000000000000000;
	sram_mem[99731] = 16'b0000000000000000;
	sram_mem[99732] = 16'b0000000000000000;
	sram_mem[99733] = 16'b0000000000000000;
	sram_mem[99734] = 16'b0000000000000000;
	sram_mem[99735] = 16'b0000000000000000;
	sram_mem[99736] = 16'b0000000000000000;
	sram_mem[99737] = 16'b0000000000000000;
	sram_mem[99738] = 16'b0000000000000000;
	sram_mem[99739] = 16'b0000000000000000;
	sram_mem[99740] = 16'b0000000000000000;
	sram_mem[99741] = 16'b0000000000000000;
	sram_mem[99742] = 16'b0000000000000000;
	sram_mem[99743] = 16'b0000000000000000;
	sram_mem[99744] = 16'b0000000000000000;
	sram_mem[99745] = 16'b0000000000000000;
	sram_mem[99746] = 16'b0000000000000000;
	sram_mem[99747] = 16'b0000000000000000;
	sram_mem[99748] = 16'b0000000000000000;
	sram_mem[99749] = 16'b0000000000000000;
	sram_mem[99750] = 16'b0000000000000000;
	sram_mem[99751] = 16'b0000000000000000;
	sram_mem[99752] = 16'b0000000000000000;
	sram_mem[99753] = 16'b0000000000000000;
	sram_mem[99754] = 16'b0000000000000000;
	sram_mem[99755] = 16'b0000000000000000;
	sram_mem[99756] = 16'b0000000000000000;
	sram_mem[99757] = 16'b0000000000000000;
	sram_mem[99758] = 16'b0000000000000000;
	sram_mem[99759] = 16'b0000000000000000;
	sram_mem[99760] = 16'b0000000000000000;
	sram_mem[99761] = 16'b0000000000000000;
	sram_mem[99762] = 16'b0000000000000000;
	sram_mem[99763] = 16'b0000000000000000;
	sram_mem[99764] = 16'b0000000000000000;
	sram_mem[99765] = 16'b0000000000000000;
	sram_mem[99766] = 16'b0000000000000000;
	sram_mem[99767] = 16'b0000000000000000;
	sram_mem[99768] = 16'b0000000000000000;
	sram_mem[99769] = 16'b0000000000000000;
	sram_mem[99770] = 16'b0000000000000000;
	sram_mem[99771] = 16'b0000000000000000;
	sram_mem[99772] = 16'b0000000000000000;
	sram_mem[99773] = 16'b0000000000000000;
	sram_mem[99774] = 16'b0000000000000000;
	sram_mem[99775] = 16'b0000000000000000;
	sram_mem[99776] = 16'b0000000000000000;
	sram_mem[99777] = 16'b0000000000000000;
	sram_mem[99778] = 16'b0000000000000000;
	sram_mem[99779] = 16'b0000000000000000;
	sram_mem[99780] = 16'b0000000000000000;
	sram_mem[99781] = 16'b0000000000000000;
	sram_mem[99782] = 16'b0000000000000000;
	sram_mem[99783] = 16'b0000000000000000;
	sram_mem[99784] = 16'b0000000000000000;
	sram_mem[99785] = 16'b0000000000000000;
	sram_mem[99786] = 16'b0000000000000000;
	sram_mem[99787] = 16'b0000000000000000;
	sram_mem[99788] = 16'b0000000000000000;
	sram_mem[99789] = 16'b0000000000000000;
	sram_mem[99790] = 16'b0000000000000000;
	sram_mem[99791] = 16'b0000000000000000;
	sram_mem[99792] = 16'b0000000000000000;
	sram_mem[99793] = 16'b0000000000000000;
	sram_mem[99794] = 16'b0000000000000000;
	sram_mem[99795] = 16'b0000000000000000;
	sram_mem[99796] = 16'b0000000000000000;
	sram_mem[99797] = 16'b0000000000000000;
	sram_mem[99798] = 16'b0000000000000000;
	sram_mem[99799] = 16'b0000000000000000;
	sram_mem[99800] = 16'b0000000000000000;
	sram_mem[99801] = 16'b0000000000000000;
	sram_mem[99802] = 16'b0000000000000000;
	sram_mem[99803] = 16'b0000000000000000;
	sram_mem[99804] = 16'b0000000000000000;
	sram_mem[99805] = 16'b0000000000000000;
	sram_mem[99806] = 16'b0000000000000000;
	sram_mem[99807] = 16'b0000000000000000;
	sram_mem[99808] = 16'b0000000000000000;
	sram_mem[99809] = 16'b0000000000000000;
	sram_mem[99810] = 16'b0000000000000000;
	sram_mem[99811] = 16'b0000000000000000;
	sram_mem[99812] = 16'b0000000000000000;
	sram_mem[99813] = 16'b0000000000000000;
	sram_mem[99814] = 16'b0000000000000000;
	sram_mem[99815] = 16'b0000000000000000;
	sram_mem[99816] = 16'b0000000000000000;
	sram_mem[99817] = 16'b0000000000000000;
	sram_mem[99818] = 16'b0000000000000000;
	sram_mem[99819] = 16'b0000000000000000;
	sram_mem[99820] = 16'b0000000000000000;
	sram_mem[99821] = 16'b0000000000000000;
	sram_mem[99822] = 16'b0000000000000000;
	sram_mem[99823] = 16'b0000000000000000;
	sram_mem[99824] = 16'b0000000000000000;
	sram_mem[99825] = 16'b0000000000000000;
	sram_mem[99826] = 16'b0000000000000000;
	sram_mem[99827] = 16'b0000000000000000;
	sram_mem[99828] = 16'b0000000000000000;
	sram_mem[99829] = 16'b0000000000000000;
	sram_mem[99830] = 16'b0000000000000000;
	sram_mem[99831] = 16'b0000000000000000;
	sram_mem[99832] = 16'b0000000000000000;
	sram_mem[99833] = 16'b0000000000000000;
	sram_mem[99834] = 16'b0000000000000000;
	sram_mem[99835] = 16'b0000000000000000;
	sram_mem[99836] = 16'b0000000000000000;
	sram_mem[99837] = 16'b0000000000000000;
	sram_mem[99838] = 16'b0000000000000000;
	sram_mem[99839] = 16'b0000000000000000;
	sram_mem[99840] = 16'b0000000000000000;
	sram_mem[99841] = 16'b0000000000000000;
	sram_mem[99842] = 16'b0000000000000000;
	sram_mem[99843] = 16'b0000000000000000;
	sram_mem[99844] = 16'b0000000000000000;
	sram_mem[99845] = 16'b0000000000000000;
	sram_mem[99846] = 16'b0000000000000000;
	sram_mem[99847] = 16'b0000000000000000;
	sram_mem[99848] = 16'b0000000000000000;
	sram_mem[99849] = 16'b0000000000000000;
	sram_mem[99850] = 16'b0000000000000000;
	sram_mem[99851] = 16'b0000000000000000;
	sram_mem[99852] = 16'b0000000000000000;
	sram_mem[99853] = 16'b0000000000000000;
	sram_mem[99854] = 16'b0000000000000000;
	sram_mem[99855] = 16'b0000000000000000;
	sram_mem[99856] = 16'b0000000000000000;
	sram_mem[99857] = 16'b0000000000000000;
	sram_mem[99858] = 16'b0000000000000000;
	sram_mem[99859] = 16'b0000000000000000;
	sram_mem[99860] = 16'b0000000000000000;
	sram_mem[99861] = 16'b0000000000000000;
	sram_mem[99862] = 16'b0000000000000000;
	sram_mem[99863] = 16'b0000000000000000;
	sram_mem[99864] = 16'b0000000000000000;
	sram_mem[99865] = 16'b0000000000000000;
	sram_mem[99866] = 16'b0000000000000000;
	sram_mem[99867] = 16'b0000000000000000;
	sram_mem[99868] = 16'b0000000000000000;
	sram_mem[99869] = 16'b0000000000000000;
	sram_mem[99870] = 16'b0000000000000000;
	sram_mem[99871] = 16'b0000000000000000;
	sram_mem[99872] = 16'b0000000000000000;
	sram_mem[99873] = 16'b0000000000000000;
	sram_mem[99874] = 16'b0000000000000000;
	sram_mem[99875] = 16'b0000000000000000;
	sram_mem[99876] = 16'b0000000000000000;
	sram_mem[99877] = 16'b0000000000000000;
	sram_mem[99878] = 16'b0000000000000000;
	sram_mem[99879] = 16'b0000000000000000;
	sram_mem[99880] = 16'b0000000000000000;
	sram_mem[99881] = 16'b0000000000000000;
	sram_mem[99882] = 16'b0000000000000000;
	sram_mem[99883] = 16'b0000000000000000;
	sram_mem[99884] = 16'b0000000000000000;
	sram_mem[99885] = 16'b0000000000000000;
	sram_mem[99886] = 16'b0000000000000000;
	sram_mem[99887] = 16'b0000000000000000;
	sram_mem[99888] = 16'b0000000000000000;
	sram_mem[99889] = 16'b0000000000000000;
	sram_mem[99890] = 16'b0000000000000000;
	sram_mem[99891] = 16'b0000000000000000;
	sram_mem[99892] = 16'b0000000000000000;
	sram_mem[99893] = 16'b0000000000000000;
	sram_mem[99894] = 16'b0000000000000000;
	sram_mem[99895] = 16'b0000000000000000;
	sram_mem[99896] = 16'b0000000000000000;
	sram_mem[99897] = 16'b0000000000000000;
	sram_mem[99898] = 16'b0000000000000000;
	sram_mem[99899] = 16'b0000000000000000;
	sram_mem[99900] = 16'b0000000000000000;
	sram_mem[99901] = 16'b0000000000000000;
	sram_mem[99902] = 16'b0000000000000000;
	sram_mem[99903] = 16'b0000000000000000;
	sram_mem[99904] = 16'b0000000000000000;
	sram_mem[99905] = 16'b0000000000000000;
	sram_mem[99906] = 16'b0000000000000000;
	sram_mem[99907] = 16'b0000000000000000;
	sram_mem[99908] = 16'b0000000000000000;
	sram_mem[99909] = 16'b0000000000000000;
	sram_mem[99910] = 16'b0000000000000000;
	sram_mem[99911] = 16'b0000000000000000;
	sram_mem[99912] = 16'b0000000000000000;
	sram_mem[99913] = 16'b0000000000000000;
	sram_mem[99914] = 16'b0000000000000000;
	sram_mem[99915] = 16'b0000000000000000;
	sram_mem[99916] = 16'b0000000000000000;
	sram_mem[99917] = 16'b0000000000000000;
	sram_mem[99918] = 16'b0000000000000000;
	sram_mem[99919] = 16'b0000000000000000;
	sram_mem[99920] = 16'b0000000000000000;
	sram_mem[99921] = 16'b0000000000000000;
	sram_mem[99922] = 16'b0000000000000000;
	sram_mem[99923] = 16'b0000000000000000;
	sram_mem[99924] = 16'b0000000000000000;
	sram_mem[99925] = 16'b0000000000000000;
	sram_mem[99926] = 16'b0000000000000000;
	sram_mem[99927] = 16'b0000000000000000;
	sram_mem[99928] = 16'b0000000000000000;
	sram_mem[99929] = 16'b0000000000000000;
	sram_mem[99930] = 16'b0000000000000000;
	sram_mem[99931] = 16'b0000000000000000;
	sram_mem[99932] = 16'b0000000000000000;
	sram_mem[99933] = 16'b0000000000000000;
	sram_mem[99934] = 16'b0000000000000000;
	sram_mem[99935] = 16'b0000000000000000;
	sram_mem[99936] = 16'b0000000000000000;
	sram_mem[99937] = 16'b0000000000000000;
	sram_mem[99938] = 16'b0000000000000000;
	sram_mem[99939] = 16'b0000000000000000;
	sram_mem[99940] = 16'b0000000000000000;
	sram_mem[99941] = 16'b0000000000000000;
	sram_mem[99942] = 16'b0000000000000000;
	sram_mem[99943] = 16'b0000000000000000;
	sram_mem[99944] = 16'b0000000000000000;
	sram_mem[99945] = 16'b0000000000000000;
	sram_mem[99946] = 16'b0000000000000000;
	sram_mem[99947] = 16'b0000000000000000;
	sram_mem[99948] = 16'b0000000000000000;
	sram_mem[99949] = 16'b0000000000000000;
	sram_mem[99950] = 16'b0000000000000000;
	sram_mem[99951] = 16'b0000000000000000;
	sram_mem[99952] = 16'b0000000000000000;
	sram_mem[99953] = 16'b0000000000000000;
	sram_mem[99954] = 16'b0000000000000000;
	sram_mem[99955] = 16'b0000000000000000;
	sram_mem[99956] = 16'b0000000000000000;
	sram_mem[99957] = 16'b0000000000000000;
	sram_mem[99958] = 16'b0000000000000000;
	sram_mem[99959] = 16'b0000000000000000;
	sram_mem[99960] = 16'b0000000000000000;
	sram_mem[99961] = 16'b0000000000000000;
	sram_mem[99962] = 16'b0000000000000000;
	sram_mem[99963] = 16'b0000000000000000;
	sram_mem[99964] = 16'b0000000000000000;
	sram_mem[99965] = 16'b0000000000000000;
	sram_mem[99966] = 16'b0000000000000000;
	sram_mem[99967] = 16'b0000000000000000;
	sram_mem[99968] = 16'b0000000000000000;
	sram_mem[99969] = 16'b0000000000000000;
	sram_mem[99970] = 16'b0000000000000000;
	sram_mem[99971] = 16'b0000000000000000;
	sram_mem[99972] = 16'b0000000000000000;
	sram_mem[99973] = 16'b0000000000000000;
	sram_mem[99974] = 16'b0000000000000000;
	sram_mem[99975] = 16'b0000000000000000;
	sram_mem[99976] = 16'b0000000000000000;
	sram_mem[99977] = 16'b0000000000000000;
	sram_mem[99978] = 16'b0000000000000000;
	sram_mem[99979] = 16'b0000000000000000;
	sram_mem[99980] = 16'b0000000000000000;
	sram_mem[99981] = 16'b0000000000000000;
	sram_mem[99982] = 16'b0000000000000000;
	sram_mem[99983] = 16'b0000000000000000;
	sram_mem[99984] = 16'b0000000000000000;
	sram_mem[99985] = 16'b0000000000000000;
	sram_mem[99986] = 16'b0000000000000000;
	sram_mem[99987] = 16'b0000000000000000;
	sram_mem[99988] = 16'b0000000000000000;
	sram_mem[99989] = 16'b0000000000000000;
	sram_mem[99990] = 16'b0000000000000000;
	sram_mem[99991] = 16'b0000000000000000;
	sram_mem[99992] = 16'b0000000000000000;
	sram_mem[99993] = 16'b0000000000000000;
	sram_mem[99994] = 16'b0000000000000000;
	sram_mem[99995] = 16'b0000000000000000;
	sram_mem[99996] = 16'b0000000000000000;
	sram_mem[99997] = 16'b0000000000000000;
	sram_mem[99998] = 16'b0000000000000000;
	sram_mem[99999] = 16'b0000000000000000;
	sram_mem[100000] = 16'b0000000000000000;
	sram_mem[100001] = 16'b0000000000000000;
	sram_mem[100002] = 16'b0000000000000000;
	sram_mem[100003] = 16'b0000000000000000;
	sram_mem[100004] = 16'b0000000000000000;
	sram_mem[100005] = 16'b0000000000000000;
	sram_mem[100006] = 16'b0000000000000000;
	sram_mem[100007] = 16'b0000000000000000;
	sram_mem[100008] = 16'b0000000000000000;
	sram_mem[100009] = 16'b0000000000000000;
	sram_mem[100010] = 16'b0000000000000000;
	sram_mem[100011] = 16'b0000000000000000;
	sram_mem[100012] = 16'b0000000000000000;
	sram_mem[100013] = 16'b0000000000000000;
	sram_mem[100014] = 16'b0000000000000000;
	sram_mem[100015] = 16'b0000000000000000;
	sram_mem[100016] = 16'b0000000000000000;
	sram_mem[100017] = 16'b0000000000000000;
	sram_mem[100018] = 16'b0000000000000000;
	sram_mem[100019] = 16'b0000000000000000;
	sram_mem[100020] = 16'b0000000000000000;
	sram_mem[100021] = 16'b0000000000000000;
	sram_mem[100022] = 16'b0000000000000000;
	sram_mem[100023] = 16'b0000000000000000;
	sram_mem[100024] = 16'b0000000000000000;
	sram_mem[100025] = 16'b0000000000000000;
	sram_mem[100026] = 16'b0000000000000000;
	sram_mem[100027] = 16'b0000000000000000;
	sram_mem[100028] = 16'b0000000000000000;
	sram_mem[100029] = 16'b0000000000000000;
	sram_mem[100030] = 16'b0000000000000000;
	sram_mem[100031] = 16'b0000000000000000;
	sram_mem[100032] = 16'b0000000000000000;
	sram_mem[100033] = 16'b0000000000000000;
	sram_mem[100034] = 16'b0000000000000000;
	sram_mem[100035] = 16'b0000000000000000;
	sram_mem[100036] = 16'b0000000000000000;
	sram_mem[100037] = 16'b0000000000000000;
	sram_mem[100038] = 16'b0000000000000000;
	sram_mem[100039] = 16'b0000000000000000;
	sram_mem[100040] = 16'b0000000000000000;
	sram_mem[100041] = 16'b0000000000000000;
	sram_mem[100042] = 16'b0000000000000000;
	sram_mem[100043] = 16'b0000000000000000;
	sram_mem[100044] = 16'b0000000000000000;
	sram_mem[100045] = 16'b0000000000000000;
	sram_mem[100046] = 16'b0000000000000000;
	sram_mem[100047] = 16'b0000000000000000;
	sram_mem[100048] = 16'b0000000000000000;
	sram_mem[100049] = 16'b0000000000000000;
	sram_mem[100050] = 16'b0000000000000000;
	sram_mem[100051] = 16'b0000000000000000;
	sram_mem[100052] = 16'b0000000000000000;
	sram_mem[100053] = 16'b0000000000000000;
	sram_mem[100054] = 16'b0000000000000000;
	sram_mem[100055] = 16'b0000000000000000;
	sram_mem[100056] = 16'b0000000000000000;
	sram_mem[100057] = 16'b0000000000000000;
	sram_mem[100058] = 16'b0000000000000000;
	sram_mem[100059] = 16'b0000000000000000;
	sram_mem[100060] = 16'b0000000000000000;
	sram_mem[100061] = 16'b0000000000000000;
	sram_mem[100062] = 16'b0000000000000000;
	sram_mem[100063] = 16'b0000000000000000;
	sram_mem[100064] = 16'b0000000000000000;
	sram_mem[100065] = 16'b0000000000000000;
	sram_mem[100066] = 16'b0000000000000000;
	sram_mem[100067] = 16'b0000000000000000;
	sram_mem[100068] = 16'b0000000000000000;
	sram_mem[100069] = 16'b0000000000000000;
	sram_mem[100070] = 16'b0000000000000000;
	sram_mem[100071] = 16'b0000000000000000;
	sram_mem[100072] = 16'b0000000000000000;
	sram_mem[100073] = 16'b0000000000000000;
	sram_mem[100074] = 16'b0000000000000000;
	sram_mem[100075] = 16'b0000000000000000;
	sram_mem[100076] = 16'b0000000000000000;
	sram_mem[100077] = 16'b0000000000000000;
	sram_mem[100078] = 16'b0000000000000000;
	sram_mem[100079] = 16'b0000000000000000;
	sram_mem[100080] = 16'b0000000000000000;
	sram_mem[100081] = 16'b0000000000000000;
	sram_mem[100082] = 16'b0000000000000000;
	sram_mem[100083] = 16'b0000000000000000;
	sram_mem[100084] = 16'b0000000000000000;
	sram_mem[100085] = 16'b0000000000000000;
	sram_mem[100086] = 16'b0000000000000000;
	sram_mem[100087] = 16'b0000000000000000;
	sram_mem[100088] = 16'b0000000000000000;
	sram_mem[100089] = 16'b0000000000000000;
	sram_mem[100090] = 16'b0000000000000000;
	sram_mem[100091] = 16'b0000000000000000;
	sram_mem[100092] = 16'b0000000000000000;
	sram_mem[100093] = 16'b0000000000000000;
	sram_mem[100094] = 16'b0000000000000000;
	sram_mem[100095] = 16'b0000000000000000;
	sram_mem[100096] = 16'b0000000000000000;
	sram_mem[100097] = 16'b0000000000000000;
	sram_mem[100098] = 16'b0000000000000000;
	sram_mem[100099] = 16'b0000000000000000;
	sram_mem[100100] = 16'b0000000000000000;
	sram_mem[100101] = 16'b0000000000000000;
	sram_mem[100102] = 16'b0000000000000000;
	sram_mem[100103] = 16'b0000000000000000;
	sram_mem[100104] = 16'b0000000000000000;
	sram_mem[100105] = 16'b0000000000000000;
	sram_mem[100106] = 16'b0000000000000000;
	sram_mem[100107] = 16'b0000000000000000;
	sram_mem[100108] = 16'b0000000000000000;
	sram_mem[100109] = 16'b0000000000000000;
	sram_mem[100110] = 16'b0000000000000000;
	sram_mem[100111] = 16'b0000000000000000;
	sram_mem[100112] = 16'b0000000000000000;
	sram_mem[100113] = 16'b0000000000000000;
	sram_mem[100114] = 16'b0000000000000000;
	sram_mem[100115] = 16'b0000000000000000;
	sram_mem[100116] = 16'b0000000000000000;
	sram_mem[100117] = 16'b0000000000000000;
	sram_mem[100118] = 16'b0000000000000000;
	sram_mem[100119] = 16'b0000000000000000;
	sram_mem[100120] = 16'b0000000000000000;
	sram_mem[100121] = 16'b0000000000000000;
	sram_mem[100122] = 16'b0000000000000000;
	sram_mem[100123] = 16'b0000000000000000;
	sram_mem[100124] = 16'b0000000000000000;
	sram_mem[100125] = 16'b0000000000000000;
	sram_mem[100126] = 16'b0000000000000000;
	sram_mem[100127] = 16'b0000000000000000;
	sram_mem[100128] = 16'b0000000000000000;
	sram_mem[100129] = 16'b0000000000000000;
	sram_mem[100130] = 16'b0000000000000000;
	sram_mem[100131] = 16'b0000000000000000;
	sram_mem[100132] = 16'b0000000000000000;
	sram_mem[100133] = 16'b0000000000000000;
	sram_mem[100134] = 16'b0000000000000000;
	sram_mem[100135] = 16'b0000000000000000;
	sram_mem[100136] = 16'b0000000000000000;
	sram_mem[100137] = 16'b0000000000000000;
	sram_mem[100138] = 16'b0000000000000000;
	sram_mem[100139] = 16'b0000000000000000;
	sram_mem[100140] = 16'b0000000000000000;
	sram_mem[100141] = 16'b0000000000000000;
	sram_mem[100142] = 16'b0000000000000000;
	sram_mem[100143] = 16'b0000000000000000;
	sram_mem[100144] = 16'b0000000000000000;
	sram_mem[100145] = 16'b0000000000000000;
	sram_mem[100146] = 16'b0000000000000000;
	sram_mem[100147] = 16'b0000000000000000;
	sram_mem[100148] = 16'b0000000000000000;
	sram_mem[100149] = 16'b0000000000000000;
	sram_mem[100150] = 16'b0000000000000000;
	sram_mem[100151] = 16'b0000000000000000;
	sram_mem[100152] = 16'b0000000000000000;
	sram_mem[100153] = 16'b0000000000000000;
	sram_mem[100154] = 16'b0000000000000000;
	sram_mem[100155] = 16'b0000000000000000;
	sram_mem[100156] = 16'b0000000000000000;
	sram_mem[100157] = 16'b0000000000000000;
	sram_mem[100158] = 16'b0000000000000000;
	sram_mem[100159] = 16'b0000000000000000;
	sram_mem[100160] = 16'b0000000000000000;
	sram_mem[100161] = 16'b0000000000000000;
	sram_mem[100162] = 16'b0000000000000000;
	sram_mem[100163] = 16'b0000000000000000;
	sram_mem[100164] = 16'b0000000000000000;
	sram_mem[100165] = 16'b0000000000000000;
	sram_mem[100166] = 16'b0000000000000000;
	sram_mem[100167] = 16'b0000000000000000;
	sram_mem[100168] = 16'b0000000000000000;
	sram_mem[100169] = 16'b0000000000000000;
	sram_mem[100170] = 16'b0000000000000000;
	sram_mem[100171] = 16'b0000000000000000;
	sram_mem[100172] = 16'b0000000000000000;
	sram_mem[100173] = 16'b0000000000000000;
	sram_mem[100174] = 16'b0000000000000000;
	sram_mem[100175] = 16'b0000000000000000;
	sram_mem[100176] = 16'b0000000000000000;
	sram_mem[100177] = 16'b0000000000000000;
	sram_mem[100178] = 16'b0000000000000000;
	sram_mem[100179] = 16'b0000000000000000;
	sram_mem[100180] = 16'b0000000000000000;
	sram_mem[100181] = 16'b0000000000000000;
	sram_mem[100182] = 16'b0000000000000000;
	sram_mem[100183] = 16'b0000000000000000;
	sram_mem[100184] = 16'b0000000000000000;
	sram_mem[100185] = 16'b0000000000000000;
	sram_mem[100186] = 16'b0000000000000000;
	sram_mem[100187] = 16'b0000000000000000;
	sram_mem[100188] = 16'b0000000000000000;
	sram_mem[100189] = 16'b0000000000000000;
	sram_mem[100190] = 16'b0000000000000000;
	sram_mem[100191] = 16'b0000000000000000;
	sram_mem[100192] = 16'b0000000000000000;
	sram_mem[100193] = 16'b0000000000000000;
	sram_mem[100194] = 16'b0000000000000000;
	sram_mem[100195] = 16'b0000000000000000;
	sram_mem[100196] = 16'b0000000000000000;
	sram_mem[100197] = 16'b0000000000000000;
	sram_mem[100198] = 16'b0000000000000000;
	sram_mem[100199] = 16'b0000000000000000;
	sram_mem[100200] = 16'b0000000000000000;
	sram_mem[100201] = 16'b0000000000000000;
	sram_mem[100202] = 16'b0000000000000000;
	sram_mem[100203] = 16'b0000000000000000;
	sram_mem[100204] = 16'b0000000000000000;
	sram_mem[100205] = 16'b0000000000000000;
	sram_mem[100206] = 16'b0000000000000000;
	sram_mem[100207] = 16'b0000000000000000;
	sram_mem[100208] = 16'b0000000000000000;
	sram_mem[100209] = 16'b0000000000000000;
	sram_mem[100210] = 16'b0000000000000000;
	sram_mem[100211] = 16'b0000000000000000;
	sram_mem[100212] = 16'b0000000000000000;
	sram_mem[100213] = 16'b0000000000000000;
	sram_mem[100214] = 16'b0000000000000000;
	sram_mem[100215] = 16'b0000000000000000;
	sram_mem[100216] = 16'b0000000000000000;
	sram_mem[100217] = 16'b0000000000000000;
	sram_mem[100218] = 16'b0000000000000000;
	sram_mem[100219] = 16'b0000000000000000;
	sram_mem[100220] = 16'b0000000000000000;
	sram_mem[100221] = 16'b0000000000000000;
	sram_mem[100222] = 16'b0000000000000000;
	sram_mem[100223] = 16'b0000000000000000;
	sram_mem[100224] = 16'b0000000000000000;
	sram_mem[100225] = 16'b0000000000000000;
	sram_mem[100226] = 16'b0000000000000000;
	sram_mem[100227] = 16'b0000000000000000;
	sram_mem[100228] = 16'b0000000000000000;
	sram_mem[100229] = 16'b0000000000000000;
	sram_mem[100230] = 16'b0000000000000000;
	sram_mem[100231] = 16'b0000000000000000;
	sram_mem[100232] = 16'b0000000000000000;
	sram_mem[100233] = 16'b0000000000000000;
	sram_mem[100234] = 16'b0000000000000000;
	sram_mem[100235] = 16'b0000000000000000;
	sram_mem[100236] = 16'b0000000000000000;
	sram_mem[100237] = 16'b0000000000000000;
	sram_mem[100238] = 16'b0000000000000000;
	sram_mem[100239] = 16'b0000000000000000;
	sram_mem[100240] = 16'b0000000000000000;
	sram_mem[100241] = 16'b0000000000000000;
	sram_mem[100242] = 16'b0000000000000000;
	sram_mem[100243] = 16'b0000000000000000;
	sram_mem[100244] = 16'b0000000000000000;
	sram_mem[100245] = 16'b0000000000000000;
	sram_mem[100246] = 16'b0000000000000000;
	sram_mem[100247] = 16'b0000000000000000;
	sram_mem[100248] = 16'b0000000000000000;
	sram_mem[100249] = 16'b0000000000000000;
	sram_mem[100250] = 16'b0000000000000000;
	sram_mem[100251] = 16'b0000000000000000;
	sram_mem[100252] = 16'b0000000000000000;
	sram_mem[100253] = 16'b0000000000000000;
	sram_mem[100254] = 16'b0000000000000000;
	sram_mem[100255] = 16'b0000000000000000;
	sram_mem[100256] = 16'b0000000000000000;
	sram_mem[100257] = 16'b0000000000000000;
	sram_mem[100258] = 16'b0000000000000000;
	sram_mem[100259] = 16'b0000000000000000;
	sram_mem[100260] = 16'b0000000000000000;
	sram_mem[100261] = 16'b0000000000000000;
	sram_mem[100262] = 16'b0000000000000000;
	sram_mem[100263] = 16'b0000000000000000;
	sram_mem[100264] = 16'b0000000000000000;
	sram_mem[100265] = 16'b0000000000000000;
	sram_mem[100266] = 16'b0000000000000000;
	sram_mem[100267] = 16'b0000000000000000;
	sram_mem[100268] = 16'b0000000000000000;
	sram_mem[100269] = 16'b0000000000000000;
	sram_mem[100270] = 16'b0000000000000000;
	sram_mem[100271] = 16'b0000000000000000;
	sram_mem[100272] = 16'b0000000000000000;
	sram_mem[100273] = 16'b0000000000000000;
	sram_mem[100274] = 16'b0000000000000000;
	sram_mem[100275] = 16'b0000000000000000;
	sram_mem[100276] = 16'b0000000000000000;
	sram_mem[100277] = 16'b0000000000000000;
	sram_mem[100278] = 16'b0000000000000000;
	sram_mem[100279] = 16'b0000000000000000;
	sram_mem[100280] = 16'b0000000000000000;
	sram_mem[100281] = 16'b0000000000000000;
	sram_mem[100282] = 16'b0000000000000000;
	sram_mem[100283] = 16'b0000000000000000;
	sram_mem[100284] = 16'b0000000000000000;
	sram_mem[100285] = 16'b0000000000000000;
	sram_mem[100286] = 16'b0000000000000000;
	sram_mem[100287] = 16'b0000000000000000;
	sram_mem[100288] = 16'b0000000000000000;
	sram_mem[100289] = 16'b0000000000000000;
	sram_mem[100290] = 16'b0000000000000000;
	sram_mem[100291] = 16'b0000000000000000;
	sram_mem[100292] = 16'b0000000000000000;
	sram_mem[100293] = 16'b0000000000000000;
	sram_mem[100294] = 16'b0000000000000000;
	sram_mem[100295] = 16'b0000000000000000;
	sram_mem[100296] = 16'b0000000000000000;
	sram_mem[100297] = 16'b0000000000000000;
	sram_mem[100298] = 16'b0000000000000000;
	sram_mem[100299] = 16'b0000000000000000;
	sram_mem[100300] = 16'b0000000000000000;
	sram_mem[100301] = 16'b0000000000000000;
	sram_mem[100302] = 16'b0000000000000000;
	sram_mem[100303] = 16'b0000000000000000;
	sram_mem[100304] = 16'b0000000000000000;
	sram_mem[100305] = 16'b0000000000000000;
	sram_mem[100306] = 16'b0000000000000000;
	sram_mem[100307] = 16'b0000000000000000;
	sram_mem[100308] = 16'b0000000000000000;
	sram_mem[100309] = 16'b0000000000000000;
	sram_mem[100310] = 16'b0000000000000000;
	sram_mem[100311] = 16'b0000000000000000;
	sram_mem[100312] = 16'b0000000000000000;
	sram_mem[100313] = 16'b0000000000000000;
	sram_mem[100314] = 16'b0000000000000000;
	sram_mem[100315] = 16'b0000000000000000;
	sram_mem[100316] = 16'b0000000000000000;
	sram_mem[100317] = 16'b0000000000000000;
	sram_mem[100318] = 16'b0000000000000000;
	sram_mem[100319] = 16'b0000000000000000;
	sram_mem[100320] = 16'b0000000000000000;
	sram_mem[100321] = 16'b0000000000000000;
	sram_mem[100322] = 16'b0000000000000000;
	sram_mem[100323] = 16'b0000000000000000;
	sram_mem[100324] = 16'b0000000000000000;
	sram_mem[100325] = 16'b0000000000000000;
	sram_mem[100326] = 16'b0000000000000000;
	sram_mem[100327] = 16'b0000000000000000;
	sram_mem[100328] = 16'b0000000000000000;
	sram_mem[100329] = 16'b0000000000000000;
	sram_mem[100330] = 16'b0000000000000000;
	sram_mem[100331] = 16'b0000000000000000;
	sram_mem[100332] = 16'b0000000000000000;
	sram_mem[100333] = 16'b0000000000000000;
	sram_mem[100334] = 16'b0000000000000000;
	sram_mem[100335] = 16'b0000000000000000;
	sram_mem[100336] = 16'b0000000000000000;
	sram_mem[100337] = 16'b0000000000000000;
	sram_mem[100338] = 16'b0000000000000000;
	sram_mem[100339] = 16'b0000000000000000;
	sram_mem[100340] = 16'b0000000000000000;
	sram_mem[100341] = 16'b0000000000000000;
	sram_mem[100342] = 16'b0000000000000000;
	sram_mem[100343] = 16'b0000000000000000;
	sram_mem[100344] = 16'b0000000000000000;
	sram_mem[100345] = 16'b0000000000000000;
	sram_mem[100346] = 16'b0000000000000000;
	sram_mem[100347] = 16'b0000000000000000;
	sram_mem[100348] = 16'b0000000000000000;
	sram_mem[100349] = 16'b0000000000000000;
	sram_mem[100350] = 16'b0000000000000000;
	sram_mem[100351] = 16'b0000000000000000;
	sram_mem[100352] = 16'b0000000000000000;
	sram_mem[100353] = 16'b0000000000000000;
	sram_mem[100354] = 16'b0000000000000000;
	sram_mem[100355] = 16'b0000000000000000;
	sram_mem[100356] = 16'b0000000000000000;
	sram_mem[100357] = 16'b0000000000000000;
	sram_mem[100358] = 16'b0000000000000000;
	sram_mem[100359] = 16'b0000000000000000;
	sram_mem[100360] = 16'b0000000000000000;
	sram_mem[100361] = 16'b0000000000000000;
	sram_mem[100362] = 16'b0000000000000000;
	sram_mem[100363] = 16'b0000000000000000;
	sram_mem[100364] = 16'b0000000000000000;
	sram_mem[100365] = 16'b0000000000000000;
	sram_mem[100366] = 16'b0000000000000000;
	sram_mem[100367] = 16'b0000000000000000;
	sram_mem[100368] = 16'b0000000000000000;
	sram_mem[100369] = 16'b0000000000000000;
	sram_mem[100370] = 16'b0000000000000000;
	sram_mem[100371] = 16'b0000000000000000;
	sram_mem[100372] = 16'b0000000000000000;
	sram_mem[100373] = 16'b0000000000000000;
	sram_mem[100374] = 16'b0000000000000000;
	sram_mem[100375] = 16'b0000000000000000;
	sram_mem[100376] = 16'b0000000000000000;
	sram_mem[100377] = 16'b0000000000000000;
	sram_mem[100378] = 16'b0000000000000000;
	sram_mem[100379] = 16'b0000000000000000;
	sram_mem[100380] = 16'b0000000000000000;
	sram_mem[100381] = 16'b0000000000000000;
	sram_mem[100382] = 16'b0000000000000000;
	sram_mem[100383] = 16'b0000000000000000;
	sram_mem[100384] = 16'b0000000000000000;
	sram_mem[100385] = 16'b0000000000000000;
	sram_mem[100386] = 16'b0000000000000000;
	sram_mem[100387] = 16'b0000000000000000;
	sram_mem[100388] = 16'b0000000000000000;
	sram_mem[100389] = 16'b0000000000000000;
	sram_mem[100390] = 16'b0000000000000000;
	sram_mem[100391] = 16'b0000000000000000;
	sram_mem[100392] = 16'b0000000000000000;
	sram_mem[100393] = 16'b0000000000000000;
	sram_mem[100394] = 16'b0000000000000000;
	sram_mem[100395] = 16'b0000000000000000;
	sram_mem[100396] = 16'b0000000000000000;
	sram_mem[100397] = 16'b0000000000000000;
	sram_mem[100398] = 16'b0000000000000000;
	sram_mem[100399] = 16'b0000000000000000;
	sram_mem[100400] = 16'b0000000000000000;
	sram_mem[100401] = 16'b0000000000000000;
	sram_mem[100402] = 16'b0000000000000000;
	sram_mem[100403] = 16'b0000000000000000;
	sram_mem[100404] = 16'b0000000000000000;
	sram_mem[100405] = 16'b0000000000000000;
	sram_mem[100406] = 16'b0000000000000000;
	sram_mem[100407] = 16'b0000000000000000;
	sram_mem[100408] = 16'b0000000000000000;
	sram_mem[100409] = 16'b0000000000000000;
	sram_mem[100410] = 16'b0000000000000000;
	sram_mem[100411] = 16'b0000000000000000;
	sram_mem[100412] = 16'b0000000000000000;
	sram_mem[100413] = 16'b0000000000000000;
	sram_mem[100414] = 16'b0000000000000000;
	sram_mem[100415] = 16'b0000000000000000;
	sram_mem[100416] = 16'b0000000000000000;
	sram_mem[100417] = 16'b0000000000000000;
	sram_mem[100418] = 16'b0000000000000000;
	sram_mem[100419] = 16'b0000000000000000;
	sram_mem[100420] = 16'b0000000000000000;
	sram_mem[100421] = 16'b0000000000000000;
	sram_mem[100422] = 16'b0000000000000000;
	sram_mem[100423] = 16'b0000000000000000;
	sram_mem[100424] = 16'b0000000000000000;
	sram_mem[100425] = 16'b0000000000000000;
	sram_mem[100426] = 16'b0000000000000000;
	sram_mem[100427] = 16'b0000000000000000;
	sram_mem[100428] = 16'b0000000000000000;
	sram_mem[100429] = 16'b0000000000000000;
	sram_mem[100430] = 16'b0000000000000000;
	sram_mem[100431] = 16'b0000000000000000;
	sram_mem[100432] = 16'b0000000000000000;
	sram_mem[100433] = 16'b0000000000000000;
	sram_mem[100434] = 16'b0000000000000000;
	sram_mem[100435] = 16'b0000000000000000;
	sram_mem[100436] = 16'b0000000000000000;
	sram_mem[100437] = 16'b0000000000000000;
	sram_mem[100438] = 16'b0000000000000000;
	sram_mem[100439] = 16'b0000000000000000;
	sram_mem[100440] = 16'b0000000000000000;
	sram_mem[100441] = 16'b0000000000000000;
	sram_mem[100442] = 16'b0000000000000000;
	sram_mem[100443] = 16'b0000000000000000;
	sram_mem[100444] = 16'b0000000000000000;
	sram_mem[100445] = 16'b0000000000000000;
	sram_mem[100446] = 16'b0000000000000000;
	sram_mem[100447] = 16'b0000000000000000;
	sram_mem[100448] = 16'b0000000000000000;
	sram_mem[100449] = 16'b0000000000000000;
	sram_mem[100450] = 16'b0000000000000000;
	sram_mem[100451] = 16'b0000000000000000;
	sram_mem[100452] = 16'b0000000000000000;
	sram_mem[100453] = 16'b0000000000000000;
	sram_mem[100454] = 16'b0000000000000000;
	sram_mem[100455] = 16'b0000000000000000;
	sram_mem[100456] = 16'b0000000000000000;
	sram_mem[100457] = 16'b0000000000000000;
	sram_mem[100458] = 16'b0000000000000000;
	sram_mem[100459] = 16'b0000000000000000;
	sram_mem[100460] = 16'b0000000000000000;
	sram_mem[100461] = 16'b0000000000000000;
	sram_mem[100462] = 16'b0000000000000000;
	sram_mem[100463] = 16'b0000000000000000;
	sram_mem[100464] = 16'b0000000000000000;
	sram_mem[100465] = 16'b0000000000000000;
	sram_mem[100466] = 16'b0000000000000000;
	sram_mem[100467] = 16'b0000000000000000;
	sram_mem[100468] = 16'b0000000000000000;
	sram_mem[100469] = 16'b0000000000000000;
	sram_mem[100470] = 16'b0000000000000000;
	sram_mem[100471] = 16'b0000000000000000;
	sram_mem[100472] = 16'b0000000000000000;
	sram_mem[100473] = 16'b0000000000000000;
	sram_mem[100474] = 16'b0000000000000000;
	sram_mem[100475] = 16'b0000000000000000;
	sram_mem[100476] = 16'b0000000000000000;
	sram_mem[100477] = 16'b0000000000000000;
	sram_mem[100478] = 16'b0000000000000000;
	sram_mem[100479] = 16'b0000000000000000;
	sram_mem[100480] = 16'b0000000000000000;
	sram_mem[100481] = 16'b0000000000000000;
	sram_mem[100482] = 16'b0000000000000000;
	sram_mem[100483] = 16'b0000000000000000;
	sram_mem[100484] = 16'b0000000000000000;
	sram_mem[100485] = 16'b0000000000000000;
	sram_mem[100486] = 16'b0000000000000000;
	sram_mem[100487] = 16'b0000000000000000;
	sram_mem[100488] = 16'b0000000000000000;
	sram_mem[100489] = 16'b0000000000000000;
	sram_mem[100490] = 16'b0000000000000000;
	sram_mem[100491] = 16'b0000000000000000;
	sram_mem[100492] = 16'b0000000000000000;
	sram_mem[100493] = 16'b0000000000000000;
	sram_mem[100494] = 16'b0000000000000000;
	sram_mem[100495] = 16'b0000000000000000;
	sram_mem[100496] = 16'b0000000000000000;
	sram_mem[100497] = 16'b0000000000000000;
	sram_mem[100498] = 16'b0000000000000000;
	sram_mem[100499] = 16'b0000000000000000;
	sram_mem[100500] = 16'b0000000000000000;
	sram_mem[100501] = 16'b0000000000000000;
	sram_mem[100502] = 16'b0000000000000000;
	sram_mem[100503] = 16'b0000000000000000;
	sram_mem[100504] = 16'b0000000000000000;
	sram_mem[100505] = 16'b0000000000000000;
	sram_mem[100506] = 16'b0000000000000000;
	sram_mem[100507] = 16'b0000000000000000;
	sram_mem[100508] = 16'b0000000000000000;
	sram_mem[100509] = 16'b0000000000000000;
	sram_mem[100510] = 16'b0000000000000000;
	sram_mem[100511] = 16'b0000000000000000;
	sram_mem[100512] = 16'b0000000000000000;
	sram_mem[100513] = 16'b0000000000000000;
	sram_mem[100514] = 16'b0000000000000000;
	sram_mem[100515] = 16'b0000000000000000;
	sram_mem[100516] = 16'b0000000000000000;
	sram_mem[100517] = 16'b0000000000000000;
	sram_mem[100518] = 16'b0000000000000000;
	sram_mem[100519] = 16'b0000000000000000;
	sram_mem[100520] = 16'b0000000000000000;
	sram_mem[100521] = 16'b0000000000000000;
	sram_mem[100522] = 16'b0000000000000000;
	sram_mem[100523] = 16'b0000000000000000;
	sram_mem[100524] = 16'b0000000000000000;
	sram_mem[100525] = 16'b0000000000000000;
	sram_mem[100526] = 16'b0000000000000000;
	sram_mem[100527] = 16'b0000000000000000;
	sram_mem[100528] = 16'b0000000000000000;
	sram_mem[100529] = 16'b0000000000000000;
	sram_mem[100530] = 16'b0000000000000000;
	sram_mem[100531] = 16'b0000000000000000;
	sram_mem[100532] = 16'b0000000000000000;
	sram_mem[100533] = 16'b0000000000000000;
	sram_mem[100534] = 16'b0000000000000000;
	sram_mem[100535] = 16'b0000000000000000;
	sram_mem[100536] = 16'b0000000000000000;
	sram_mem[100537] = 16'b0000000000000000;
	sram_mem[100538] = 16'b0000000000000000;
	sram_mem[100539] = 16'b0000000000000000;
	sram_mem[100540] = 16'b0000000000000000;
	sram_mem[100541] = 16'b0000000000000000;
	sram_mem[100542] = 16'b0000000000000000;
	sram_mem[100543] = 16'b0000000000000000;
	sram_mem[100544] = 16'b0000000000000000;
	sram_mem[100545] = 16'b0000000000000000;
	sram_mem[100546] = 16'b0000000000000000;
	sram_mem[100547] = 16'b0000000000000000;
	sram_mem[100548] = 16'b0000000000000000;
	sram_mem[100549] = 16'b0000000000000000;
	sram_mem[100550] = 16'b0000000000000000;
	sram_mem[100551] = 16'b0000000000000000;
	sram_mem[100552] = 16'b0000000000000000;
	sram_mem[100553] = 16'b0000000000000000;
	sram_mem[100554] = 16'b0000000000000000;
	sram_mem[100555] = 16'b0000000000000000;
	sram_mem[100556] = 16'b0000000000000000;
	sram_mem[100557] = 16'b0000000000000000;
	sram_mem[100558] = 16'b0000000000000000;
	sram_mem[100559] = 16'b0000000000000000;
	sram_mem[100560] = 16'b0000000000000000;
	sram_mem[100561] = 16'b0000000000000000;
	sram_mem[100562] = 16'b0000000000000000;
	sram_mem[100563] = 16'b0000000000000000;
	sram_mem[100564] = 16'b0000000000000000;
	sram_mem[100565] = 16'b0000000000000000;
	sram_mem[100566] = 16'b0000000000000000;
	sram_mem[100567] = 16'b0000000000000000;
	sram_mem[100568] = 16'b0000000000000000;
	sram_mem[100569] = 16'b0000000000000000;
	sram_mem[100570] = 16'b0000000000000000;
	sram_mem[100571] = 16'b0000000000000000;
	sram_mem[100572] = 16'b0000000000000000;
	sram_mem[100573] = 16'b0000000000000000;
	sram_mem[100574] = 16'b0000000000000000;
	sram_mem[100575] = 16'b0000000000000000;
	sram_mem[100576] = 16'b0000000000000000;
	sram_mem[100577] = 16'b0000000000000000;
	sram_mem[100578] = 16'b0000000000000000;
	sram_mem[100579] = 16'b0000000000000000;
	sram_mem[100580] = 16'b0000000000000000;
	sram_mem[100581] = 16'b0000000000000000;
	sram_mem[100582] = 16'b0000000000000000;
	sram_mem[100583] = 16'b0000000000000000;
	sram_mem[100584] = 16'b0000000000000000;
	sram_mem[100585] = 16'b0000000000000000;
	sram_mem[100586] = 16'b0000000000000000;
	sram_mem[100587] = 16'b0000000000000000;
	sram_mem[100588] = 16'b0000000000000000;
	sram_mem[100589] = 16'b0000000000000000;
	sram_mem[100590] = 16'b0000000000000000;
	sram_mem[100591] = 16'b0000000000000000;
	sram_mem[100592] = 16'b0000000000000000;
	sram_mem[100593] = 16'b0000000000000000;
	sram_mem[100594] = 16'b0000000000000000;
	sram_mem[100595] = 16'b0000000000000000;
	sram_mem[100596] = 16'b0000000000000000;
	sram_mem[100597] = 16'b0000000000000000;
	sram_mem[100598] = 16'b0000000000000000;
	sram_mem[100599] = 16'b0000000000000000;
	sram_mem[100600] = 16'b0000000000000000;
	sram_mem[100601] = 16'b0000000000000000;
	sram_mem[100602] = 16'b0000000000000000;
	sram_mem[100603] = 16'b0000000000000000;
	sram_mem[100604] = 16'b0000000000000000;
	sram_mem[100605] = 16'b0000000000000000;
	sram_mem[100606] = 16'b0000000000000000;
	sram_mem[100607] = 16'b0000000000000000;
	sram_mem[100608] = 16'b0000000000000000;
	sram_mem[100609] = 16'b0000000000000000;
	sram_mem[100610] = 16'b0000000000000000;
	sram_mem[100611] = 16'b0000000000000000;
	sram_mem[100612] = 16'b0000000000000000;
	sram_mem[100613] = 16'b0000000000000000;
	sram_mem[100614] = 16'b0000000000000000;
	sram_mem[100615] = 16'b0000000000000000;
	sram_mem[100616] = 16'b0000000000000000;
	sram_mem[100617] = 16'b0000000000000000;
	sram_mem[100618] = 16'b0000000000000000;
	sram_mem[100619] = 16'b0000000000000000;
	sram_mem[100620] = 16'b0000000000000000;
	sram_mem[100621] = 16'b0000000000000000;
	sram_mem[100622] = 16'b0000000000000000;
	sram_mem[100623] = 16'b0000000000000000;
	sram_mem[100624] = 16'b0000000000000000;
	sram_mem[100625] = 16'b0000000000000000;
	sram_mem[100626] = 16'b0000000000000000;
	sram_mem[100627] = 16'b0000000000000000;
	sram_mem[100628] = 16'b0000000000000000;
	sram_mem[100629] = 16'b0000000000000000;
	sram_mem[100630] = 16'b0000000000000000;
	sram_mem[100631] = 16'b0000000000000000;
	sram_mem[100632] = 16'b0000000000000000;
	sram_mem[100633] = 16'b0000000000000000;
	sram_mem[100634] = 16'b0000000000000000;
	sram_mem[100635] = 16'b0000000000000000;
	sram_mem[100636] = 16'b0000000000000000;
	sram_mem[100637] = 16'b0000000000000000;
	sram_mem[100638] = 16'b0000000000000000;
	sram_mem[100639] = 16'b0000000000000000;
	sram_mem[100640] = 16'b0000000000000000;
	sram_mem[100641] = 16'b0000000000000000;
	sram_mem[100642] = 16'b0000000000000000;
	sram_mem[100643] = 16'b0000000000000000;
	sram_mem[100644] = 16'b0000000000000000;
	sram_mem[100645] = 16'b0000000000000000;
	sram_mem[100646] = 16'b0000000000000000;
	sram_mem[100647] = 16'b0000000000000000;
	sram_mem[100648] = 16'b0000000000000000;
	sram_mem[100649] = 16'b0000000000000000;
	sram_mem[100650] = 16'b0000000000000000;
	sram_mem[100651] = 16'b0000000000000000;
	sram_mem[100652] = 16'b0000000000000000;
	sram_mem[100653] = 16'b0000000000000000;
	sram_mem[100654] = 16'b0000000000000000;
	sram_mem[100655] = 16'b0000000000000000;
	sram_mem[100656] = 16'b0000000000000000;
	sram_mem[100657] = 16'b0000000000000000;
	sram_mem[100658] = 16'b0000000000000000;
	sram_mem[100659] = 16'b0000000000000000;
	sram_mem[100660] = 16'b0000000000000000;
	sram_mem[100661] = 16'b0000000000000000;
	sram_mem[100662] = 16'b0000000000000000;
	sram_mem[100663] = 16'b0000000000000000;
	sram_mem[100664] = 16'b0000000000000000;
	sram_mem[100665] = 16'b0000000000000000;
	sram_mem[100666] = 16'b0000000000000000;
	sram_mem[100667] = 16'b0000000000000000;
	sram_mem[100668] = 16'b0000000000000000;
	sram_mem[100669] = 16'b0000000000000000;
	sram_mem[100670] = 16'b0000000000000000;
	sram_mem[100671] = 16'b0000000000000000;
	sram_mem[100672] = 16'b0000000000000000;
	sram_mem[100673] = 16'b0000000000000000;
	sram_mem[100674] = 16'b0000000000000000;
	sram_mem[100675] = 16'b0000000000000000;
	sram_mem[100676] = 16'b0000000000000000;
	sram_mem[100677] = 16'b0000000000000000;
	sram_mem[100678] = 16'b0000000000000000;
	sram_mem[100679] = 16'b0000000000000000;
	sram_mem[100680] = 16'b0000000000000000;
	sram_mem[100681] = 16'b0000000000000000;
	sram_mem[100682] = 16'b0000000000000000;
	sram_mem[100683] = 16'b0000000000000000;
	sram_mem[100684] = 16'b0000000000000000;
	sram_mem[100685] = 16'b0000000000000000;
	sram_mem[100686] = 16'b0000000000000000;
	sram_mem[100687] = 16'b0000000000000000;
	sram_mem[100688] = 16'b0000000000000000;
	sram_mem[100689] = 16'b0000000000000000;
	sram_mem[100690] = 16'b0000000000000000;
	sram_mem[100691] = 16'b0000000000000000;
	sram_mem[100692] = 16'b0000000000000000;
	sram_mem[100693] = 16'b0000000000000000;
	sram_mem[100694] = 16'b0000000000000000;
	sram_mem[100695] = 16'b0000000000000000;
	sram_mem[100696] = 16'b0000000000000000;
	sram_mem[100697] = 16'b0000000000000000;
	sram_mem[100698] = 16'b0000000000000000;
	sram_mem[100699] = 16'b0000000000000000;
	sram_mem[100700] = 16'b0000000000000000;
	sram_mem[100701] = 16'b0000000000000000;
	sram_mem[100702] = 16'b0000000000000000;
	sram_mem[100703] = 16'b0000000000000000;
	sram_mem[100704] = 16'b0000000000000000;
	sram_mem[100705] = 16'b0000000000000000;
	sram_mem[100706] = 16'b0000000000000000;
	sram_mem[100707] = 16'b0000000000000000;
	sram_mem[100708] = 16'b0000000000000000;
	sram_mem[100709] = 16'b0000000000000000;
	sram_mem[100710] = 16'b0000000000000000;
	sram_mem[100711] = 16'b0000000000000000;
	sram_mem[100712] = 16'b0000000000000000;
	sram_mem[100713] = 16'b0000000000000000;
	sram_mem[100714] = 16'b0000000000000000;
	sram_mem[100715] = 16'b0000000000000000;
	sram_mem[100716] = 16'b0000000000000000;
	sram_mem[100717] = 16'b0000000000000000;
	sram_mem[100718] = 16'b0000000000000000;
	sram_mem[100719] = 16'b0000000000000000;
	sram_mem[100720] = 16'b0000000000000000;
	sram_mem[100721] = 16'b0000000000000000;
	sram_mem[100722] = 16'b0000000000000000;
	sram_mem[100723] = 16'b0000000000000000;
	sram_mem[100724] = 16'b0000000000000000;
	sram_mem[100725] = 16'b0000000000000000;
	sram_mem[100726] = 16'b0000000000000000;
	sram_mem[100727] = 16'b0000000000000000;
	sram_mem[100728] = 16'b0000000000000000;
	sram_mem[100729] = 16'b0000000000000000;
	sram_mem[100730] = 16'b0000000000000000;
	sram_mem[100731] = 16'b0000000000000000;
	sram_mem[100732] = 16'b0000000000000000;
	sram_mem[100733] = 16'b0000000000000000;
	sram_mem[100734] = 16'b0000000000000000;
	sram_mem[100735] = 16'b0000000000000000;
	sram_mem[100736] = 16'b0000000000000000;
	sram_mem[100737] = 16'b0000000000000000;
	sram_mem[100738] = 16'b0000000000000000;
	sram_mem[100739] = 16'b0000000000000000;
	sram_mem[100740] = 16'b0000000000000000;
	sram_mem[100741] = 16'b0000000000000000;
	sram_mem[100742] = 16'b0000000000000000;
	sram_mem[100743] = 16'b0000000000000000;
	sram_mem[100744] = 16'b0000000000000000;
	sram_mem[100745] = 16'b0000000000000000;
	sram_mem[100746] = 16'b0000000000000000;
	sram_mem[100747] = 16'b0000000000000000;
	sram_mem[100748] = 16'b0000000000000000;
	sram_mem[100749] = 16'b0000000000000000;
	sram_mem[100750] = 16'b0000000000000000;
	sram_mem[100751] = 16'b0000000000000000;
	sram_mem[100752] = 16'b0000000000000000;
	sram_mem[100753] = 16'b0000000000000000;
	sram_mem[100754] = 16'b0000000000000000;
	sram_mem[100755] = 16'b0000000000000000;
	sram_mem[100756] = 16'b0000000000000000;
	sram_mem[100757] = 16'b0000000000000000;
	sram_mem[100758] = 16'b0000000000000000;
	sram_mem[100759] = 16'b0000000000000000;
	sram_mem[100760] = 16'b0000000000000000;
	sram_mem[100761] = 16'b0000000000000000;
	sram_mem[100762] = 16'b0000000000000000;
	sram_mem[100763] = 16'b0000000000000000;
	sram_mem[100764] = 16'b0000000000000000;
	sram_mem[100765] = 16'b0000000000000000;
	sram_mem[100766] = 16'b0000000000000000;
	sram_mem[100767] = 16'b0000000000000000;
	sram_mem[100768] = 16'b0000000000000000;
	sram_mem[100769] = 16'b0000000000000000;
	sram_mem[100770] = 16'b0000000000000000;
	sram_mem[100771] = 16'b0000000000000000;
	sram_mem[100772] = 16'b0000000000000000;
	sram_mem[100773] = 16'b0000000000000000;
	sram_mem[100774] = 16'b0000000000000000;
	sram_mem[100775] = 16'b0000000000000000;
	sram_mem[100776] = 16'b0000000000000000;
	sram_mem[100777] = 16'b0000000000000000;
	sram_mem[100778] = 16'b0000000000000000;
	sram_mem[100779] = 16'b0000000000000000;
	sram_mem[100780] = 16'b0000000000000000;
	sram_mem[100781] = 16'b0000000000000000;
	sram_mem[100782] = 16'b0000000000000000;
	sram_mem[100783] = 16'b0000000000000000;
	sram_mem[100784] = 16'b0000000000000000;
	sram_mem[100785] = 16'b0000000000000000;
	sram_mem[100786] = 16'b0000000000000000;
	sram_mem[100787] = 16'b0000000000000000;
	sram_mem[100788] = 16'b0000000000000000;
	sram_mem[100789] = 16'b0000000000000000;
	sram_mem[100790] = 16'b0000000000000000;
	sram_mem[100791] = 16'b0000000000000000;
	sram_mem[100792] = 16'b0000000000000000;
	sram_mem[100793] = 16'b0000000000000000;
	sram_mem[100794] = 16'b0000000000000000;
	sram_mem[100795] = 16'b0000000000000000;
	sram_mem[100796] = 16'b0000000000000000;
	sram_mem[100797] = 16'b0000000000000000;
	sram_mem[100798] = 16'b0000000000000000;
	sram_mem[100799] = 16'b0000000000000000;
	sram_mem[100800] = 16'b0000000000000000;
	sram_mem[100801] = 16'b0000000000000000;
	sram_mem[100802] = 16'b0000000000000000;
	sram_mem[100803] = 16'b0000000000000000;
	sram_mem[100804] = 16'b0000000000000000;
	sram_mem[100805] = 16'b0000000000000000;
	sram_mem[100806] = 16'b0000000000000000;
	sram_mem[100807] = 16'b0000000000000000;
	sram_mem[100808] = 16'b0000000000000000;
	sram_mem[100809] = 16'b0000000000000000;
	sram_mem[100810] = 16'b0000000000000000;
	sram_mem[100811] = 16'b0000000000000000;
	sram_mem[100812] = 16'b0000000000000000;
	sram_mem[100813] = 16'b0000000000000000;
	sram_mem[100814] = 16'b0000000000000000;
	sram_mem[100815] = 16'b0000000000000000;
	sram_mem[100816] = 16'b0000000000000000;
	sram_mem[100817] = 16'b0000000000000000;
	sram_mem[100818] = 16'b0000000000000000;
	sram_mem[100819] = 16'b0000000000000000;
	sram_mem[100820] = 16'b0000000000000000;
	sram_mem[100821] = 16'b0000000000000000;
	sram_mem[100822] = 16'b0000000000000000;
	sram_mem[100823] = 16'b0000000000000000;
	sram_mem[100824] = 16'b0000000000000000;
	sram_mem[100825] = 16'b0000000000000000;
	sram_mem[100826] = 16'b0000000000000000;
	sram_mem[100827] = 16'b0000000000000000;
	sram_mem[100828] = 16'b0000000000000000;
	sram_mem[100829] = 16'b0000000000000000;
	sram_mem[100830] = 16'b0000000000000000;
	sram_mem[100831] = 16'b0000000000000000;
	sram_mem[100832] = 16'b0000000000000000;
	sram_mem[100833] = 16'b0000000000000000;
	sram_mem[100834] = 16'b0000000000000000;
	sram_mem[100835] = 16'b0000000000000000;
	sram_mem[100836] = 16'b0000000000000000;
	sram_mem[100837] = 16'b0000000000000000;
	sram_mem[100838] = 16'b0000000000000000;
	sram_mem[100839] = 16'b0000000000000000;
	sram_mem[100840] = 16'b0000000000000000;
	sram_mem[100841] = 16'b0000000000000000;
	sram_mem[100842] = 16'b0000000000000000;
	sram_mem[100843] = 16'b0000000000000000;
	sram_mem[100844] = 16'b0000000000000000;
	sram_mem[100845] = 16'b0000000000000000;
	sram_mem[100846] = 16'b0000000000000000;
	sram_mem[100847] = 16'b0000000000000000;
	sram_mem[100848] = 16'b0000000000000000;
	sram_mem[100849] = 16'b0000000000000000;
	sram_mem[100850] = 16'b0000000000000000;
	sram_mem[100851] = 16'b0000000000000000;
	sram_mem[100852] = 16'b0000000000000000;
	sram_mem[100853] = 16'b0000000000000000;
	sram_mem[100854] = 16'b0000000000000000;
	sram_mem[100855] = 16'b0000000000000000;
	sram_mem[100856] = 16'b0000000000000000;
	sram_mem[100857] = 16'b0000000000000000;
	sram_mem[100858] = 16'b0000000000000000;
	sram_mem[100859] = 16'b0000000000000000;
	sram_mem[100860] = 16'b0000000000000000;
	sram_mem[100861] = 16'b0000000000000000;
	sram_mem[100862] = 16'b0000000000000000;
	sram_mem[100863] = 16'b0000000000000000;
	sram_mem[100864] = 16'b0000000000000000;
	sram_mem[100865] = 16'b0000000000000000;
	sram_mem[100866] = 16'b0000000000000000;
	sram_mem[100867] = 16'b0000000000000000;
	sram_mem[100868] = 16'b0000000000000000;
	sram_mem[100869] = 16'b0000000000000000;
	sram_mem[100870] = 16'b0000000000000000;
	sram_mem[100871] = 16'b0000000000000000;
	sram_mem[100872] = 16'b0000000000000000;
	sram_mem[100873] = 16'b0000000000000000;
	sram_mem[100874] = 16'b0000000000000000;
	sram_mem[100875] = 16'b0000000000000000;
	sram_mem[100876] = 16'b0000000000000000;
	sram_mem[100877] = 16'b0000000000000000;
	sram_mem[100878] = 16'b0000000000000000;
	sram_mem[100879] = 16'b0000000000000000;
	sram_mem[100880] = 16'b0000000000000000;
	sram_mem[100881] = 16'b0000000000000000;
	sram_mem[100882] = 16'b0000000000000000;
	sram_mem[100883] = 16'b0000000000000000;
	sram_mem[100884] = 16'b0000000000000000;
	sram_mem[100885] = 16'b0000000000000000;
	sram_mem[100886] = 16'b0000000000000000;
	sram_mem[100887] = 16'b0000000000000000;
	sram_mem[100888] = 16'b0000000000000000;
	sram_mem[100889] = 16'b0000000000000000;
	sram_mem[100890] = 16'b0000000000000000;
	sram_mem[100891] = 16'b0000000000000000;
	sram_mem[100892] = 16'b0000000000000000;
	sram_mem[100893] = 16'b0000000000000000;
	sram_mem[100894] = 16'b0000000000000000;
	sram_mem[100895] = 16'b0000000000000000;
	sram_mem[100896] = 16'b0000000000000000;
	sram_mem[100897] = 16'b0000000000000000;
	sram_mem[100898] = 16'b0000000000000000;
	sram_mem[100899] = 16'b0000000000000000;
	sram_mem[100900] = 16'b0000000000000000;
	sram_mem[100901] = 16'b0000000000000000;
	sram_mem[100902] = 16'b0000000000000000;
	sram_mem[100903] = 16'b0000000000000000;
	sram_mem[100904] = 16'b0000000000000000;
	sram_mem[100905] = 16'b0000000000000000;
	sram_mem[100906] = 16'b0000000000000000;
	sram_mem[100907] = 16'b0000000000000000;
	sram_mem[100908] = 16'b0000000000000000;
	sram_mem[100909] = 16'b0000000000000000;
	sram_mem[100910] = 16'b0000000000000000;
	sram_mem[100911] = 16'b0000000000000000;
	sram_mem[100912] = 16'b0000000000000000;
	sram_mem[100913] = 16'b0000000000000000;
	sram_mem[100914] = 16'b0000000000000000;
	sram_mem[100915] = 16'b0000000000000000;
	sram_mem[100916] = 16'b0000000000000000;
	sram_mem[100917] = 16'b0000000000000000;
	sram_mem[100918] = 16'b0000000000000000;
	sram_mem[100919] = 16'b0000000000000000;
	sram_mem[100920] = 16'b0000000000000000;
	sram_mem[100921] = 16'b0000000000000000;
	sram_mem[100922] = 16'b0000000000000000;
	sram_mem[100923] = 16'b0000000000000000;
	sram_mem[100924] = 16'b0000000000000000;
	sram_mem[100925] = 16'b0000000000000000;
	sram_mem[100926] = 16'b0000000000000000;
	sram_mem[100927] = 16'b0000000000000000;
	sram_mem[100928] = 16'b0000000000000000;
	sram_mem[100929] = 16'b0000000000000000;
	sram_mem[100930] = 16'b0000000000000000;
	sram_mem[100931] = 16'b0000000000000000;
	sram_mem[100932] = 16'b0000000000000000;
	sram_mem[100933] = 16'b0000000000000000;
	sram_mem[100934] = 16'b0000000000000000;
	sram_mem[100935] = 16'b0000000000000000;
	sram_mem[100936] = 16'b0000000000000000;
	sram_mem[100937] = 16'b0000000000000000;
	sram_mem[100938] = 16'b0000000000000000;
	sram_mem[100939] = 16'b0000000000000000;
	sram_mem[100940] = 16'b0000000000000000;
	sram_mem[100941] = 16'b0000000000000000;
	sram_mem[100942] = 16'b0000000000000000;
	sram_mem[100943] = 16'b0000000000000000;
	sram_mem[100944] = 16'b0000000000000000;
	sram_mem[100945] = 16'b0000000000000000;
	sram_mem[100946] = 16'b0000000000000000;
	sram_mem[100947] = 16'b0000000000000000;
	sram_mem[100948] = 16'b0000000000000000;
	sram_mem[100949] = 16'b0000000000000000;
	sram_mem[100950] = 16'b0000000000000000;
	sram_mem[100951] = 16'b0000000000000000;
	sram_mem[100952] = 16'b0000000000000000;
	sram_mem[100953] = 16'b0000000000000000;
	sram_mem[100954] = 16'b0000000000000000;
	sram_mem[100955] = 16'b0000000000000000;
	sram_mem[100956] = 16'b0000000000000000;
	sram_mem[100957] = 16'b0000000000000000;
	sram_mem[100958] = 16'b0000000000000000;
	sram_mem[100959] = 16'b0000000000000000;
	sram_mem[100960] = 16'b0000000000000000;
	sram_mem[100961] = 16'b0000000000000000;
	sram_mem[100962] = 16'b0000000000000000;
	sram_mem[100963] = 16'b0000000000000000;
	sram_mem[100964] = 16'b0000000000000000;
	sram_mem[100965] = 16'b0000000000000000;
	sram_mem[100966] = 16'b0000000000000000;
	sram_mem[100967] = 16'b0000000000000000;
	sram_mem[100968] = 16'b0000000000000000;
	sram_mem[100969] = 16'b0000000000000000;
	sram_mem[100970] = 16'b0000000000000000;
	sram_mem[100971] = 16'b0000000000000000;
	sram_mem[100972] = 16'b0000000000000000;
	sram_mem[100973] = 16'b0000000000000000;
	sram_mem[100974] = 16'b0000000000000000;
	sram_mem[100975] = 16'b0000000000000000;
	sram_mem[100976] = 16'b0000000000000000;
	sram_mem[100977] = 16'b0000000000000000;
	sram_mem[100978] = 16'b0000000000000000;
	sram_mem[100979] = 16'b0000000000000000;
	sram_mem[100980] = 16'b0000000000000000;
	sram_mem[100981] = 16'b0000000000000000;
	sram_mem[100982] = 16'b0000000000000000;
	sram_mem[100983] = 16'b0000000000000000;
	sram_mem[100984] = 16'b0000000000000000;
	sram_mem[100985] = 16'b0000000000000000;
	sram_mem[100986] = 16'b0000000000000000;
	sram_mem[100987] = 16'b0000000000000000;
	sram_mem[100988] = 16'b0000000000000000;
	sram_mem[100989] = 16'b0000000000000000;
	sram_mem[100990] = 16'b0000000000000000;
	sram_mem[100991] = 16'b0000000000000000;
	sram_mem[100992] = 16'b0000000000000000;
	sram_mem[100993] = 16'b0000000000000000;
	sram_mem[100994] = 16'b0000000000000000;
	sram_mem[100995] = 16'b0000000000000000;
	sram_mem[100996] = 16'b0000000000000000;
	sram_mem[100997] = 16'b0000000000000000;
	sram_mem[100998] = 16'b0000000000000000;
	sram_mem[100999] = 16'b0000000000000000;
	sram_mem[101000] = 16'b0000000000000000;
	sram_mem[101001] = 16'b0000000000000000;
	sram_mem[101002] = 16'b0000000000000000;
	sram_mem[101003] = 16'b0000000000000000;
	sram_mem[101004] = 16'b0000000000000000;
	sram_mem[101005] = 16'b0000000000000000;
	sram_mem[101006] = 16'b0000000000000000;
	sram_mem[101007] = 16'b0000000000000000;
	sram_mem[101008] = 16'b0000000000000000;
	sram_mem[101009] = 16'b0000000000000000;
	sram_mem[101010] = 16'b0000000000000000;
	sram_mem[101011] = 16'b0000000000000000;
	sram_mem[101012] = 16'b0000000000000000;
	sram_mem[101013] = 16'b0000000000000000;
	sram_mem[101014] = 16'b0000000000000000;
	sram_mem[101015] = 16'b0000000000000000;
	sram_mem[101016] = 16'b0000000000000000;
	sram_mem[101017] = 16'b0000000000000000;
	sram_mem[101018] = 16'b0000000000000000;
	sram_mem[101019] = 16'b0000000000000000;
	sram_mem[101020] = 16'b0000000000000000;
	sram_mem[101021] = 16'b0000000000000000;
	sram_mem[101022] = 16'b0000000000000000;
	sram_mem[101023] = 16'b0000000000000000;
	sram_mem[101024] = 16'b0000000000000000;
	sram_mem[101025] = 16'b0000000000000000;
	sram_mem[101026] = 16'b0000000000000000;
	sram_mem[101027] = 16'b0000000000000000;
	sram_mem[101028] = 16'b0000000000000000;
	sram_mem[101029] = 16'b0000000000000000;
	sram_mem[101030] = 16'b0000000000000000;
	sram_mem[101031] = 16'b0000000000000000;
	sram_mem[101032] = 16'b0000000000000000;
	sram_mem[101033] = 16'b0000000000000000;
	sram_mem[101034] = 16'b0000000000000000;
	sram_mem[101035] = 16'b0000000000000000;
	sram_mem[101036] = 16'b0000000000000000;
	sram_mem[101037] = 16'b0000000000000000;
	sram_mem[101038] = 16'b0000000000000000;
	sram_mem[101039] = 16'b0000000000000000;
	sram_mem[101040] = 16'b0000000000000000;
	sram_mem[101041] = 16'b0000000000000000;
	sram_mem[101042] = 16'b0000000000000000;
	sram_mem[101043] = 16'b0000000000000000;
	sram_mem[101044] = 16'b0000000000000000;
	sram_mem[101045] = 16'b0000000000000000;
	sram_mem[101046] = 16'b0000000000000000;
	sram_mem[101047] = 16'b0000000000000000;
	sram_mem[101048] = 16'b0000000000000000;
	sram_mem[101049] = 16'b0000000000000000;
	sram_mem[101050] = 16'b0000000000000000;
	sram_mem[101051] = 16'b0000000000000000;
	sram_mem[101052] = 16'b0000000000000000;
	sram_mem[101053] = 16'b0000000000000000;
	sram_mem[101054] = 16'b0000000000000000;
	sram_mem[101055] = 16'b0000000000000000;
	sram_mem[101056] = 16'b0000000000000000;
	sram_mem[101057] = 16'b0000000000000000;
	sram_mem[101058] = 16'b0000000000000000;
	sram_mem[101059] = 16'b0000000000000000;
	sram_mem[101060] = 16'b0000000000000000;
	sram_mem[101061] = 16'b0000000000000000;
	sram_mem[101062] = 16'b0000000000000000;
	sram_mem[101063] = 16'b0000000000000000;
	sram_mem[101064] = 16'b0000000000000000;
	sram_mem[101065] = 16'b0000000000000000;
	sram_mem[101066] = 16'b0000000000000000;
	sram_mem[101067] = 16'b0000000000000000;
	sram_mem[101068] = 16'b0000000000000000;
	sram_mem[101069] = 16'b0000000000000000;
	sram_mem[101070] = 16'b0000000000000000;
	sram_mem[101071] = 16'b0000000000000000;
	sram_mem[101072] = 16'b0000000000000000;
	sram_mem[101073] = 16'b0000000000000000;
	sram_mem[101074] = 16'b0000000000000000;
	sram_mem[101075] = 16'b0000000000000000;
	sram_mem[101076] = 16'b0000000000000000;
	sram_mem[101077] = 16'b0000000000000000;
	sram_mem[101078] = 16'b0000000000000000;
	sram_mem[101079] = 16'b0000000000000000;
	sram_mem[101080] = 16'b0000000000000000;
	sram_mem[101081] = 16'b0000000000000000;
	sram_mem[101082] = 16'b0000000000000000;
	sram_mem[101083] = 16'b0000000000000000;
	sram_mem[101084] = 16'b0000000000000000;
	sram_mem[101085] = 16'b0000000000000000;
	sram_mem[101086] = 16'b0000000000000000;
	sram_mem[101087] = 16'b0000000000000000;
	sram_mem[101088] = 16'b0000000000000000;
	sram_mem[101089] = 16'b0000000000000000;
	sram_mem[101090] = 16'b0000000000000000;
	sram_mem[101091] = 16'b0000000000000000;
	sram_mem[101092] = 16'b0000000000000000;
	sram_mem[101093] = 16'b0000000000000000;
	sram_mem[101094] = 16'b0000000000000000;
	sram_mem[101095] = 16'b0000000000000000;
	sram_mem[101096] = 16'b0000000000000000;
	sram_mem[101097] = 16'b0000000000000000;
	sram_mem[101098] = 16'b0000000000000000;
	sram_mem[101099] = 16'b0000000000000000;
	sram_mem[101100] = 16'b0000000000000000;
	sram_mem[101101] = 16'b0000000000000000;
	sram_mem[101102] = 16'b0000000000000000;
	sram_mem[101103] = 16'b0000000000000000;
	sram_mem[101104] = 16'b0000000000000000;
	sram_mem[101105] = 16'b0000000000000000;
	sram_mem[101106] = 16'b0000000000000000;
	sram_mem[101107] = 16'b0000000000000000;
	sram_mem[101108] = 16'b0000000000000000;
	sram_mem[101109] = 16'b0000000000000000;
	sram_mem[101110] = 16'b0000000000000000;
	sram_mem[101111] = 16'b0000000000000000;
	sram_mem[101112] = 16'b0000000000000000;
	sram_mem[101113] = 16'b0000000000000000;
	sram_mem[101114] = 16'b0000000000000000;
	sram_mem[101115] = 16'b0000000000000000;
	sram_mem[101116] = 16'b0000000000000000;
	sram_mem[101117] = 16'b0000000000000000;
	sram_mem[101118] = 16'b0000000000000000;
	sram_mem[101119] = 16'b0000000000000000;
	sram_mem[101120] = 16'b0000000000000000;
	sram_mem[101121] = 16'b0000000000000000;
	sram_mem[101122] = 16'b0000000000000000;
	sram_mem[101123] = 16'b0000000000000000;
	sram_mem[101124] = 16'b0000000000000000;
	sram_mem[101125] = 16'b0000000000000000;
	sram_mem[101126] = 16'b0000000000000000;
	sram_mem[101127] = 16'b0000000000000000;
	sram_mem[101128] = 16'b0000000000000000;
	sram_mem[101129] = 16'b0000000000000000;
	sram_mem[101130] = 16'b0000000000000000;
	sram_mem[101131] = 16'b0000000000000000;
	sram_mem[101132] = 16'b0000000000000000;
	sram_mem[101133] = 16'b0000000000000000;
	sram_mem[101134] = 16'b0000000000000000;
	sram_mem[101135] = 16'b0000000000000000;
	sram_mem[101136] = 16'b0000000000000000;
	sram_mem[101137] = 16'b0000000000000000;
	sram_mem[101138] = 16'b0000000000000000;
	sram_mem[101139] = 16'b0000000000000000;
	sram_mem[101140] = 16'b0000000000000000;
	sram_mem[101141] = 16'b0000000000000000;
	sram_mem[101142] = 16'b0000000000000000;
	sram_mem[101143] = 16'b0000000000000000;
	sram_mem[101144] = 16'b0000000000000000;
	sram_mem[101145] = 16'b0000000000000000;
	sram_mem[101146] = 16'b0000000000000000;
	sram_mem[101147] = 16'b0000000000000000;
	sram_mem[101148] = 16'b0000000000000000;
	sram_mem[101149] = 16'b0000000000000000;
	sram_mem[101150] = 16'b0000000000000000;
	sram_mem[101151] = 16'b0000000000000000;
	sram_mem[101152] = 16'b0000000000000000;
	sram_mem[101153] = 16'b0000000000000000;
	sram_mem[101154] = 16'b0000000000000000;
	sram_mem[101155] = 16'b0000000000000000;
	sram_mem[101156] = 16'b0000000000000000;
	sram_mem[101157] = 16'b0000000000000000;
	sram_mem[101158] = 16'b0000000000000000;
	sram_mem[101159] = 16'b0000000000000000;
	sram_mem[101160] = 16'b0000000000000000;
	sram_mem[101161] = 16'b0000000000000000;
	sram_mem[101162] = 16'b0000000000000000;
	sram_mem[101163] = 16'b0000000000000000;
	sram_mem[101164] = 16'b0000000000000000;
	sram_mem[101165] = 16'b0000000000000000;
	sram_mem[101166] = 16'b0000000000000000;
	sram_mem[101167] = 16'b0000000000000000;
	sram_mem[101168] = 16'b0000000000000000;
	sram_mem[101169] = 16'b0000000000000000;
	sram_mem[101170] = 16'b0000000000000000;
	sram_mem[101171] = 16'b0000000000000000;
	sram_mem[101172] = 16'b0000000000000000;
	sram_mem[101173] = 16'b0000000000000000;
	sram_mem[101174] = 16'b0000000000000000;
	sram_mem[101175] = 16'b0000000000000000;
	sram_mem[101176] = 16'b0000000000000000;
	sram_mem[101177] = 16'b0000000000000000;
	sram_mem[101178] = 16'b0000000000000000;
	sram_mem[101179] = 16'b0000000000000000;
	sram_mem[101180] = 16'b0000000000000000;
	sram_mem[101181] = 16'b0000000000000000;
	sram_mem[101182] = 16'b0000000000000000;
	sram_mem[101183] = 16'b0000000000000000;
	sram_mem[101184] = 16'b0000000000000000;
	sram_mem[101185] = 16'b0000000000000000;
	sram_mem[101186] = 16'b0000000000000000;
	sram_mem[101187] = 16'b0000000000000000;
	sram_mem[101188] = 16'b0000000000000000;
	sram_mem[101189] = 16'b0000000000000000;
	sram_mem[101190] = 16'b0000000000000000;
	sram_mem[101191] = 16'b0000000000000000;
	sram_mem[101192] = 16'b0000000000000000;
	sram_mem[101193] = 16'b0000000000000000;
	sram_mem[101194] = 16'b0000000000000000;
	sram_mem[101195] = 16'b0000000000000000;
	sram_mem[101196] = 16'b0000000000000000;
	sram_mem[101197] = 16'b0000000000000000;
	sram_mem[101198] = 16'b0000000000000000;
	sram_mem[101199] = 16'b0000000000000000;
	sram_mem[101200] = 16'b0000000000000000;
	sram_mem[101201] = 16'b0000000000000000;
	sram_mem[101202] = 16'b0000000000000000;
	sram_mem[101203] = 16'b0000000000000000;
	sram_mem[101204] = 16'b0000000000000000;
	sram_mem[101205] = 16'b0000000000000000;
	sram_mem[101206] = 16'b0000000000000000;
	sram_mem[101207] = 16'b0000000000000000;
	sram_mem[101208] = 16'b0000000000000000;
	sram_mem[101209] = 16'b0000000000000000;
	sram_mem[101210] = 16'b0000000000000000;
	sram_mem[101211] = 16'b0000000000000000;
	sram_mem[101212] = 16'b0000000000000000;
	sram_mem[101213] = 16'b0000000000000000;
	sram_mem[101214] = 16'b0000000000000000;
	sram_mem[101215] = 16'b0000000000000000;
	sram_mem[101216] = 16'b0000000000000000;
	sram_mem[101217] = 16'b0000000000000000;
	sram_mem[101218] = 16'b0000000000000000;
	sram_mem[101219] = 16'b0000000000000000;
	sram_mem[101220] = 16'b0000000000000000;
	sram_mem[101221] = 16'b0000000000000000;
	sram_mem[101222] = 16'b0000000000000000;
	sram_mem[101223] = 16'b0000000000000000;
	sram_mem[101224] = 16'b0000000000000000;
	sram_mem[101225] = 16'b0000000000000000;
	sram_mem[101226] = 16'b0000000000000000;
	sram_mem[101227] = 16'b0000000000000000;
	sram_mem[101228] = 16'b0000000000000000;
	sram_mem[101229] = 16'b0000000000000000;
	sram_mem[101230] = 16'b0000000000000000;
	sram_mem[101231] = 16'b0000000000000000;
	sram_mem[101232] = 16'b0000000000000000;
	sram_mem[101233] = 16'b0000000000000000;
	sram_mem[101234] = 16'b0000000000000000;
	sram_mem[101235] = 16'b0000000000000000;
	sram_mem[101236] = 16'b0000000000000000;
	sram_mem[101237] = 16'b0000000000000000;
	sram_mem[101238] = 16'b0000000000000000;
	sram_mem[101239] = 16'b0000000000000000;
	sram_mem[101240] = 16'b0000000000000000;
	sram_mem[101241] = 16'b0000000000000000;
	sram_mem[101242] = 16'b0000000000000000;
	sram_mem[101243] = 16'b0000000000000000;
	sram_mem[101244] = 16'b0000000000000000;
	sram_mem[101245] = 16'b0000000000000000;
	sram_mem[101246] = 16'b0000000000000000;
	sram_mem[101247] = 16'b0000000000000000;
	sram_mem[101248] = 16'b0000000000000000;
	sram_mem[101249] = 16'b0000000000000000;
	sram_mem[101250] = 16'b0000000000000000;
	sram_mem[101251] = 16'b0000000000000000;
	sram_mem[101252] = 16'b0000000000000000;
	sram_mem[101253] = 16'b0000000000000000;
	sram_mem[101254] = 16'b0000000000000000;
	sram_mem[101255] = 16'b0000000000000000;
	sram_mem[101256] = 16'b0000000000000000;
	sram_mem[101257] = 16'b0000000000000000;
	sram_mem[101258] = 16'b0000000000000000;
	sram_mem[101259] = 16'b0000000000000000;
	sram_mem[101260] = 16'b0000000000000000;
	sram_mem[101261] = 16'b0000000000000000;
	sram_mem[101262] = 16'b0000000000000000;
	sram_mem[101263] = 16'b0000000000000000;
	sram_mem[101264] = 16'b0000000000000000;
	sram_mem[101265] = 16'b0000000000000000;
	sram_mem[101266] = 16'b0000000000000000;
	sram_mem[101267] = 16'b0000000000000000;
	sram_mem[101268] = 16'b0000000000000000;
	sram_mem[101269] = 16'b0000000000000000;
	sram_mem[101270] = 16'b0000000000000000;
	sram_mem[101271] = 16'b0000000000000000;
	sram_mem[101272] = 16'b0000000000000000;
	sram_mem[101273] = 16'b0000000000000000;
	sram_mem[101274] = 16'b0000000000000000;
	sram_mem[101275] = 16'b0000000000000000;
	sram_mem[101276] = 16'b0000000000000000;
	sram_mem[101277] = 16'b0000000000000000;
	sram_mem[101278] = 16'b0000000000000000;
	sram_mem[101279] = 16'b0000000000000000;
	sram_mem[101280] = 16'b0000000000000000;
	sram_mem[101281] = 16'b0000000000000000;
	sram_mem[101282] = 16'b0000000000000000;
	sram_mem[101283] = 16'b0000000000000000;
	sram_mem[101284] = 16'b0000000000000000;
	sram_mem[101285] = 16'b0000000000000000;
	sram_mem[101286] = 16'b0000000000000000;
	sram_mem[101287] = 16'b0000000000000000;
	sram_mem[101288] = 16'b0000000000000000;
	sram_mem[101289] = 16'b0000000000000000;
	sram_mem[101290] = 16'b0000000000000000;
	sram_mem[101291] = 16'b0000000000000000;
	sram_mem[101292] = 16'b0000000000000000;
	sram_mem[101293] = 16'b0000000000000000;
	sram_mem[101294] = 16'b0000000000000000;
	sram_mem[101295] = 16'b0000000000000000;
	sram_mem[101296] = 16'b0000000000000000;
	sram_mem[101297] = 16'b0000000000000000;
	sram_mem[101298] = 16'b0000000000000000;
	sram_mem[101299] = 16'b0000000000000000;
	sram_mem[101300] = 16'b0000000000000000;
	sram_mem[101301] = 16'b0000000000000000;
	sram_mem[101302] = 16'b0000000000000000;
	sram_mem[101303] = 16'b0000000000000000;
	sram_mem[101304] = 16'b0000000000000000;
	sram_mem[101305] = 16'b0000000000000000;
	sram_mem[101306] = 16'b0000000000000000;
	sram_mem[101307] = 16'b0000000000000000;
	sram_mem[101308] = 16'b0000000000000000;
	sram_mem[101309] = 16'b0000000000000000;
	sram_mem[101310] = 16'b0000000000000000;
	sram_mem[101311] = 16'b0000000000000000;
	sram_mem[101312] = 16'b0000000000000000;
	sram_mem[101313] = 16'b0000000000000000;
	sram_mem[101314] = 16'b0000000000000000;
	sram_mem[101315] = 16'b0000000000000000;
	sram_mem[101316] = 16'b0000000000000000;
	sram_mem[101317] = 16'b0000000000000000;
	sram_mem[101318] = 16'b0000000000000000;
	sram_mem[101319] = 16'b0000000000000000;
	sram_mem[101320] = 16'b0000000000000000;
	sram_mem[101321] = 16'b0000000000000000;
	sram_mem[101322] = 16'b0000000000000000;
	sram_mem[101323] = 16'b0000000000000000;
	sram_mem[101324] = 16'b0000000000000000;
	sram_mem[101325] = 16'b0000000000000000;
	sram_mem[101326] = 16'b0000000000000000;
	sram_mem[101327] = 16'b0000000000000000;
	sram_mem[101328] = 16'b0000000000000000;
	sram_mem[101329] = 16'b0000000000000000;
	sram_mem[101330] = 16'b0000000000000000;
	sram_mem[101331] = 16'b0000000000000000;
	sram_mem[101332] = 16'b0000000000000000;
	sram_mem[101333] = 16'b0000000000000000;
	sram_mem[101334] = 16'b0000000000000000;
	sram_mem[101335] = 16'b0000000000000000;
	sram_mem[101336] = 16'b0000000000000000;
	sram_mem[101337] = 16'b0000000000000000;
	sram_mem[101338] = 16'b0000000000000000;
	sram_mem[101339] = 16'b0000000000000000;
	sram_mem[101340] = 16'b0000000000000000;
	sram_mem[101341] = 16'b0000000000000000;
	sram_mem[101342] = 16'b0000000000000000;
	sram_mem[101343] = 16'b0000000000000000;
	sram_mem[101344] = 16'b0000000000000000;
	sram_mem[101345] = 16'b0000000000000000;
	sram_mem[101346] = 16'b0000000000000000;
	sram_mem[101347] = 16'b0000000000000000;
	sram_mem[101348] = 16'b0000000000000000;
	sram_mem[101349] = 16'b0000000000000000;
	sram_mem[101350] = 16'b0000000000000000;
	sram_mem[101351] = 16'b0000000000000000;
	sram_mem[101352] = 16'b0000000000000000;
	sram_mem[101353] = 16'b0000000000000000;
	sram_mem[101354] = 16'b0000000000000000;
	sram_mem[101355] = 16'b0000000000000000;
	sram_mem[101356] = 16'b0000000000000000;
	sram_mem[101357] = 16'b0000000000000000;
	sram_mem[101358] = 16'b0000000000000000;
	sram_mem[101359] = 16'b0000000000000000;
	sram_mem[101360] = 16'b0000000000000000;
	sram_mem[101361] = 16'b0000000000000000;
	sram_mem[101362] = 16'b0000000000000000;
	sram_mem[101363] = 16'b0000000000000000;
	sram_mem[101364] = 16'b0000000000000000;
	sram_mem[101365] = 16'b0000000000000000;
	sram_mem[101366] = 16'b0000000000000000;
	sram_mem[101367] = 16'b0000000000000000;
	sram_mem[101368] = 16'b0000000000000000;
	sram_mem[101369] = 16'b0000000000000000;
	sram_mem[101370] = 16'b0000000000000000;
	sram_mem[101371] = 16'b0000000000000000;
	sram_mem[101372] = 16'b0000000000000000;
	sram_mem[101373] = 16'b0000000000000000;
	sram_mem[101374] = 16'b0000000000000000;
	sram_mem[101375] = 16'b0000000000000000;
	sram_mem[101376] = 16'b0000000000000000;
	sram_mem[101377] = 16'b0000000000000000;
	sram_mem[101378] = 16'b0000000000000000;
	sram_mem[101379] = 16'b0000000000000000;
	sram_mem[101380] = 16'b0000000000000000;
	sram_mem[101381] = 16'b0000000000000000;
	sram_mem[101382] = 16'b0000000000000000;
	sram_mem[101383] = 16'b0000000000000000;
	sram_mem[101384] = 16'b0000000000000000;
	sram_mem[101385] = 16'b0000000000000000;
	sram_mem[101386] = 16'b0000000000000000;
	sram_mem[101387] = 16'b0000000000000000;
	sram_mem[101388] = 16'b0000000000000000;
	sram_mem[101389] = 16'b0000000000000000;
	sram_mem[101390] = 16'b0000000000000000;
	sram_mem[101391] = 16'b0000000000000000;
	sram_mem[101392] = 16'b0000000000000000;
	sram_mem[101393] = 16'b0000000000000000;
	sram_mem[101394] = 16'b0000000000000000;
	sram_mem[101395] = 16'b0000000000000000;
	sram_mem[101396] = 16'b0000000000000000;
	sram_mem[101397] = 16'b0000000000000000;
	sram_mem[101398] = 16'b0000000000000000;
	sram_mem[101399] = 16'b0000000000000000;
	sram_mem[101400] = 16'b0000000000000000;
	sram_mem[101401] = 16'b0000000000000000;
	sram_mem[101402] = 16'b0000000000000000;
	sram_mem[101403] = 16'b0000000000000000;
	sram_mem[101404] = 16'b0000000000000000;
	sram_mem[101405] = 16'b0000000000000000;
	sram_mem[101406] = 16'b0000000000000000;
	sram_mem[101407] = 16'b0000000000000000;
	sram_mem[101408] = 16'b0000000000000000;
	sram_mem[101409] = 16'b0000000000000000;
	sram_mem[101410] = 16'b0000000000000000;
	sram_mem[101411] = 16'b0000000000000000;
	sram_mem[101412] = 16'b0000000000000000;
	sram_mem[101413] = 16'b0000000000000000;
	sram_mem[101414] = 16'b0000000000000000;
	sram_mem[101415] = 16'b0000000000000000;
	sram_mem[101416] = 16'b0000000000000000;
	sram_mem[101417] = 16'b0000000000000000;
	sram_mem[101418] = 16'b0000000000000000;
	sram_mem[101419] = 16'b0000000000000000;
	sram_mem[101420] = 16'b0000000000000000;
	sram_mem[101421] = 16'b0000000000000000;
	sram_mem[101422] = 16'b0000000000000000;
	sram_mem[101423] = 16'b0000000000000000;
	sram_mem[101424] = 16'b0000000000000000;
	sram_mem[101425] = 16'b0000000000000000;
	sram_mem[101426] = 16'b0000000000000000;
	sram_mem[101427] = 16'b0000000000000000;
	sram_mem[101428] = 16'b0000000000000000;
	sram_mem[101429] = 16'b0000000000000000;
	sram_mem[101430] = 16'b0000000000000000;
	sram_mem[101431] = 16'b0000000000000000;
	sram_mem[101432] = 16'b0000000000000000;
	sram_mem[101433] = 16'b0000000000000000;
	sram_mem[101434] = 16'b0000000000000000;
	sram_mem[101435] = 16'b0000000000000000;
	sram_mem[101436] = 16'b0000000000000000;
	sram_mem[101437] = 16'b0000000000000000;
	sram_mem[101438] = 16'b0000000000000000;
	sram_mem[101439] = 16'b0000000000000000;
	sram_mem[101440] = 16'b0000000000000000;
	sram_mem[101441] = 16'b0000000000000000;
	sram_mem[101442] = 16'b0000000000000000;
	sram_mem[101443] = 16'b0000000000000000;
	sram_mem[101444] = 16'b0000000000000000;
	sram_mem[101445] = 16'b0000000000000000;
	sram_mem[101446] = 16'b0000000000000000;
	sram_mem[101447] = 16'b0000000000000000;
	sram_mem[101448] = 16'b0000000000000000;
	sram_mem[101449] = 16'b0000000000000000;
	sram_mem[101450] = 16'b0000000000000000;
	sram_mem[101451] = 16'b0000000000000000;
	sram_mem[101452] = 16'b0000000000000000;
	sram_mem[101453] = 16'b0000000000000000;
	sram_mem[101454] = 16'b0000000000000000;
	sram_mem[101455] = 16'b0000000000000000;
	sram_mem[101456] = 16'b0000000000000000;
	sram_mem[101457] = 16'b0000000000000000;
	sram_mem[101458] = 16'b0000000000000000;
	sram_mem[101459] = 16'b0000000000000000;
	sram_mem[101460] = 16'b0000000000000000;
	sram_mem[101461] = 16'b0000000000000000;
	sram_mem[101462] = 16'b0000000000000000;
	sram_mem[101463] = 16'b0000000000000000;
	sram_mem[101464] = 16'b0000000000000000;
	sram_mem[101465] = 16'b0000000000000000;
	sram_mem[101466] = 16'b0000000000000000;
	sram_mem[101467] = 16'b0000000000000000;
	sram_mem[101468] = 16'b0000000000000000;
	sram_mem[101469] = 16'b0000000000000000;
	sram_mem[101470] = 16'b0000000000000000;
	sram_mem[101471] = 16'b0000000000000000;
	sram_mem[101472] = 16'b0000000000000000;
	sram_mem[101473] = 16'b0000000000000000;
	sram_mem[101474] = 16'b0000000000000000;
	sram_mem[101475] = 16'b0000000000000000;
	sram_mem[101476] = 16'b0000000000000000;
	sram_mem[101477] = 16'b0000000000000000;
	sram_mem[101478] = 16'b0000000000000000;
	sram_mem[101479] = 16'b0000000000000000;
	sram_mem[101480] = 16'b0000000000000000;
	sram_mem[101481] = 16'b0000000000000000;
	sram_mem[101482] = 16'b0000000000000000;
	sram_mem[101483] = 16'b0000000000000000;
	sram_mem[101484] = 16'b0000000000000000;
	sram_mem[101485] = 16'b0000000000000000;
	sram_mem[101486] = 16'b0000000000000000;
	sram_mem[101487] = 16'b0000000000000000;
	sram_mem[101488] = 16'b0000000000000000;
	sram_mem[101489] = 16'b0000000000000000;
	sram_mem[101490] = 16'b0000000000000000;
	sram_mem[101491] = 16'b0000000000000000;
	sram_mem[101492] = 16'b0000000000000000;
	sram_mem[101493] = 16'b0000000000000000;
	sram_mem[101494] = 16'b0000000000000000;
	sram_mem[101495] = 16'b0000000000000000;
	sram_mem[101496] = 16'b0000000000000000;
	sram_mem[101497] = 16'b0000000000000000;
	sram_mem[101498] = 16'b0000000000000000;
	sram_mem[101499] = 16'b0000000000000000;
	sram_mem[101500] = 16'b0000000000000000;
	sram_mem[101501] = 16'b0000000000000000;
	sram_mem[101502] = 16'b0000000000000000;
	sram_mem[101503] = 16'b0000000000000000;
	sram_mem[101504] = 16'b0000000000000000;
	sram_mem[101505] = 16'b0000000000000000;
	sram_mem[101506] = 16'b0000000000000000;
	sram_mem[101507] = 16'b0000000000000000;
	sram_mem[101508] = 16'b0000000000000000;
	sram_mem[101509] = 16'b0000000000000000;
	sram_mem[101510] = 16'b0000000000000000;
	sram_mem[101511] = 16'b0000000000000000;
	sram_mem[101512] = 16'b0000000000000000;
	sram_mem[101513] = 16'b0000000000000000;
	sram_mem[101514] = 16'b0000000000000000;
	sram_mem[101515] = 16'b0000000000000000;
	sram_mem[101516] = 16'b0000000000000000;
	sram_mem[101517] = 16'b0000000000000000;
	sram_mem[101518] = 16'b0000000000000000;
	sram_mem[101519] = 16'b0000000000000000;
	sram_mem[101520] = 16'b0000000000000000;
	sram_mem[101521] = 16'b0000000000000000;
	sram_mem[101522] = 16'b0000000000000000;
	sram_mem[101523] = 16'b0000000000000000;
	sram_mem[101524] = 16'b0000000000000000;
	sram_mem[101525] = 16'b0000000000000000;
	sram_mem[101526] = 16'b0000000000000000;
	sram_mem[101527] = 16'b0000000000000000;
	sram_mem[101528] = 16'b0000000000000000;
	sram_mem[101529] = 16'b0000000000000000;
	sram_mem[101530] = 16'b0000000000000000;
	sram_mem[101531] = 16'b0000000000000000;
	sram_mem[101532] = 16'b0000000000000000;
	sram_mem[101533] = 16'b0000000000000000;
	sram_mem[101534] = 16'b0000000000000000;
	sram_mem[101535] = 16'b0000000000000000;
	sram_mem[101536] = 16'b0000000000000000;
	sram_mem[101537] = 16'b0000000000000000;
	sram_mem[101538] = 16'b0000000000000000;
	sram_mem[101539] = 16'b0000000000000000;
	sram_mem[101540] = 16'b0000000000000000;
	sram_mem[101541] = 16'b0000000000000000;
	sram_mem[101542] = 16'b0000000000000000;
	sram_mem[101543] = 16'b0000000000000000;
	sram_mem[101544] = 16'b0000000000000000;
	sram_mem[101545] = 16'b0000000000000000;
	sram_mem[101546] = 16'b0000000000000000;
	sram_mem[101547] = 16'b0000000000000000;
	sram_mem[101548] = 16'b0000000000000000;
	sram_mem[101549] = 16'b0000000000000000;
	sram_mem[101550] = 16'b0000000000000000;
	sram_mem[101551] = 16'b0000000000000000;
	sram_mem[101552] = 16'b0000000000000000;
	sram_mem[101553] = 16'b0000000000000000;
	sram_mem[101554] = 16'b0000000000000000;
	sram_mem[101555] = 16'b0000000000000000;
	sram_mem[101556] = 16'b0000000000000000;
	sram_mem[101557] = 16'b0000000000000000;
	sram_mem[101558] = 16'b0000000000000000;
	sram_mem[101559] = 16'b0000000000000000;
	sram_mem[101560] = 16'b0000000000000000;
	sram_mem[101561] = 16'b0000000000000000;
	sram_mem[101562] = 16'b0000000000000000;
	sram_mem[101563] = 16'b0000000000000000;
	sram_mem[101564] = 16'b0000000000000000;
	sram_mem[101565] = 16'b0000000000000000;
	sram_mem[101566] = 16'b0000000000000000;
	sram_mem[101567] = 16'b0000000000000000;
	sram_mem[101568] = 16'b0000000000000000;
	sram_mem[101569] = 16'b0000000000000000;
	sram_mem[101570] = 16'b0000000000000000;
	sram_mem[101571] = 16'b0000000000000000;
	sram_mem[101572] = 16'b0000000000000000;
	sram_mem[101573] = 16'b0000000000000000;
	sram_mem[101574] = 16'b0000000000000000;
	sram_mem[101575] = 16'b0000000000000000;
	sram_mem[101576] = 16'b0000000000000000;
	sram_mem[101577] = 16'b0000000000000000;
	sram_mem[101578] = 16'b0000000000000000;
	sram_mem[101579] = 16'b0000000000000000;
	sram_mem[101580] = 16'b0000000000000000;
	sram_mem[101581] = 16'b0000000000000000;
	sram_mem[101582] = 16'b0000000000000000;
	sram_mem[101583] = 16'b0000000000000000;
	sram_mem[101584] = 16'b0000000000000000;
	sram_mem[101585] = 16'b0000000000000000;
	sram_mem[101586] = 16'b0000000000000000;
	sram_mem[101587] = 16'b0000000000000000;
	sram_mem[101588] = 16'b0000000000000000;
	sram_mem[101589] = 16'b0000000000000000;
	sram_mem[101590] = 16'b0000000000000000;
	sram_mem[101591] = 16'b0000000000000000;
	sram_mem[101592] = 16'b0000000000000000;
	sram_mem[101593] = 16'b0000000000000000;
	sram_mem[101594] = 16'b0000000000000000;
	sram_mem[101595] = 16'b0000000000000000;
	sram_mem[101596] = 16'b0000000000000000;
	sram_mem[101597] = 16'b0000000000000000;
	sram_mem[101598] = 16'b0000000000000000;
	sram_mem[101599] = 16'b0000000000000000;
	sram_mem[101600] = 16'b0000000000000000;
	sram_mem[101601] = 16'b0000000000000000;
	sram_mem[101602] = 16'b0000000000000000;
	sram_mem[101603] = 16'b0000000000000000;
	sram_mem[101604] = 16'b0000000000000000;
	sram_mem[101605] = 16'b0000000000000000;
	sram_mem[101606] = 16'b0000000000000000;
	sram_mem[101607] = 16'b0000000000000000;
	sram_mem[101608] = 16'b0000000000000000;
	sram_mem[101609] = 16'b0000000000000000;
	sram_mem[101610] = 16'b0000000000000000;
	sram_mem[101611] = 16'b0000000000000000;
	sram_mem[101612] = 16'b0000000000000000;
	sram_mem[101613] = 16'b0000000000000000;
	sram_mem[101614] = 16'b0000000000000000;
	sram_mem[101615] = 16'b0000000000000000;
	sram_mem[101616] = 16'b0000000000000000;
	sram_mem[101617] = 16'b0000000000000000;
	sram_mem[101618] = 16'b0000000000000000;
	sram_mem[101619] = 16'b0000000000000000;
	sram_mem[101620] = 16'b0000000000000000;
	sram_mem[101621] = 16'b0000000000000000;
	sram_mem[101622] = 16'b0000000000000000;
	sram_mem[101623] = 16'b0000000000000000;
	sram_mem[101624] = 16'b0000000000000000;
	sram_mem[101625] = 16'b0000000000000000;
	sram_mem[101626] = 16'b0000000000000000;
	sram_mem[101627] = 16'b0000000000000000;
	sram_mem[101628] = 16'b0000000000000000;
	sram_mem[101629] = 16'b0000000000000000;
	sram_mem[101630] = 16'b0000000000000000;
	sram_mem[101631] = 16'b0000000000000000;
	sram_mem[101632] = 16'b0000000000000000;
	sram_mem[101633] = 16'b0000000000000000;
	sram_mem[101634] = 16'b0000000000000000;
	sram_mem[101635] = 16'b0000000000000000;
	sram_mem[101636] = 16'b0000000000000000;
	sram_mem[101637] = 16'b0000000000000000;
	sram_mem[101638] = 16'b0000000000000000;
	sram_mem[101639] = 16'b0000000000000000;
	sram_mem[101640] = 16'b0000000000000000;
	sram_mem[101641] = 16'b0000000000000000;
	sram_mem[101642] = 16'b0000000000000000;
	sram_mem[101643] = 16'b0000000000000000;
	sram_mem[101644] = 16'b0000000000000000;
	sram_mem[101645] = 16'b0000000000000000;
	sram_mem[101646] = 16'b0000000000000000;
	sram_mem[101647] = 16'b0000000000000000;
	sram_mem[101648] = 16'b0000000000000000;
	sram_mem[101649] = 16'b0000000000000000;
	sram_mem[101650] = 16'b0000000000000000;
	sram_mem[101651] = 16'b0000000000000000;
	sram_mem[101652] = 16'b0000000000000000;
	sram_mem[101653] = 16'b0000000000000000;
	sram_mem[101654] = 16'b0000000000000000;
	sram_mem[101655] = 16'b0000000000000000;
	sram_mem[101656] = 16'b0000000000000000;
	sram_mem[101657] = 16'b0000000000000000;
	sram_mem[101658] = 16'b0000000000000000;
	sram_mem[101659] = 16'b0000000000000000;
	sram_mem[101660] = 16'b0000000000000000;
	sram_mem[101661] = 16'b0000000000000000;
	sram_mem[101662] = 16'b0000000000000000;
	sram_mem[101663] = 16'b0000000000000000;
	sram_mem[101664] = 16'b0000000000000000;
	sram_mem[101665] = 16'b0000000000000000;
	sram_mem[101666] = 16'b0000000000000000;
	sram_mem[101667] = 16'b0000000000000000;
	sram_mem[101668] = 16'b0000000000000000;
	sram_mem[101669] = 16'b0000000000000000;
	sram_mem[101670] = 16'b0000000000000000;
	sram_mem[101671] = 16'b0000000000000000;
	sram_mem[101672] = 16'b0000000000000000;
	sram_mem[101673] = 16'b0000000000000000;
	sram_mem[101674] = 16'b0000000000000000;
	sram_mem[101675] = 16'b0000000000000000;
	sram_mem[101676] = 16'b0000000000000000;
	sram_mem[101677] = 16'b0000000000000000;
	sram_mem[101678] = 16'b0000000000000000;
	sram_mem[101679] = 16'b0000000000000000;
	sram_mem[101680] = 16'b0000000000000000;
	sram_mem[101681] = 16'b0000000000000000;
	sram_mem[101682] = 16'b0000000000000000;
	sram_mem[101683] = 16'b0000000000000000;
	sram_mem[101684] = 16'b0000000000000000;
	sram_mem[101685] = 16'b0000000000000000;
	sram_mem[101686] = 16'b0000000000000000;
	sram_mem[101687] = 16'b0000000000000000;
	sram_mem[101688] = 16'b0000000000000000;
	sram_mem[101689] = 16'b0000000000000000;
	sram_mem[101690] = 16'b0000000000000000;
	sram_mem[101691] = 16'b0000000000000000;
	sram_mem[101692] = 16'b0000000000000000;
	sram_mem[101693] = 16'b0000000000000000;
	sram_mem[101694] = 16'b0000000000000000;
	sram_mem[101695] = 16'b0000000000000000;
	sram_mem[101696] = 16'b0000000000000000;
	sram_mem[101697] = 16'b0000000000000000;
	sram_mem[101698] = 16'b0000000000000000;
	sram_mem[101699] = 16'b0000000000000000;
	sram_mem[101700] = 16'b0000000000000000;
	sram_mem[101701] = 16'b0000000000000000;
	sram_mem[101702] = 16'b0000000000000000;
	sram_mem[101703] = 16'b0000000000000000;
	sram_mem[101704] = 16'b0000000000000000;
	sram_mem[101705] = 16'b0000000000000000;
	sram_mem[101706] = 16'b0000000000000000;
	sram_mem[101707] = 16'b0000000000000000;
	sram_mem[101708] = 16'b0000000000000000;
	sram_mem[101709] = 16'b0000000000000000;
	sram_mem[101710] = 16'b0000000000000000;
	sram_mem[101711] = 16'b0000000000000000;
	sram_mem[101712] = 16'b0000000000000000;
	sram_mem[101713] = 16'b0000000000000000;
	sram_mem[101714] = 16'b0000000000000000;
	sram_mem[101715] = 16'b0000000000000000;
	sram_mem[101716] = 16'b0000000000000000;
	sram_mem[101717] = 16'b0000000000000000;
	sram_mem[101718] = 16'b0000000000000000;
	sram_mem[101719] = 16'b0000000000000000;
	sram_mem[101720] = 16'b0000000000000000;
	sram_mem[101721] = 16'b0000000000000000;
	sram_mem[101722] = 16'b0000000000000000;
	sram_mem[101723] = 16'b0000000000000000;
	sram_mem[101724] = 16'b0000000000000000;
	sram_mem[101725] = 16'b0000000000000000;
	sram_mem[101726] = 16'b0000000000000000;
	sram_mem[101727] = 16'b0000000000000000;
	sram_mem[101728] = 16'b0000000000000000;
	sram_mem[101729] = 16'b0000000000000000;
	sram_mem[101730] = 16'b0000000000000000;
	sram_mem[101731] = 16'b0000000000000000;
	sram_mem[101732] = 16'b0000000000000000;
	sram_mem[101733] = 16'b0000000000000000;
	sram_mem[101734] = 16'b0000000000000000;
	sram_mem[101735] = 16'b0000000000000000;
	sram_mem[101736] = 16'b0000000000000000;
	sram_mem[101737] = 16'b0000000000000000;
	sram_mem[101738] = 16'b0000000000000000;
	sram_mem[101739] = 16'b0000000000000000;
	sram_mem[101740] = 16'b0000000000000000;
	sram_mem[101741] = 16'b0000000000000000;
	sram_mem[101742] = 16'b0000000000000000;
	sram_mem[101743] = 16'b0000000000000000;
	sram_mem[101744] = 16'b0000000000000000;
	sram_mem[101745] = 16'b0000000000000000;
	sram_mem[101746] = 16'b0000000000000000;
	sram_mem[101747] = 16'b0000000000000000;
	sram_mem[101748] = 16'b0000000000000000;
	sram_mem[101749] = 16'b0000000000000000;
	sram_mem[101750] = 16'b0000000000000000;
	sram_mem[101751] = 16'b0000000000000000;
	sram_mem[101752] = 16'b0000000000000000;
	sram_mem[101753] = 16'b0000000000000000;
	sram_mem[101754] = 16'b0000000000000000;
	sram_mem[101755] = 16'b0000000000000000;
	sram_mem[101756] = 16'b0000000000000000;
	sram_mem[101757] = 16'b0000000000000000;
	sram_mem[101758] = 16'b0000000000000000;
	sram_mem[101759] = 16'b0000000000000000;
	sram_mem[101760] = 16'b0000000000000000;
	sram_mem[101761] = 16'b0000000000000000;
	sram_mem[101762] = 16'b0000000000000000;
	sram_mem[101763] = 16'b0000000000000000;
	sram_mem[101764] = 16'b0000000000000000;
	sram_mem[101765] = 16'b0000000000000000;
	sram_mem[101766] = 16'b0000000000000000;
	sram_mem[101767] = 16'b0000000000000000;
	sram_mem[101768] = 16'b0000000000000000;
	sram_mem[101769] = 16'b0000000000000000;
	sram_mem[101770] = 16'b0000000000000000;
	sram_mem[101771] = 16'b0000000000000000;
	sram_mem[101772] = 16'b0000000000000000;
	sram_mem[101773] = 16'b0000000000000000;
	sram_mem[101774] = 16'b0000000000000000;
	sram_mem[101775] = 16'b0000000000000000;
	sram_mem[101776] = 16'b0000000000000000;
	sram_mem[101777] = 16'b0000000000000000;
	sram_mem[101778] = 16'b0000000000000000;
	sram_mem[101779] = 16'b0000000000000000;
	sram_mem[101780] = 16'b0000000000000000;
	sram_mem[101781] = 16'b0000000000000000;
	sram_mem[101782] = 16'b0000000000000000;
	sram_mem[101783] = 16'b0000000000000000;
	sram_mem[101784] = 16'b0000000000000000;
	sram_mem[101785] = 16'b0000000000000000;
	sram_mem[101786] = 16'b0000000000000000;
	sram_mem[101787] = 16'b0000000000000000;
	sram_mem[101788] = 16'b0000000000000000;
	sram_mem[101789] = 16'b0000000000000000;
	sram_mem[101790] = 16'b0000000000000000;
	sram_mem[101791] = 16'b0000000000000000;
	sram_mem[101792] = 16'b0000000000000000;
	sram_mem[101793] = 16'b0000000000000000;
	sram_mem[101794] = 16'b0000000000000000;
	sram_mem[101795] = 16'b0000000000000000;
	sram_mem[101796] = 16'b0000000000000000;
	sram_mem[101797] = 16'b0000000000000000;
	sram_mem[101798] = 16'b0000000000000000;
	sram_mem[101799] = 16'b0000000000000000;
	sram_mem[101800] = 16'b0000000000000000;
	sram_mem[101801] = 16'b0000000000000000;
	sram_mem[101802] = 16'b0000000000000000;
	sram_mem[101803] = 16'b0000000000000000;
	sram_mem[101804] = 16'b0000000000000000;
	sram_mem[101805] = 16'b0000000000000000;
	sram_mem[101806] = 16'b0000000000000000;
	sram_mem[101807] = 16'b0000000000000000;
	sram_mem[101808] = 16'b0000000000000000;
	sram_mem[101809] = 16'b0000000000000000;
	sram_mem[101810] = 16'b0000000000000000;
	sram_mem[101811] = 16'b0000000000000000;
	sram_mem[101812] = 16'b0000000000000000;
	sram_mem[101813] = 16'b0000000000000000;
	sram_mem[101814] = 16'b0000000000000000;
	sram_mem[101815] = 16'b0000000000000000;
	sram_mem[101816] = 16'b0000000000000000;
	sram_mem[101817] = 16'b0000000000000000;
	sram_mem[101818] = 16'b0000000000000000;
	sram_mem[101819] = 16'b0000000000000000;
	sram_mem[101820] = 16'b0000000000000000;
	sram_mem[101821] = 16'b0000000000000000;
	sram_mem[101822] = 16'b0000000000000000;
	sram_mem[101823] = 16'b0000000000000000;
	sram_mem[101824] = 16'b0000000000000000;
	sram_mem[101825] = 16'b0000000000000000;
	sram_mem[101826] = 16'b0000000000000000;
	sram_mem[101827] = 16'b0000000000000000;
	sram_mem[101828] = 16'b0000000000000000;
	sram_mem[101829] = 16'b0000000000000000;
	sram_mem[101830] = 16'b0000000000000000;
	sram_mem[101831] = 16'b0000000000000000;
	sram_mem[101832] = 16'b0000000000000000;
	sram_mem[101833] = 16'b0000000000000000;
	sram_mem[101834] = 16'b0000000000000000;
	sram_mem[101835] = 16'b0000000000000000;
	sram_mem[101836] = 16'b0000000000000000;
	sram_mem[101837] = 16'b0000000000000000;
	sram_mem[101838] = 16'b0000000000000000;
	sram_mem[101839] = 16'b0000000000000000;
	sram_mem[101840] = 16'b0000000000000000;
	sram_mem[101841] = 16'b0000000000000000;
	sram_mem[101842] = 16'b0000000000000000;
	sram_mem[101843] = 16'b0000000000000000;
	sram_mem[101844] = 16'b0000000000000000;
	sram_mem[101845] = 16'b0000000000000000;
	sram_mem[101846] = 16'b0000000000000000;
	sram_mem[101847] = 16'b0000000000000000;
	sram_mem[101848] = 16'b0000000000000000;
	sram_mem[101849] = 16'b0000000000000000;
	sram_mem[101850] = 16'b0000000000000000;
	sram_mem[101851] = 16'b0000000000000000;
	sram_mem[101852] = 16'b0000000000000000;
	sram_mem[101853] = 16'b0000000000000000;
	sram_mem[101854] = 16'b0000000000000000;
	sram_mem[101855] = 16'b0000000000000000;
	sram_mem[101856] = 16'b0000000000000000;
	sram_mem[101857] = 16'b0000000000000000;
	sram_mem[101858] = 16'b0000000000000000;
	sram_mem[101859] = 16'b0000000000000000;
	sram_mem[101860] = 16'b0000000000000000;
	sram_mem[101861] = 16'b0000000000000000;
	sram_mem[101862] = 16'b0000000000000000;
	sram_mem[101863] = 16'b0000000000000000;
	sram_mem[101864] = 16'b0000000000000000;
	sram_mem[101865] = 16'b0000000000000000;
	sram_mem[101866] = 16'b0000000000000000;
	sram_mem[101867] = 16'b0000000000000000;
	sram_mem[101868] = 16'b0000000000000000;
	sram_mem[101869] = 16'b0000000000000000;
	sram_mem[101870] = 16'b0000000000000000;
	sram_mem[101871] = 16'b0000000000000000;
	sram_mem[101872] = 16'b0000000000000000;
	sram_mem[101873] = 16'b0000000000000000;
	sram_mem[101874] = 16'b0000000000000000;
	sram_mem[101875] = 16'b0000000000000000;
	sram_mem[101876] = 16'b0000000000000000;
	sram_mem[101877] = 16'b0000000000000000;
	sram_mem[101878] = 16'b0000000000000000;
	sram_mem[101879] = 16'b0000000000000000;
	sram_mem[101880] = 16'b0000000000000000;
	sram_mem[101881] = 16'b0000000000000000;
	sram_mem[101882] = 16'b0000000000000000;
	sram_mem[101883] = 16'b0000000000000000;
	sram_mem[101884] = 16'b0000000000000000;
	sram_mem[101885] = 16'b0000000000000000;
	sram_mem[101886] = 16'b0000000000000000;
	sram_mem[101887] = 16'b0000000000000000;
	sram_mem[101888] = 16'b0000000000000000;
	sram_mem[101889] = 16'b0000000000000000;
	sram_mem[101890] = 16'b0000000000000000;
	sram_mem[101891] = 16'b0000000000000000;
	sram_mem[101892] = 16'b0000000000000000;
	sram_mem[101893] = 16'b0000000000000000;
	sram_mem[101894] = 16'b0000000000000000;
	sram_mem[101895] = 16'b0000000000000000;
	sram_mem[101896] = 16'b0000000000000000;
	sram_mem[101897] = 16'b0000000000000000;
	sram_mem[101898] = 16'b0000000000000000;
	sram_mem[101899] = 16'b0000000000000000;
	sram_mem[101900] = 16'b0000000000000000;
	sram_mem[101901] = 16'b0000000000000000;
	sram_mem[101902] = 16'b0000000000000000;
	sram_mem[101903] = 16'b0000000000000000;
	sram_mem[101904] = 16'b0000000000000000;
	sram_mem[101905] = 16'b0000000000000000;
	sram_mem[101906] = 16'b0000000000000000;
	sram_mem[101907] = 16'b0000000000000000;
	sram_mem[101908] = 16'b0000000000000000;
	sram_mem[101909] = 16'b0000000000000000;
	sram_mem[101910] = 16'b0000000000000000;
	sram_mem[101911] = 16'b0000000000000000;
	sram_mem[101912] = 16'b0000000000000000;
	sram_mem[101913] = 16'b0000000000000000;
	sram_mem[101914] = 16'b0000000000000000;
	sram_mem[101915] = 16'b0000000000000000;
	sram_mem[101916] = 16'b0000000000000000;
	sram_mem[101917] = 16'b0000000000000000;
	sram_mem[101918] = 16'b0000000000000000;
	sram_mem[101919] = 16'b0000000000000000;
	sram_mem[101920] = 16'b0000000000000000;
	sram_mem[101921] = 16'b0000000000000000;
	sram_mem[101922] = 16'b0000000000000000;
	sram_mem[101923] = 16'b0000000000000000;
	sram_mem[101924] = 16'b0000000000000000;
	sram_mem[101925] = 16'b0000000000000000;
	sram_mem[101926] = 16'b0000000000000000;
	sram_mem[101927] = 16'b0000000000000000;
	sram_mem[101928] = 16'b0000000000000000;
	sram_mem[101929] = 16'b0000000000000000;
	sram_mem[101930] = 16'b0000000000000000;
	sram_mem[101931] = 16'b0000000000000000;
	sram_mem[101932] = 16'b0000000000000000;
	sram_mem[101933] = 16'b0000000000000000;
	sram_mem[101934] = 16'b0000000000000000;
	sram_mem[101935] = 16'b0000000000000000;
	sram_mem[101936] = 16'b0000000000000000;
	sram_mem[101937] = 16'b0000000000000000;
	sram_mem[101938] = 16'b0000000000000000;
	sram_mem[101939] = 16'b0000000000000000;
	sram_mem[101940] = 16'b0000000000000000;
	sram_mem[101941] = 16'b0000000000000000;
	sram_mem[101942] = 16'b0000000000000000;
	sram_mem[101943] = 16'b0000000000000000;
	sram_mem[101944] = 16'b0000000000000000;
	sram_mem[101945] = 16'b0000000000000000;
	sram_mem[101946] = 16'b0000000000000000;
	sram_mem[101947] = 16'b0000000000000000;
	sram_mem[101948] = 16'b0000000000000000;
	sram_mem[101949] = 16'b0000000000000000;
	sram_mem[101950] = 16'b0000000000000000;
	sram_mem[101951] = 16'b0000000000000000;
	sram_mem[101952] = 16'b0000000000000000;
	sram_mem[101953] = 16'b0000000000000000;
	sram_mem[101954] = 16'b0000000000000000;
	sram_mem[101955] = 16'b0000000000000000;
	sram_mem[101956] = 16'b0000000000000000;
	sram_mem[101957] = 16'b0000000000000000;
	sram_mem[101958] = 16'b0000000000000000;
	sram_mem[101959] = 16'b0000000000000000;
	sram_mem[101960] = 16'b0000000000000000;
	sram_mem[101961] = 16'b0000000000000000;
	sram_mem[101962] = 16'b0000000000000000;
	sram_mem[101963] = 16'b0000000000000000;
	sram_mem[101964] = 16'b0000000000000000;
	sram_mem[101965] = 16'b0000000000000000;
	sram_mem[101966] = 16'b0000000000000000;
	sram_mem[101967] = 16'b0000000000000000;
	sram_mem[101968] = 16'b0000000000000000;
	sram_mem[101969] = 16'b0000000000000000;
	sram_mem[101970] = 16'b0000000000000000;
	sram_mem[101971] = 16'b0000000000000000;
	sram_mem[101972] = 16'b0000000000000000;
	sram_mem[101973] = 16'b0000000000000000;
	sram_mem[101974] = 16'b0000000000000000;
	sram_mem[101975] = 16'b0000000000000000;
	sram_mem[101976] = 16'b0000000000000000;
	sram_mem[101977] = 16'b0000000000000000;
	sram_mem[101978] = 16'b0000000000000000;
	sram_mem[101979] = 16'b0000000000000000;
	sram_mem[101980] = 16'b0000000000000000;
	sram_mem[101981] = 16'b0000000000000000;
	sram_mem[101982] = 16'b0000000000000000;
	sram_mem[101983] = 16'b0000000000000000;
	sram_mem[101984] = 16'b0000000000000000;
	sram_mem[101985] = 16'b0000000000000000;
	sram_mem[101986] = 16'b0000000000000000;
	sram_mem[101987] = 16'b0000000000000000;
	sram_mem[101988] = 16'b0000000000000000;
	sram_mem[101989] = 16'b0000000000000000;
	sram_mem[101990] = 16'b0000000000000000;
	sram_mem[101991] = 16'b0000000000000000;
	sram_mem[101992] = 16'b0000000000000000;
	sram_mem[101993] = 16'b0000000000000000;
	sram_mem[101994] = 16'b0000000000000000;
	sram_mem[101995] = 16'b0000000000000000;
	sram_mem[101996] = 16'b0000000000000000;
	sram_mem[101997] = 16'b0000000000000000;
	sram_mem[101998] = 16'b0000000000000000;
	sram_mem[101999] = 16'b0000000000000000;
	sram_mem[102000] = 16'b0000000000000000;
	sram_mem[102001] = 16'b0000000000000000;
	sram_mem[102002] = 16'b0000000000000000;
	sram_mem[102003] = 16'b0000000000000000;
	sram_mem[102004] = 16'b0000000000000000;
	sram_mem[102005] = 16'b0000000000000000;
	sram_mem[102006] = 16'b0000000000000000;
	sram_mem[102007] = 16'b0000000000000000;
	sram_mem[102008] = 16'b0000000000000000;
	sram_mem[102009] = 16'b0000000000000000;
	sram_mem[102010] = 16'b0000000000000000;
	sram_mem[102011] = 16'b0000000000000000;
	sram_mem[102012] = 16'b0000000000000000;
	sram_mem[102013] = 16'b0000000000000000;
	sram_mem[102014] = 16'b0000000000000000;
	sram_mem[102015] = 16'b0000000000000000;
	sram_mem[102016] = 16'b0000000000000000;
	sram_mem[102017] = 16'b0000000000000000;
	sram_mem[102018] = 16'b0000000000000000;
	sram_mem[102019] = 16'b0000000000000000;
	sram_mem[102020] = 16'b0000000000000000;
	sram_mem[102021] = 16'b0000000000000000;
	sram_mem[102022] = 16'b0000000000000000;
	sram_mem[102023] = 16'b0000000000000000;
	sram_mem[102024] = 16'b0000000000000000;
	sram_mem[102025] = 16'b0000000000000000;
	sram_mem[102026] = 16'b0000000000000000;
	sram_mem[102027] = 16'b0000000000000000;
	sram_mem[102028] = 16'b0000000000000000;
	sram_mem[102029] = 16'b0000000000000000;
	sram_mem[102030] = 16'b0000000000000000;
	sram_mem[102031] = 16'b0000000000000000;
	sram_mem[102032] = 16'b0000000000000000;
	sram_mem[102033] = 16'b0000000000000000;
	sram_mem[102034] = 16'b0000000000000000;
	sram_mem[102035] = 16'b0000000000000000;
	sram_mem[102036] = 16'b0000000000000000;
	sram_mem[102037] = 16'b0000000000000000;
	sram_mem[102038] = 16'b0000000000000000;
	sram_mem[102039] = 16'b0000000000000000;
	sram_mem[102040] = 16'b0000000000000000;
	sram_mem[102041] = 16'b0000000000000000;
	sram_mem[102042] = 16'b0000000000000000;
	sram_mem[102043] = 16'b0000000000000000;
	sram_mem[102044] = 16'b0000000000000000;
	sram_mem[102045] = 16'b0000000000000000;
	sram_mem[102046] = 16'b0000000000000000;
	sram_mem[102047] = 16'b0000000000000000;
	sram_mem[102048] = 16'b0000000000000000;
	sram_mem[102049] = 16'b0000000000000000;
	sram_mem[102050] = 16'b0000000000000000;
	sram_mem[102051] = 16'b0000000000000000;
	sram_mem[102052] = 16'b0000000000000000;
	sram_mem[102053] = 16'b0000000000000000;
	sram_mem[102054] = 16'b0000000000000000;
	sram_mem[102055] = 16'b0000000000000000;
	sram_mem[102056] = 16'b0000000000000000;
	sram_mem[102057] = 16'b0000000000000000;
	sram_mem[102058] = 16'b0000000000000000;
	sram_mem[102059] = 16'b0000000000000000;
	sram_mem[102060] = 16'b0000000000000000;
	sram_mem[102061] = 16'b0000000000000000;
	sram_mem[102062] = 16'b0000000000000000;
	sram_mem[102063] = 16'b0000000000000000;
	sram_mem[102064] = 16'b0000000000000000;
	sram_mem[102065] = 16'b0000000000000000;
	sram_mem[102066] = 16'b0000000000000000;
	sram_mem[102067] = 16'b0000000000000000;
	sram_mem[102068] = 16'b0000000000000000;
	sram_mem[102069] = 16'b0000000000000000;
	sram_mem[102070] = 16'b0000000000000000;
	sram_mem[102071] = 16'b0000000000000000;
	sram_mem[102072] = 16'b0000000000000000;
	sram_mem[102073] = 16'b0000000000000000;
	sram_mem[102074] = 16'b0000000000000000;
	sram_mem[102075] = 16'b0000000000000000;
	sram_mem[102076] = 16'b0000000000000000;
	sram_mem[102077] = 16'b0000000000000000;
	sram_mem[102078] = 16'b0000000000000000;
	sram_mem[102079] = 16'b0000000000000000;
	sram_mem[102080] = 16'b0000000000000000;
	sram_mem[102081] = 16'b0000000000000000;
	sram_mem[102082] = 16'b0000000000000000;
	sram_mem[102083] = 16'b0000000000000000;
	sram_mem[102084] = 16'b0000000000000000;
	sram_mem[102085] = 16'b0000000000000000;
	sram_mem[102086] = 16'b0000000000000000;
	sram_mem[102087] = 16'b0000000000000000;
	sram_mem[102088] = 16'b0000000000000000;
	sram_mem[102089] = 16'b0000000000000000;
	sram_mem[102090] = 16'b0000000000000000;
	sram_mem[102091] = 16'b0000000000000000;
	sram_mem[102092] = 16'b0000000000000000;
	sram_mem[102093] = 16'b0000000000000000;
	sram_mem[102094] = 16'b0000000000000000;
	sram_mem[102095] = 16'b0000000000000000;
	sram_mem[102096] = 16'b0000000000000000;
	sram_mem[102097] = 16'b0000000000000000;
	sram_mem[102098] = 16'b0000000000000000;
	sram_mem[102099] = 16'b0000000000000000;
	sram_mem[102100] = 16'b0000000000000000;
	sram_mem[102101] = 16'b0000000000000000;
	sram_mem[102102] = 16'b0000000000000000;
	sram_mem[102103] = 16'b0000000000000000;
	sram_mem[102104] = 16'b0000000000000000;
	sram_mem[102105] = 16'b0000000000000000;
	sram_mem[102106] = 16'b0000000000000000;
	sram_mem[102107] = 16'b0000000000000000;
	sram_mem[102108] = 16'b0000000000000000;
	sram_mem[102109] = 16'b0000000000000000;
	sram_mem[102110] = 16'b0000000000000000;
	sram_mem[102111] = 16'b0000000000000000;
	sram_mem[102112] = 16'b0000000000000000;
	sram_mem[102113] = 16'b0000000000000000;
	sram_mem[102114] = 16'b0000000000000000;
	sram_mem[102115] = 16'b0000000000000000;
	sram_mem[102116] = 16'b0000000000000000;
	sram_mem[102117] = 16'b0000000000000000;
	sram_mem[102118] = 16'b0000000000000000;
	sram_mem[102119] = 16'b0000000000000000;
	sram_mem[102120] = 16'b0000000000000000;
	sram_mem[102121] = 16'b0000000000000000;
	sram_mem[102122] = 16'b0000000000000000;
	sram_mem[102123] = 16'b0000000000000000;
	sram_mem[102124] = 16'b0000000000000000;
	sram_mem[102125] = 16'b0000000000000000;
	sram_mem[102126] = 16'b0000000000000000;
	sram_mem[102127] = 16'b0000000000000000;
	sram_mem[102128] = 16'b0000000000000000;
	sram_mem[102129] = 16'b0000000000000000;
	sram_mem[102130] = 16'b0000000000000000;
	sram_mem[102131] = 16'b0000000000000000;
	sram_mem[102132] = 16'b0000000000000000;
	sram_mem[102133] = 16'b0000000000000000;
	sram_mem[102134] = 16'b0000000000000000;
	sram_mem[102135] = 16'b0000000000000000;
	sram_mem[102136] = 16'b0000000000000000;
	sram_mem[102137] = 16'b0000000000000000;
	sram_mem[102138] = 16'b0000000000000000;
	sram_mem[102139] = 16'b0000000000000000;
	sram_mem[102140] = 16'b0000000000000000;
	sram_mem[102141] = 16'b0000000000000000;
	sram_mem[102142] = 16'b0000000000000000;
	sram_mem[102143] = 16'b0000000000000000;
	sram_mem[102144] = 16'b0000000000000000;
	sram_mem[102145] = 16'b0000000000000000;
	sram_mem[102146] = 16'b0000000000000000;
	sram_mem[102147] = 16'b0000000000000000;
	sram_mem[102148] = 16'b0000000000000000;
	sram_mem[102149] = 16'b0000000000000000;
	sram_mem[102150] = 16'b0000000000000000;
	sram_mem[102151] = 16'b0000000000000000;
	sram_mem[102152] = 16'b0000000000000000;
	sram_mem[102153] = 16'b0000000000000000;
	sram_mem[102154] = 16'b0000000000000000;
	sram_mem[102155] = 16'b0000000000000000;
	sram_mem[102156] = 16'b0000000000000000;
	sram_mem[102157] = 16'b0000000000000000;
	sram_mem[102158] = 16'b0000000000000000;
	sram_mem[102159] = 16'b0000000000000000;
	sram_mem[102160] = 16'b0000000000000000;
	sram_mem[102161] = 16'b0000000000000000;
	sram_mem[102162] = 16'b0000000000000000;
	sram_mem[102163] = 16'b0000000000000000;
	sram_mem[102164] = 16'b0000000000000000;
	sram_mem[102165] = 16'b0000000000000000;
	sram_mem[102166] = 16'b0000000000000000;
	sram_mem[102167] = 16'b0000000000000000;
	sram_mem[102168] = 16'b0000000000000000;
	sram_mem[102169] = 16'b0000000000000000;
	sram_mem[102170] = 16'b0000000000000000;
	sram_mem[102171] = 16'b0000000000000000;
	sram_mem[102172] = 16'b0000000000000000;
	sram_mem[102173] = 16'b0000000000000000;
	sram_mem[102174] = 16'b0000000000000000;
	sram_mem[102175] = 16'b0000000000000000;
	sram_mem[102176] = 16'b0000000000000000;
	sram_mem[102177] = 16'b0000000000000000;
	sram_mem[102178] = 16'b0000000000000000;
	sram_mem[102179] = 16'b0000000000000000;
	sram_mem[102180] = 16'b0000000000000000;
	sram_mem[102181] = 16'b0000000000000000;
	sram_mem[102182] = 16'b0000000000000000;
	sram_mem[102183] = 16'b0000000000000000;
	sram_mem[102184] = 16'b0000000000000000;
	sram_mem[102185] = 16'b0000000000000000;
	sram_mem[102186] = 16'b0000000000000000;
	sram_mem[102187] = 16'b0000000000000000;
	sram_mem[102188] = 16'b0000000000000000;
	sram_mem[102189] = 16'b0000000000000000;
	sram_mem[102190] = 16'b0000000000000000;
	sram_mem[102191] = 16'b0000000000000000;
	sram_mem[102192] = 16'b0000000000000000;
	sram_mem[102193] = 16'b0000000000000000;
	sram_mem[102194] = 16'b0000000000000000;
	sram_mem[102195] = 16'b0000000000000000;
	sram_mem[102196] = 16'b0000000000000000;
	sram_mem[102197] = 16'b0000000000000000;
	sram_mem[102198] = 16'b0000000000000000;
	sram_mem[102199] = 16'b0000000000000000;
	sram_mem[102200] = 16'b0000000000000000;
	sram_mem[102201] = 16'b0000000000000000;
	sram_mem[102202] = 16'b0000000000000000;
	sram_mem[102203] = 16'b0000000000000000;
	sram_mem[102204] = 16'b0000000000000000;
	sram_mem[102205] = 16'b0000000000000000;
	sram_mem[102206] = 16'b0000000000000000;
	sram_mem[102207] = 16'b0000000000000000;
	sram_mem[102208] = 16'b0000000000000000;
	sram_mem[102209] = 16'b0000000000000000;
	sram_mem[102210] = 16'b0000000000000000;
	sram_mem[102211] = 16'b0000000000000000;
	sram_mem[102212] = 16'b0000000000000000;
	sram_mem[102213] = 16'b0000000000000000;
	sram_mem[102214] = 16'b0000000000000000;
	sram_mem[102215] = 16'b0000000000000000;
	sram_mem[102216] = 16'b0000000000000000;
	sram_mem[102217] = 16'b0000000000000000;
	sram_mem[102218] = 16'b0000000000000000;
	sram_mem[102219] = 16'b0000000000000000;
	sram_mem[102220] = 16'b0000000000000000;
	sram_mem[102221] = 16'b0000000000000000;
	sram_mem[102222] = 16'b0000000000000000;
	sram_mem[102223] = 16'b0000000000000000;
	sram_mem[102224] = 16'b0000000000000000;
	sram_mem[102225] = 16'b0000000000000000;
	sram_mem[102226] = 16'b0000000000000000;
	sram_mem[102227] = 16'b0000000000000000;
	sram_mem[102228] = 16'b0000000000000000;
	sram_mem[102229] = 16'b0000000000000000;
	sram_mem[102230] = 16'b0000000000000000;
	sram_mem[102231] = 16'b0000000000000000;
	sram_mem[102232] = 16'b0000000000000000;
	sram_mem[102233] = 16'b0000000000000000;
	sram_mem[102234] = 16'b0000000000000000;
	sram_mem[102235] = 16'b0000000000000000;
	sram_mem[102236] = 16'b0000000000000000;
	sram_mem[102237] = 16'b0000000000000000;
	sram_mem[102238] = 16'b0000000000000000;
	sram_mem[102239] = 16'b0000000000000000;
	sram_mem[102240] = 16'b0000000000000000;
	sram_mem[102241] = 16'b0000000000000000;
	sram_mem[102242] = 16'b0000000000000000;
	sram_mem[102243] = 16'b0000000000000000;
	sram_mem[102244] = 16'b0000000000000000;
	sram_mem[102245] = 16'b0000000000000000;
	sram_mem[102246] = 16'b0000000000000000;
	sram_mem[102247] = 16'b0000000000000000;
	sram_mem[102248] = 16'b0000000000000000;
	sram_mem[102249] = 16'b0000000000000000;
	sram_mem[102250] = 16'b0000000000000000;
	sram_mem[102251] = 16'b0000000000000000;
	sram_mem[102252] = 16'b0000000000000000;
	sram_mem[102253] = 16'b0000000000000000;
	sram_mem[102254] = 16'b0000000000000000;
	sram_mem[102255] = 16'b0000000000000000;
	sram_mem[102256] = 16'b0000000000000000;
	sram_mem[102257] = 16'b0000000000000000;
	sram_mem[102258] = 16'b0000000000000000;
	sram_mem[102259] = 16'b0000000000000000;
	sram_mem[102260] = 16'b0000000000000000;
	sram_mem[102261] = 16'b0000000000000000;
	sram_mem[102262] = 16'b0000000000000000;
	sram_mem[102263] = 16'b0000000000000000;
	sram_mem[102264] = 16'b0000000000000000;
	sram_mem[102265] = 16'b0000000000000000;
	sram_mem[102266] = 16'b0000000000000000;
	sram_mem[102267] = 16'b0000000000000000;
	sram_mem[102268] = 16'b0000000000000000;
	sram_mem[102269] = 16'b0000000000000000;
	sram_mem[102270] = 16'b0000000000000000;
	sram_mem[102271] = 16'b0000000000000000;
	sram_mem[102272] = 16'b0000000000000000;
	sram_mem[102273] = 16'b0000000000000000;
	sram_mem[102274] = 16'b0000000000000000;
	sram_mem[102275] = 16'b0000000000000000;
	sram_mem[102276] = 16'b0000000000000000;
	sram_mem[102277] = 16'b0000000000000000;
	sram_mem[102278] = 16'b0000000000000000;
	sram_mem[102279] = 16'b0000000000000000;
	sram_mem[102280] = 16'b0000000000000000;
	sram_mem[102281] = 16'b0000000000000000;
	sram_mem[102282] = 16'b0000000000000000;
	sram_mem[102283] = 16'b0000000000000000;
	sram_mem[102284] = 16'b0000000000000000;
	sram_mem[102285] = 16'b0000000000000000;
	sram_mem[102286] = 16'b0000000000000000;
	sram_mem[102287] = 16'b0000000000000000;
	sram_mem[102288] = 16'b0000000000000000;
	sram_mem[102289] = 16'b0000000000000000;
	sram_mem[102290] = 16'b0000000000000000;
	sram_mem[102291] = 16'b0000000000000000;
	sram_mem[102292] = 16'b0000000000000000;
	sram_mem[102293] = 16'b0000000000000000;
	sram_mem[102294] = 16'b0000000000000000;
	sram_mem[102295] = 16'b0000000000000000;
	sram_mem[102296] = 16'b0000000000000000;
	sram_mem[102297] = 16'b0000000000000000;
	sram_mem[102298] = 16'b0000000000000000;
	sram_mem[102299] = 16'b0000000000000000;
	sram_mem[102300] = 16'b0000000000000000;
	sram_mem[102301] = 16'b0000000000000000;
	sram_mem[102302] = 16'b0000000000000000;
	sram_mem[102303] = 16'b0000000000000000;
	sram_mem[102304] = 16'b0000000000000000;
	sram_mem[102305] = 16'b0000000000000000;
	sram_mem[102306] = 16'b0000000000000000;
	sram_mem[102307] = 16'b0000000000000000;
	sram_mem[102308] = 16'b0000000000000000;
	sram_mem[102309] = 16'b0000000000000000;
	sram_mem[102310] = 16'b0000000000000000;
	sram_mem[102311] = 16'b0000000000000000;
	sram_mem[102312] = 16'b0000000000000000;
	sram_mem[102313] = 16'b0000000000000000;
	sram_mem[102314] = 16'b0000000000000000;
	sram_mem[102315] = 16'b0000000000000000;
	sram_mem[102316] = 16'b0000000000000000;
	sram_mem[102317] = 16'b0000000000000000;
	sram_mem[102318] = 16'b0000000000000000;
	sram_mem[102319] = 16'b0000000000000000;
	sram_mem[102320] = 16'b0000000000000000;
	sram_mem[102321] = 16'b0000000000000000;
	sram_mem[102322] = 16'b0000000000000000;
	sram_mem[102323] = 16'b0000000000000000;
	sram_mem[102324] = 16'b0000000000000000;
	sram_mem[102325] = 16'b0000000000000000;
	sram_mem[102326] = 16'b0000000000000000;
	sram_mem[102327] = 16'b0000000000000000;
	sram_mem[102328] = 16'b0000000000000000;
	sram_mem[102329] = 16'b0000000000000000;
	sram_mem[102330] = 16'b0000000000000000;
	sram_mem[102331] = 16'b0000000000000000;
	sram_mem[102332] = 16'b0000000000000000;
	sram_mem[102333] = 16'b0000000000000000;
	sram_mem[102334] = 16'b0000000000000000;
	sram_mem[102335] = 16'b0000000000000000;
	sram_mem[102336] = 16'b0000000000000000;
	sram_mem[102337] = 16'b0000000000000000;
	sram_mem[102338] = 16'b0000000000000000;
	sram_mem[102339] = 16'b0000000000000000;
	sram_mem[102340] = 16'b0000000000000000;
	sram_mem[102341] = 16'b0000000000000000;
	sram_mem[102342] = 16'b0000000000000000;
	sram_mem[102343] = 16'b0000000000000000;
	sram_mem[102344] = 16'b0000000000000000;
	sram_mem[102345] = 16'b0000000000000000;
	sram_mem[102346] = 16'b0000000000000000;
	sram_mem[102347] = 16'b0000000000000000;
	sram_mem[102348] = 16'b0000000000000000;
	sram_mem[102349] = 16'b0000000000000000;
	sram_mem[102350] = 16'b0000000000000000;
	sram_mem[102351] = 16'b0000000000000000;
	sram_mem[102352] = 16'b0000000000000000;
	sram_mem[102353] = 16'b0000000000000000;
	sram_mem[102354] = 16'b0000000000000000;
	sram_mem[102355] = 16'b0000000000000000;
	sram_mem[102356] = 16'b0000000000000000;
	sram_mem[102357] = 16'b0000000000000000;
	sram_mem[102358] = 16'b0000000000000000;
	sram_mem[102359] = 16'b0000000000000000;
	sram_mem[102360] = 16'b0000000000000000;
	sram_mem[102361] = 16'b0000000000000000;
	sram_mem[102362] = 16'b0000000000000000;
	sram_mem[102363] = 16'b0000000000000000;
	sram_mem[102364] = 16'b0000000000000000;
	sram_mem[102365] = 16'b0000000000000000;
	sram_mem[102366] = 16'b0000000000000000;
	sram_mem[102367] = 16'b0000000000000000;
	sram_mem[102368] = 16'b0000000000000000;
	sram_mem[102369] = 16'b0000000000000000;
	sram_mem[102370] = 16'b0000000000000000;
	sram_mem[102371] = 16'b0000000000000000;
	sram_mem[102372] = 16'b0000000000000000;
	sram_mem[102373] = 16'b0000000000000000;
	sram_mem[102374] = 16'b0000000000000000;
	sram_mem[102375] = 16'b0000000000000000;
	sram_mem[102376] = 16'b0000000000000000;
	sram_mem[102377] = 16'b0000000000000000;
	sram_mem[102378] = 16'b0000000000000000;
	sram_mem[102379] = 16'b0000000000000000;
	sram_mem[102380] = 16'b0000000000000000;
	sram_mem[102381] = 16'b0000000000000000;
	sram_mem[102382] = 16'b0000000000000000;
	sram_mem[102383] = 16'b0000000000000000;
	sram_mem[102384] = 16'b0000000000000000;
	sram_mem[102385] = 16'b0000000000000000;
	sram_mem[102386] = 16'b0000000000000000;
	sram_mem[102387] = 16'b0000000000000000;
	sram_mem[102388] = 16'b0000000000000000;
	sram_mem[102389] = 16'b0000000000000000;
	sram_mem[102390] = 16'b0000000000000000;
	sram_mem[102391] = 16'b0000000000000000;
	sram_mem[102392] = 16'b0000000000000000;
	sram_mem[102393] = 16'b0000000000000000;
	sram_mem[102394] = 16'b0000000000000000;
	sram_mem[102395] = 16'b0000000000000000;
	sram_mem[102396] = 16'b0000000000000000;
	sram_mem[102397] = 16'b0000000000000000;
	sram_mem[102398] = 16'b0000000000000000;
	sram_mem[102399] = 16'b0000000000000000;
	sram_mem[102400] = 16'b0000000000000000;
	sram_mem[102401] = 16'b0000000000000000;
	sram_mem[102402] = 16'b0000000000000000;
	sram_mem[102403] = 16'b0000000000000000;
	sram_mem[102404] = 16'b0000000000000000;
	sram_mem[102405] = 16'b0000000000000000;
	sram_mem[102406] = 16'b0000000000000000;
	sram_mem[102407] = 16'b0000000000000000;
	sram_mem[102408] = 16'b0000000000000000;
	sram_mem[102409] = 16'b0000000000000000;
	sram_mem[102410] = 16'b0000000000000000;
	sram_mem[102411] = 16'b0000000000000000;
	sram_mem[102412] = 16'b0000000000000000;
	sram_mem[102413] = 16'b0000000000000000;
	sram_mem[102414] = 16'b0000000000000000;
	sram_mem[102415] = 16'b0000000000000000;
	sram_mem[102416] = 16'b0000000000000000;
	sram_mem[102417] = 16'b0000000000000000;
	sram_mem[102418] = 16'b0000000000000000;
	sram_mem[102419] = 16'b0000000000000000;
	sram_mem[102420] = 16'b0000000000000000;
	sram_mem[102421] = 16'b0000000000000000;
	sram_mem[102422] = 16'b0000000000000000;
	sram_mem[102423] = 16'b0000000000000000;
	sram_mem[102424] = 16'b0000000000000000;
	sram_mem[102425] = 16'b0000000000000000;
	sram_mem[102426] = 16'b0000000000000000;
	sram_mem[102427] = 16'b0000000000000000;
	sram_mem[102428] = 16'b0000000000000000;
	sram_mem[102429] = 16'b0000000000000000;
	sram_mem[102430] = 16'b0000000000000000;
	sram_mem[102431] = 16'b0000000000000000;
	sram_mem[102432] = 16'b0000000000000000;
	sram_mem[102433] = 16'b0000000000000000;
	sram_mem[102434] = 16'b0000000000000000;
	sram_mem[102435] = 16'b0000000000000000;
	sram_mem[102436] = 16'b0000000000000000;
	sram_mem[102437] = 16'b0000000000000000;
	sram_mem[102438] = 16'b0000000000000000;
	sram_mem[102439] = 16'b0000000000000000;
	sram_mem[102440] = 16'b0000000000000000;
	sram_mem[102441] = 16'b0000000000000000;
	sram_mem[102442] = 16'b0000000000000000;
	sram_mem[102443] = 16'b0000000000000000;
	sram_mem[102444] = 16'b0000000000000000;
	sram_mem[102445] = 16'b0000000000000000;
	sram_mem[102446] = 16'b0000000000000000;
	sram_mem[102447] = 16'b0000000000000000;
	sram_mem[102448] = 16'b0000000000000000;
	sram_mem[102449] = 16'b0000000000000000;
	sram_mem[102450] = 16'b0000000000000000;
	sram_mem[102451] = 16'b0000000000000000;
	sram_mem[102452] = 16'b0000000000000000;
	sram_mem[102453] = 16'b0000000000000000;
	sram_mem[102454] = 16'b0000000000000000;
	sram_mem[102455] = 16'b0000000000000000;
	sram_mem[102456] = 16'b0000000000000000;
	sram_mem[102457] = 16'b0000000000000000;
	sram_mem[102458] = 16'b0000000000000000;
	sram_mem[102459] = 16'b0000000000000000;
	sram_mem[102460] = 16'b0000000000000000;
	sram_mem[102461] = 16'b0000000000000000;
	sram_mem[102462] = 16'b0000000000000000;
	sram_mem[102463] = 16'b0000000000000000;
	sram_mem[102464] = 16'b0000000000000000;
	sram_mem[102465] = 16'b0000000000000000;
	sram_mem[102466] = 16'b0000000000000000;
	sram_mem[102467] = 16'b0000000000000000;
	sram_mem[102468] = 16'b0000000000000000;
	sram_mem[102469] = 16'b0000000000000000;
	sram_mem[102470] = 16'b0000000000000000;
	sram_mem[102471] = 16'b0000000000000000;
	sram_mem[102472] = 16'b0000000000000000;
	sram_mem[102473] = 16'b0000000000000000;
	sram_mem[102474] = 16'b0000000000000000;
	sram_mem[102475] = 16'b0000000000000000;
	sram_mem[102476] = 16'b0000000000000000;
	sram_mem[102477] = 16'b0000000000000000;
	sram_mem[102478] = 16'b0000000000000000;
	sram_mem[102479] = 16'b0000000000000000;
	sram_mem[102480] = 16'b0000000000000000;
	sram_mem[102481] = 16'b0000000000000000;
	sram_mem[102482] = 16'b0000000000000000;
	sram_mem[102483] = 16'b0000000000000000;
	sram_mem[102484] = 16'b0000000000000000;
	sram_mem[102485] = 16'b0000000000000000;
	sram_mem[102486] = 16'b0000000000000000;
	sram_mem[102487] = 16'b0000000000000000;
	sram_mem[102488] = 16'b0000000000000000;
	sram_mem[102489] = 16'b0000000000000000;
	sram_mem[102490] = 16'b0000000000000000;
	sram_mem[102491] = 16'b0000000000000000;
	sram_mem[102492] = 16'b0000000000000000;
	sram_mem[102493] = 16'b0000000000000000;
	sram_mem[102494] = 16'b0000000000000000;
	sram_mem[102495] = 16'b0000000000000000;
	sram_mem[102496] = 16'b0000000000000000;
	sram_mem[102497] = 16'b0000000000000000;
	sram_mem[102498] = 16'b0000000000000000;
	sram_mem[102499] = 16'b0000000000000000;
	sram_mem[102500] = 16'b0000000000000000;
	sram_mem[102501] = 16'b0000000000000000;
	sram_mem[102502] = 16'b0000000000000000;
	sram_mem[102503] = 16'b0000000000000000;
	sram_mem[102504] = 16'b0000000000000000;
	sram_mem[102505] = 16'b0000000000000000;
	sram_mem[102506] = 16'b0000000000000000;
	sram_mem[102507] = 16'b0000000000000000;
	sram_mem[102508] = 16'b0000000000000000;
	sram_mem[102509] = 16'b0000000000000000;
	sram_mem[102510] = 16'b0000000000000000;
	sram_mem[102511] = 16'b0000000000000000;
	sram_mem[102512] = 16'b0000000000000000;
	sram_mem[102513] = 16'b0000000000000000;
	sram_mem[102514] = 16'b0000000000000000;
	sram_mem[102515] = 16'b0000000000000000;
	sram_mem[102516] = 16'b0000000000000000;
	sram_mem[102517] = 16'b0000000000000000;
	sram_mem[102518] = 16'b0000000000000000;
	sram_mem[102519] = 16'b0000000000000000;
	sram_mem[102520] = 16'b0000000000000000;
	sram_mem[102521] = 16'b0000000000000000;
	sram_mem[102522] = 16'b0000000000000000;
	sram_mem[102523] = 16'b0000000000000000;
	sram_mem[102524] = 16'b0000000000000000;
	sram_mem[102525] = 16'b0000000000000000;
	sram_mem[102526] = 16'b0000000000000000;
	sram_mem[102527] = 16'b0000000000000000;
	sram_mem[102528] = 16'b0000000000000000;
	sram_mem[102529] = 16'b0000000000000000;
	sram_mem[102530] = 16'b0000000000000000;
	sram_mem[102531] = 16'b0000000000000000;
	sram_mem[102532] = 16'b0000000000000000;
	sram_mem[102533] = 16'b0000000000000000;
	sram_mem[102534] = 16'b0000000000000000;
	sram_mem[102535] = 16'b0000000000000000;
	sram_mem[102536] = 16'b0000000000000000;
	sram_mem[102537] = 16'b0000000000000000;
	sram_mem[102538] = 16'b0000000000000000;
	sram_mem[102539] = 16'b0000000000000000;
	sram_mem[102540] = 16'b0000000000000000;
	sram_mem[102541] = 16'b0000000000000000;
	sram_mem[102542] = 16'b0000000000000000;
	sram_mem[102543] = 16'b0000000000000000;
	sram_mem[102544] = 16'b0000000000000000;
	sram_mem[102545] = 16'b0000000000000000;
	sram_mem[102546] = 16'b0000000000000000;
	sram_mem[102547] = 16'b0000000000000000;
	sram_mem[102548] = 16'b0000000000000000;
	sram_mem[102549] = 16'b0000000000000000;
	sram_mem[102550] = 16'b0000000000000000;
	sram_mem[102551] = 16'b0000000000000000;
	sram_mem[102552] = 16'b0000000000000000;
	sram_mem[102553] = 16'b0000000000000000;
	sram_mem[102554] = 16'b0000000000000000;
	sram_mem[102555] = 16'b0000000000000000;
	sram_mem[102556] = 16'b0000000000000000;
	sram_mem[102557] = 16'b0000000000000000;
	sram_mem[102558] = 16'b0000000000000000;
	sram_mem[102559] = 16'b0000000000000000;
	sram_mem[102560] = 16'b0000000000000000;
	sram_mem[102561] = 16'b0000000000000000;
	sram_mem[102562] = 16'b0000000000000000;
	sram_mem[102563] = 16'b0000000000000000;
	sram_mem[102564] = 16'b0000000000000000;
	sram_mem[102565] = 16'b0000000000000000;
	sram_mem[102566] = 16'b0000000000000000;
	sram_mem[102567] = 16'b0000000000000000;
	sram_mem[102568] = 16'b0000000000000000;
	sram_mem[102569] = 16'b0000000000000000;
	sram_mem[102570] = 16'b0000000000000000;
	sram_mem[102571] = 16'b0000000000000000;
	sram_mem[102572] = 16'b0000000000000000;
	sram_mem[102573] = 16'b0000000000000000;
	sram_mem[102574] = 16'b0000000000000000;
	sram_mem[102575] = 16'b0000000000000000;
	sram_mem[102576] = 16'b0000000000000000;
	sram_mem[102577] = 16'b0000000000000000;
	sram_mem[102578] = 16'b0000000000000000;
	sram_mem[102579] = 16'b0000000000000000;
	sram_mem[102580] = 16'b0000000000000000;
	sram_mem[102581] = 16'b0000000000000000;
	sram_mem[102582] = 16'b0000000000000000;
	sram_mem[102583] = 16'b0000000000000000;
	sram_mem[102584] = 16'b0000000000000000;
	sram_mem[102585] = 16'b0000000000000000;
	sram_mem[102586] = 16'b0000000000000000;
	sram_mem[102587] = 16'b0000000000000000;
	sram_mem[102588] = 16'b0000000000000000;
	sram_mem[102589] = 16'b0000000000000000;
	sram_mem[102590] = 16'b0000000000000000;
	sram_mem[102591] = 16'b0000000000000000;
	sram_mem[102592] = 16'b0000000000000000;
	sram_mem[102593] = 16'b0000000000000000;
	sram_mem[102594] = 16'b0000000000000000;
	sram_mem[102595] = 16'b0000000000000000;
	sram_mem[102596] = 16'b0000000000000000;
	sram_mem[102597] = 16'b0000000000000000;
	sram_mem[102598] = 16'b0000000000000000;
	sram_mem[102599] = 16'b0000000000000000;
	sram_mem[102600] = 16'b0000000000000000;
	sram_mem[102601] = 16'b0000000000000000;
	sram_mem[102602] = 16'b0000000000000000;
	sram_mem[102603] = 16'b0000000000000000;
	sram_mem[102604] = 16'b0000000000000000;
	sram_mem[102605] = 16'b0000000000000000;
	sram_mem[102606] = 16'b0000000000000000;
	sram_mem[102607] = 16'b0000000000000000;
	sram_mem[102608] = 16'b0000000000000000;
	sram_mem[102609] = 16'b0000000000000000;
	sram_mem[102610] = 16'b0000000000000000;
	sram_mem[102611] = 16'b0000000000000000;
	sram_mem[102612] = 16'b0000000000000000;
	sram_mem[102613] = 16'b0000000000000000;
	sram_mem[102614] = 16'b0000000000000000;
	sram_mem[102615] = 16'b0000000000000000;
	sram_mem[102616] = 16'b0000000000000000;
	sram_mem[102617] = 16'b0000000000000000;
	sram_mem[102618] = 16'b0000000000000000;
	sram_mem[102619] = 16'b0000000000000000;
	sram_mem[102620] = 16'b0000000000000000;
	sram_mem[102621] = 16'b0000000000000000;
	sram_mem[102622] = 16'b0000000000000000;
	sram_mem[102623] = 16'b0000000000000000;
	sram_mem[102624] = 16'b0000000000000000;
	sram_mem[102625] = 16'b0000000000000000;
	sram_mem[102626] = 16'b0000000000000000;
	sram_mem[102627] = 16'b0000000000000000;
	sram_mem[102628] = 16'b0000000000000000;
	sram_mem[102629] = 16'b0000000000000000;
	sram_mem[102630] = 16'b0000000000000000;
	sram_mem[102631] = 16'b0000000000000000;
	sram_mem[102632] = 16'b0000000000000000;
	sram_mem[102633] = 16'b0000000000000000;
	sram_mem[102634] = 16'b0000000000000000;
	sram_mem[102635] = 16'b0000000000000000;
	sram_mem[102636] = 16'b0000000000000000;
	sram_mem[102637] = 16'b0000000000000000;
	sram_mem[102638] = 16'b0000000000000000;
	sram_mem[102639] = 16'b0000000000000000;
	sram_mem[102640] = 16'b0000000000000000;
	sram_mem[102641] = 16'b0000000000000000;
	sram_mem[102642] = 16'b0000000000000000;
	sram_mem[102643] = 16'b0000000000000000;
	sram_mem[102644] = 16'b0000000000000000;
	sram_mem[102645] = 16'b0000000000000000;
	sram_mem[102646] = 16'b0000000000000000;
	sram_mem[102647] = 16'b0000000000000000;
	sram_mem[102648] = 16'b0000000000000000;
	sram_mem[102649] = 16'b0000000000000000;
	sram_mem[102650] = 16'b0000000000000000;
	sram_mem[102651] = 16'b0000000000000000;
	sram_mem[102652] = 16'b0000000000000000;
	sram_mem[102653] = 16'b0000000000000000;
	sram_mem[102654] = 16'b0000000000000000;
	sram_mem[102655] = 16'b0000000000000000;
	sram_mem[102656] = 16'b0000000000000000;
	sram_mem[102657] = 16'b0000000000000000;
	sram_mem[102658] = 16'b0000000000000000;
	sram_mem[102659] = 16'b0000000000000000;
	sram_mem[102660] = 16'b0000000000000000;
	sram_mem[102661] = 16'b0000000000000000;
	sram_mem[102662] = 16'b0000000000000000;
	sram_mem[102663] = 16'b0000000000000000;
	sram_mem[102664] = 16'b0000000000000000;
	sram_mem[102665] = 16'b0000000000000000;
	sram_mem[102666] = 16'b0000000000000000;
	sram_mem[102667] = 16'b0000000000000000;
	sram_mem[102668] = 16'b0000000000000000;
	sram_mem[102669] = 16'b0000000000000000;
	sram_mem[102670] = 16'b0000000000000000;
	sram_mem[102671] = 16'b0000000000000000;
	sram_mem[102672] = 16'b0000000000000000;
	sram_mem[102673] = 16'b0000000000000000;
	sram_mem[102674] = 16'b0000000000000000;
	sram_mem[102675] = 16'b0000000000000000;
	sram_mem[102676] = 16'b0000000000000000;
	sram_mem[102677] = 16'b0000000000000000;
	sram_mem[102678] = 16'b0000000000000000;
	sram_mem[102679] = 16'b0000000000000000;
	sram_mem[102680] = 16'b0000000000000000;
	sram_mem[102681] = 16'b0000000000000000;
	sram_mem[102682] = 16'b0000000000000000;
	sram_mem[102683] = 16'b0000000000000000;
	sram_mem[102684] = 16'b0000000000000000;
	sram_mem[102685] = 16'b0000000000000000;
	sram_mem[102686] = 16'b0000000000000000;
	sram_mem[102687] = 16'b0000000000000000;
	sram_mem[102688] = 16'b0000000000000000;
	sram_mem[102689] = 16'b0000000000000000;
	sram_mem[102690] = 16'b0000000000000000;
	sram_mem[102691] = 16'b0000000000000000;
	sram_mem[102692] = 16'b0000000000000000;
	sram_mem[102693] = 16'b0000000000000000;
	sram_mem[102694] = 16'b0000000000000000;
	sram_mem[102695] = 16'b0000000000000000;
	sram_mem[102696] = 16'b0000000000000000;
	sram_mem[102697] = 16'b0000000000000000;
	sram_mem[102698] = 16'b0000000000000000;
	sram_mem[102699] = 16'b0000000000000000;
	sram_mem[102700] = 16'b0000000000000000;
	sram_mem[102701] = 16'b0000000000000000;
	sram_mem[102702] = 16'b0000000000000000;
	sram_mem[102703] = 16'b0000000000000000;
	sram_mem[102704] = 16'b0000000000000000;
	sram_mem[102705] = 16'b0000000000000000;
	sram_mem[102706] = 16'b0000000000000000;
	sram_mem[102707] = 16'b0000000000000000;
	sram_mem[102708] = 16'b0000000000000000;
	sram_mem[102709] = 16'b0000000000000000;
	sram_mem[102710] = 16'b0000000000000000;
	sram_mem[102711] = 16'b0000000000000000;
	sram_mem[102712] = 16'b0000000000000000;
	sram_mem[102713] = 16'b0000000000000000;
	sram_mem[102714] = 16'b0000000000000000;
	sram_mem[102715] = 16'b0000000000000000;
	sram_mem[102716] = 16'b0000000000000000;
	sram_mem[102717] = 16'b0000000000000000;
	sram_mem[102718] = 16'b0000000000000000;
	sram_mem[102719] = 16'b0000000000000000;
	sram_mem[102720] = 16'b0000000000000000;
	sram_mem[102721] = 16'b0000000000000000;
	sram_mem[102722] = 16'b0000000000000000;
	sram_mem[102723] = 16'b0000000000000000;
	sram_mem[102724] = 16'b0000000000000000;
	sram_mem[102725] = 16'b0000000000000000;
	sram_mem[102726] = 16'b0000000000000000;
	sram_mem[102727] = 16'b0000000000000000;
	sram_mem[102728] = 16'b0000000000000000;
	sram_mem[102729] = 16'b0000000000000000;
	sram_mem[102730] = 16'b0000000000000000;
	sram_mem[102731] = 16'b0000000000000000;
	sram_mem[102732] = 16'b0000000000000000;
	sram_mem[102733] = 16'b0000000000000000;
	sram_mem[102734] = 16'b0000000000000000;
	sram_mem[102735] = 16'b0000000000000000;
	sram_mem[102736] = 16'b0000000000000000;
	sram_mem[102737] = 16'b0000000000000000;
	sram_mem[102738] = 16'b0000000000000000;
	sram_mem[102739] = 16'b0000000000000000;
	sram_mem[102740] = 16'b0000000000000000;
	sram_mem[102741] = 16'b0000000000000000;
	sram_mem[102742] = 16'b0000000000000000;
	sram_mem[102743] = 16'b0000000000000000;
	sram_mem[102744] = 16'b0000000000000000;
	sram_mem[102745] = 16'b0000000000000000;
	sram_mem[102746] = 16'b0000000000000000;
	sram_mem[102747] = 16'b0000000000000000;
	sram_mem[102748] = 16'b0000000000000000;
	sram_mem[102749] = 16'b0000000000000000;
	sram_mem[102750] = 16'b0000000000000000;
	sram_mem[102751] = 16'b0000000000000000;
	sram_mem[102752] = 16'b0000000000000000;
	sram_mem[102753] = 16'b0000000000000000;
	sram_mem[102754] = 16'b0000000000000000;
	sram_mem[102755] = 16'b0000000000000000;
	sram_mem[102756] = 16'b0000000000000000;
	sram_mem[102757] = 16'b0000000000000000;
	sram_mem[102758] = 16'b0000000000000000;
	sram_mem[102759] = 16'b0000000000000000;
	sram_mem[102760] = 16'b0000000000000000;
	sram_mem[102761] = 16'b0000000000000000;
	sram_mem[102762] = 16'b0000000000000000;
	sram_mem[102763] = 16'b0000000000000000;
	sram_mem[102764] = 16'b0000000000000000;
	sram_mem[102765] = 16'b0000000000000000;
	sram_mem[102766] = 16'b0000000000000000;
	sram_mem[102767] = 16'b0000000000000000;
	sram_mem[102768] = 16'b0000000000000000;
	sram_mem[102769] = 16'b0000000000000000;
	sram_mem[102770] = 16'b0000000000000000;
	sram_mem[102771] = 16'b0000000000000000;
	sram_mem[102772] = 16'b0000000000000000;
	sram_mem[102773] = 16'b0000000000000000;
	sram_mem[102774] = 16'b0000000000000000;
	sram_mem[102775] = 16'b0000000000000000;
	sram_mem[102776] = 16'b0000000000000000;
	sram_mem[102777] = 16'b0000000000000000;
	sram_mem[102778] = 16'b0000000000000000;
	sram_mem[102779] = 16'b0000000000000000;
	sram_mem[102780] = 16'b0000000000000000;
	sram_mem[102781] = 16'b0000000000000000;
	sram_mem[102782] = 16'b0000000000000000;
	sram_mem[102783] = 16'b0000000000000000;
	sram_mem[102784] = 16'b0000000000000000;
	sram_mem[102785] = 16'b0000000000000000;
	sram_mem[102786] = 16'b0000000000000000;
	sram_mem[102787] = 16'b0000000000000000;
	sram_mem[102788] = 16'b0000000000000000;
	sram_mem[102789] = 16'b0000000000000000;
	sram_mem[102790] = 16'b0000000000000000;
	sram_mem[102791] = 16'b0000000000000000;
	sram_mem[102792] = 16'b0000000000000000;
	sram_mem[102793] = 16'b0000000000000000;
	sram_mem[102794] = 16'b0000000000000000;
	sram_mem[102795] = 16'b0000000000000000;
	sram_mem[102796] = 16'b0000000000000000;
	sram_mem[102797] = 16'b0000000000000000;
	sram_mem[102798] = 16'b0000000000000000;
	sram_mem[102799] = 16'b0000000000000000;
	sram_mem[102800] = 16'b0000000000000000;
	sram_mem[102801] = 16'b0000000000000000;
	sram_mem[102802] = 16'b0000000000000000;
	sram_mem[102803] = 16'b0000000000000000;
	sram_mem[102804] = 16'b0000000000000000;
	sram_mem[102805] = 16'b0000000000000000;
	sram_mem[102806] = 16'b0000000000000000;
	sram_mem[102807] = 16'b0000000000000000;
	sram_mem[102808] = 16'b0000000000000000;
	sram_mem[102809] = 16'b0000000000000000;
	sram_mem[102810] = 16'b0000000000000000;
	sram_mem[102811] = 16'b0000000000000000;
	sram_mem[102812] = 16'b0000000000000000;
	sram_mem[102813] = 16'b0000000000000000;
	sram_mem[102814] = 16'b0000000000000000;
	sram_mem[102815] = 16'b0000000000000000;
	sram_mem[102816] = 16'b0000000000000000;
	sram_mem[102817] = 16'b0000000000000000;
	sram_mem[102818] = 16'b0000000000000000;
	sram_mem[102819] = 16'b0000000000000000;
	sram_mem[102820] = 16'b0000000000000000;
	sram_mem[102821] = 16'b0000000000000000;
	sram_mem[102822] = 16'b0000000000000000;
	sram_mem[102823] = 16'b0000000000000000;
	sram_mem[102824] = 16'b0000000000000000;
	sram_mem[102825] = 16'b0000000000000000;
	sram_mem[102826] = 16'b0000000000000000;
	sram_mem[102827] = 16'b0000000000000000;
	sram_mem[102828] = 16'b0000000000000000;
	sram_mem[102829] = 16'b0000000000000000;
	sram_mem[102830] = 16'b0000000000000000;
	sram_mem[102831] = 16'b0000000000000000;
	sram_mem[102832] = 16'b0000000000000000;
	sram_mem[102833] = 16'b0000000000000000;
	sram_mem[102834] = 16'b0000000000000000;
	sram_mem[102835] = 16'b0000000000000000;
	sram_mem[102836] = 16'b0000000000000000;
	sram_mem[102837] = 16'b0000000000000000;
	sram_mem[102838] = 16'b0000000000000000;
	sram_mem[102839] = 16'b0000000000000000;
	sram_mem[102840] = 16'b0000000000000000;
	sram_mem[102841] = 16'b0000000000000000;
	sram_mem[102842] = 16'b0000000000000000;
	sram_mem[102843] = 16'b0000000000000000;
	sram_mem[102844] = 16'b0000000000000000;
	sram_mem[102845] = 16'b0000000000000000;
	sram_mem[102846] = 16'b0000000000000000;
	sram_mem[102847] = 16'b0000000000000000;
	sram_mem[102848] = 16'b0000000000000000;
	sram_mem[102849] = 16'b0000000000000000;
	sram_mem[102850] = 16'b0000000000000000;
	sram_mem[102851] = 16'b0000000000000000;
	sram_mem[102852] = 16'b0000000000000000;
	sram_mem[102853] = 16'b0000000000000000;
	sram_mem[102854] = 16'b0000000000000000;
	sram_mem[102855] = 16'b0000000000000000;
	sram_mem[102856] = 16'b0000000000000000;
	sram_mem[102857] = 16'b0000000000000000;
	sram_mem[102858] = 16'b0000000000000000;
	sram_mem[102859] = 16'b0000000000000000;
	sram_mem[102860] = 16'b0000000000000000;
	sram_mem[102861] = 16'b0000000000000000;
	sram_mem[102862] = 16'b0000000000000000;
	sram_mem[102863] = 16'b0000000000000000;
	sram_mem[102864] = 16'b0000000000000000;
	sram_mem[102865] = 16'b0000000000000000;
	sram_mem[102866] = 16'b0000000000000000;
	sram_mem[102867] = 16'b0000000000000000;
	sram_mem[102868] = 16'b0000000000000000;
	sram_mem[102869] = 16'b0000000000000000;
	sram_mem[102870] = 16'b0000000000000000;
	sram_mem[102871] = 16'b0000000000000000;
	sram_mem[102872] = 16'b0000000000000000;
	sram_mem[102873] = 16'b0000000000000000;
	sram_mem[102874] = 16'b0000000000000000;
	sram_mem[102875] = 16'b0000000000000000;
	sram_mem[102876] = 16'b0000000000000000;
	sram_mem[102877] = 16'b0000000000000000;
	sram_mem[102878] = 16'b0000000000000000;
	sram_mem[102879] = 16'b0000000000000000;
	sram_mem[102880] = 16'b0000000000000000;
	sram_mem[102881] = 16'b0000000000000000;
	sram_mem[102882] = 16'b0000000000000000;
	sram_mem[102883] = 16'b0000000000000000;
	sram_mem[102884] = 16'b0000000000000000;
	sram_mem[102885] = 16'b0000000000000000;
	sram_mem[102886] = 16'b0000000000000000;
	sram_mem[102887] = 16'b0000000000000000;
	sram_mem[102888] = 16'b0000000000000000;
	sram_mem[102889] = 16'b0000000000000000;
	sram_mem[102890] = 16'b0000000000000000;
	sram_mem[102891] = 16'b0000000000000000;
	sram_mem[102892] = 16'b0000000000000000;
	sram_mem[102893] = 16'b0000000000000000;
	sram_mem[102894] = 16'b0000000000000000;
	sram_mem[102895] = 16'b0000000000000000;
	sram_mem[102896] = 16'b0000000000000000;
	sram_mem[102897] = 16'b0000000000000000;
	sram_mem[102898] = 16'b0000000000000000;
	sram_mem[102899] = 16'b0000000000000000;
	sram_mem[102900] = 16'b0000000000000000;
	sram_mem[102901] = 16'b0000000000000000;
	sram_mem[102902] = 16'b0000000000000000;
	sram_mem[102903] = 16'b0000000000000000;
	sram_mem[102904] = 16'b0000000000000000;
	sram_mem[102905] = 16'b0000000000000000;
	sram_mem[102906] = 16'b0000000000000000;
	sram_mem[102907] = 16'b0000000000000000;
	sram_mem[102908] = 16'b0000000000000000;
	sram_mem[102909] = 16'b0000000000000000;
	sram_mem[102910] = 16'b0000000000000000;
	sram_mem[102911] = 16'b0000000000000000;
	sram_mem[102912] = 16'b0000000000000000;
	sram_mem[102913] = 16'b0000000000000000;
	sram_mem[102914] = 16'b0000000000000000;
	sram_mem[102915] = 16'b0000000000000000;
	sram_mem[102916] = 16'b0000000000000000;
	sram_mem[102917] = 16'b0000000000000000;
	sram_mem[102918] = 16'b0000000000000000;
	sram_mem[102919] = 16'b0000000000000000;
	sram_mem[102920] = 16'b0000000000000000;
	sram_mem[102921] = 16'b0000000000000000;
	sram_mem[102922] = 16'b0000000000000000;
	sram_mem[102923] = 16'b0000000000000000;
	sram_mem[102924] = 16'b0000000000000000;
	sram_mem[102925] = 16'b0000000000000000;
	sram_mem[102926] = 16'b0000000000000000;
	sram_mem[102927] = 16'b0000000000000000;
	sram_mem[102928] = 16'b0000000000000000;
	sram_mem[102929] = 16'b0000000000000000;
	sram_mem[102930] = 16'b0000000000000000;
	sram_mem[102931] = 16'b0000000000000000;
	sram_mem[102932] = 16'b0000000000000000;
	sram_mem[102933] = 16'b0000000000000000;
	sram_mem[102934] = 16'b0000000000000000;
	sram_mem[102935] = 16'b0000000000000000;
	sram_mem[102936] = 16'b0000000000000000;
	sram_mem[102937] = 16'b0000000000000000;
	sram_mem[102938] = 16'b0000000000000000;
	sram_mem[102939] = 16'b0000000000000000;
	sram_mem[102940] = 16'b0000000000000000;
	sram_mem[102941] = 16'b0000000000000000;
	sram_mem[102942] = 16'b0000000000000000;
	sram_mem[102943] = 16'b0000000000000000;
	sram_mem[102944] = 16'b0000000000000000;
	sram_mem[102945] = 16'b0000000000000000;
	sram_mem[102946] = 16'b0000000000000000;
	sram_mem[102947] = 16'b0000000000000000;
	sram_mem[102948] = 16'b0000000000000000;
	sram_mem[102949] = 16'b0000000000000000;
	sram_mem[102950] = 16'b0000000000000000;
	sram_mem[102951] = 16'b0000000000000000;
	sram_mem[102952] = 16'b0000000000000000;
	sram_mem[102953] = 16'b0000000000000000;
	sram_mem[102954] = 16'b0000000000000000;
	sram_mem[102955] = 16'b0000000000000000;
	sram_mem[102956] = 16'b0000000000000000;
	sram_mem[102957] = 16'b0000000000000000;
	sram_mem[102958] = 16'b0000000000000000;
	sram_mem[102959] = 16'b0000000000000000;
	sram_mem[102960] = 16'b0000000000000000;
	sram_mem[102961] = 16'b0000000000000000;
	sram_mem[102962] = 16'b0000000000000000;
	sram_mem[102963] = 16'b0000000000000000;
	sram_mem[102964] = 16'b0000000000000000;
	sram_mem[102965] = 16'b0000000000000000;
	sram_mem[102966] = 16'b0000000000000000;
	sram_mem[102967] = 16'b0000000000000000;
	sram_mem[102968] = 16'b0000000000000000;
	sram_mem[102969] = 16'b0000000000000000;
	sram_mem[102970] = 16'b0000000000000000;
	sram_mem[102971] = 16'b0000000000000000;
	sram_mem[102972] = 16'b0000000000000000;
	sram_mem[102973] = 16'b0000000000000000;
	sram_mem[102974] = 16'b0000000000000000;
	sram_mem[102975] = 16'b0000000000000000;
	sram_mem[102976] = 16'b0000000000000000;
	sram_mem[102977] = 16'b0000000000000000;
	sram_mem[102978] = 16'b0000000000000000;
	sram_mem[102979] = 16'b0000000000000000;
	sram_mem[102980] = 16'b0000000000000000;
	sram_mem[102981] = 16'b0000000000000000;
	sram_mem[102982] = 16'b0000000000000000;
	sram_mem[102983] = 16'b0000000000000000;
	sram_mem[102984] = 16'b0000000000000000;
	sram_mem[102985] = 16'b0000000000000000;
	sram_mem[102986] = 16'b0000000000000000;
	sram_mem[102987] = 16'b0000000000000000;
	sram_mem[102988] = 16'b0000000000000000;
	sram_mem[102989] = 16'b0000000000000000;
	sram_mem[102990] = 16'b0000000000000000;
	sram_mem[102991] = 16'b0000000000000000;
	sram_mem[102992] = 16'b0000000000000000;
	sram_mem[102993] = 16'b0000000000000000;
	sram_mem[102994] = 16'b0000000000000000;
	sram_mem[102995] = 16'b0000000000000000;
	sram_mem[102996] = 16'b0000000000000000;
	sram_mem[102997] = 16'b0000000000000000;
	sram_mem[102998] = 16'b0000000000000000;
	sram_mem[102999] = 16'b0000000000000000;
	sram_mem[103000] = 16'b0000000000000000;
	sram_mem[103001] = 16'b0000000000000000;
	sram_mem[103002] = 16'b0000000000000000;
	sram_mem[103003] = 16'b0000000000000000;
	sram_mem[103004] = 16'b0000000000000000;
	sram_mem[103005] = 16'b0000000000000000;
	sram_mem[103006] = 16'b0000000000000000;
	sram_mem[103007] = 16'b0000000000000000;
	sram_mem[103008] = 16'b0000000000000000;
	sram_mem[103009] = 16'b0000000000000000;
	sram_mem[103010] = 16'b0000000000000000;
	sram_mem[103011] = 16'b0000000000000000;
	sram_mem[103012] = 16'b0000000000000000;
	sram_mem[103013] = 16'b0000000000000000;
	sram_mem[103014] = 16'b0000000000000000;
	sram_mem[103015] = 16'b0000000000000000;
	sram_mem[103016] = 16'b0000000000000000;
	sram_mem[103017] = 16'b0000000000000000;
	sram_mem[103018] = 16'b0000000000000000;
	sram_mem[103019] = 16'b0000000000000000;
	sram_mem[103020] = 16'b0000000000000000;
	sram_mem[103021] = 16'b0000000000000000;
	sram_mem[103022] = 16'b0000000000000000;
	sram_mem[103023] = 16'b0000000000000000;
	sram_mem[103024] = 16'b0000000000000000;
	sram_mem[103025] = 16'b0000000000000000;
	sram_mem[103026] = 16'b0000000000000000;
	sram_mem[103027] = 16'b0000000000000000;
	sram_mem[103028] = 16'b0000000000000000;
	sram_mem[103029] = 16'b0000000000000000;
	sram_mem[103030] = 16'b0000000000000000;
	sram_mem[103031] = 16'b0000000000000000;
	sram_mem[103032] = 16'b0000000000000000;
	sram_mem[103033] = 16'b0000000000000000;
	sram_mem[103034] = 16'b0000000000000000;
	sram_mem[103035] = 16'b0000000000000000;
	sram_mem[103036] = 16'b0000000000000000;
	sram_mem[103037] = 16'b0000000000000000;
	sram_mem[103038] = 16'b0000000000000000;
	sram_mem[103039] = 16'b0000000000000000;
	sram_mem[103040] = 16'b0000000000000000;
	sram_mem[103041] = 16'b0000000000000000;
	sram_mem[103042] = 16'b0000000000000000;
	sram_mem[103043] = 16'b0000000000000000;
	sram_mem[103044] = 16'b0000000000000000;
	sram_mem[103045] = 16'b0000000000000000;
	sram_mem[103046] = 16'b0000000000000000;
	sram_mem[103047] = 16'b0000000000000000;
	sram_mem[103048] = 16'b0000000000000000;
	sram_mem[103049] = 16'b0000000000000000;
	sram_mem[103050] = 16'b0000000000000000;
	sram_mem[103051] = 16'b0000000000000000;
	sram_mem[103052] = 16'b0000000000000000;
	sram_mem[103053] = 16'b0000000000000000;
	sram_mem[103054] = 16'b0000000000000000;
	sram_mem[103055] = 16'b0000000000000000;
	sram_mem[103056] = 16'b0000000000000000;
	sram_mem[103057] = 16'b0000000000000000;
	sram_mem[103058] = 16'b0000000000000000;
	sram_mem[103059] = 16'b0000000000000000;
	sram_mem[103060] = 16'b0000000000000000;
	sram_mem[103061] = 16'b0000000000000000;
	sram_mem[103062] = 16'b0000000000000000;
	sram_mem[103063] = 16'b0000000000000000;
	sram_mem[103064] = 16'b0000000000000000;
	sram_mem[103065] = 16'b0000000000000000;
	sram_mem[103066] = 16'b0000000000000000;
	sram_mem[103067] = 16'b0000000000000000;
	sram_mem[103068] = 16'b0000000000000000;
	sram_mem[103069] = 16'b0000000000000000;
	sram_mem[103070] = 16'b0000000000000000;
	sram_mem[103071] = 16'b0000000000000000;
	sram_mem[103072] = 16'b0000000000000000;
	sram_mem[103073] = 16'b0000000000000000;
	sram_mem[103074] = 16'b0000000000000000;
	sram_mem[103075] = 16'b0000000000000000;
	sram_mem[103076] = 16'b0000000000000000;
	sram_mem[103077] = 16'b0000000000000000;
	sram_mem[103078] = 16'b0000000000000000;
	sram_mem[103079] = 16'b0000000000000000;
	sram_mem[103080] = 16'b0000000000000000;
	sram_mem[103081] = 16'b0000000000000000;
	sram_mem[103082] = 16'b0000000000000000;
	sram_mem[103083] = 16'b0000000000000000;
	sram_mem[103084] = 16'b0000000000000000;
	sram_mem[103085] = 16'b0000000000000000;
	sram_mem[103086] = 16'b0000000000000000;
	sram_mem[103087] = 16'b0000000000000000;
	sram_mem[103088] = 16'b0000000000000000;
	sram_mem[103089] = 16'b0000000000000000;
	sram_mem[103090] = 16'b0000000000000000;
	sram_mem[103091] = 16'b0000000000000000;
	sram_mem[103092] = 16'b0000000000000000;
	sram_mem[103093] = 16'b0000000000000000;
	sram_mem[103094] = 16'b0000000000000000;
	sram_mem[103095] = 16'b0000000000000000;
	sram_mem[103096] = 16'b0000000000000000;
	sram_mem[103097] = 16'b0000000000000000;
	sram_mem[103098] = 16'b0000000000000000;
	sram_mem[103099] = 16'b0000000000000000;
	sram_mem[103100] = 16'b0000000000000000;
	sram_mem[103101] = 16'b0000000000000000;
	sram_mem[103102] = 16'b0000000000000000;
	sram_mem[103103] = 16'b0000000000000000;
	sram_mem[103104] = 16'b0000000000000000;
	sram_mem[103105] = 16'b0000000000000000;
	sram_mem[103106] = 16'b0000000000000000;
	sram_mem[103107] = 16'b0000000000000000;
	sram_mem[103108] = 16'b0000000000000000;
	sram_mem[103109] = 16'b0000000000000000;
	sram_mem[103110] = 16'b0000000000000000;
	sram_mem[103111] = 16'b0000000000000000;
	sram_mem[103112] = 16'b0000000000000000;
	sram_mem[103113] = 16'b0000000000000000;
	sram_mem[103114] = 16'b0000000000000000;
	sram_mem[103115] = 16'b0000000000000000;
	sram_mem[103116] = 16'b0000000000000000;
	sram_mem[103117] = 16'b0000000000000000;
	sram_mem[103118] = 16'b0000000000000000;
	sram_mem[103119] = 16'b0000000000000000;
	sram_mem[103120] = 16'b0000000000000000;
	sram_mem[103121] = 16'b0000000000000000;
	sram_mem[103122] = 16'b0000000000000000;
	sram_mem[103123] = 16'b0000000000000000;
	sram_mem[103124] = 16'b0000000000000000;
	sram_mem[103125] = 16'b0000000000000000;
	sram_mem[103126] = 16'b0000000000000000;
	sram_mem[103127] = 16'b0000000000000000;
	sram_mem[103128] = 16'b0000000000000000;
	sram_mem[103129] = 16'b0000000000000000;
	sram_mem[103130] = 16'b0000000000000000;
	sram_mem[103131] = 16'b0000000000000000;
	sram_mem[103132] = 16'b0000000000000000;
	sram_mem[103133] = 16'b0000000000000000;
	sram_mem[103134] = 16'b0000000000000000;
	sram_mem[103135] = 16'b0000000000000000;
	sram_mem[103136] = 16'b0000000000000000;
	sram_mem[103137] = 16'b0000000000000000;
	sram_mem[103138] = 16'b0000000000000000;
	sram_mem[103139] = 16'b0000000000000000;
	sram_mem[103140] = 16'b0000000000000000;
	sram_mem[103141] = 16'b0000000000000000;
	sram_mem[103142] = 16'b0000000000000000;
	sram_mem[103143] = 16'b0000000000000000;
	sram_mem[103144] = 16'b0000000000000000;
	sram_mem[103145] = 16'b0000000000000000;
	sram_mem[103146] = 16'b0000000000000000;
	sram_mem[103147] = 16'b0000000000000000;
	sram_mem[103148] = 16'b0000000000000000;
	sram_mem[103149] = 16'b0000000000000000;
	sram_mem[103150] = 16'b0000000000000000;
	sram_mem[103151] = 16'b0000000000000000;
	sram_mem[103152] = 16'b0000000000000000;
	sram_mem[103153] = 16'b0000000000000000;
	sram_mem[103154] = 16'b0000000000000000;
	sram_mem[103155] = 16'b0000000000000000;
	sram_mem[103156] = 16'b0000000000000000;
	sram_mem[103157] = 16'b0000000000000000;
	sram_mem[103158] = 16'b0000000000000000;
	sram_mem[103159] = 16'b0000000000000000;
	sram_mem[103160] = 16'b0000000000000000;
	sram_mem[103161] = 16'b0000000000000000;
	sram_mem[103162] = 16'b0000000000000000;
	sram_mem[103163] = 16'b0000000000000000;
	sram_mem[103164] = 16'b0000000000000000;
	sram_mem[103165] = 16'b0000000000000000;
	sram_mem[103166] = 16'b0000000000000000;
	sram_mem[103167] = 16'b0000000000000000;
	sram_mem[103168] = 16'b0000000000000000;
	sram_mem[103169] = 16'b0000000000000000;
	sram_mem[103170] = 16'b0000000000000000;
	sram_mem[103171] = 16'b0000000000000000;
	sram_mem[103172] = 16'b0000000000000000;
	sram_mem[103173] = 16'b0000000000000000;
	sram_mem[103174] = 16'b0000000000000000;
	sram_mem[103175] = 16'b0000000000000000;
	sram_mem[103176] = 16'b0000000000000000;
	sram_mem[103177] = 16'b0000000000000000;
	sram_mem[103178] = 16'b0000000000000000;
	sram_mem[103179] = 16'b0000000000000000;
	sram_mem[103180] = 16'b0000000000000000;
	sram_mem[103181] = 16'b0000000000000000;
	sram_mem[103182] = 16'b0000000000000000;
	sram_mem[103183] = 16'b0000000000000000;
	sram_mem[103184] = 16'b0000000000000000;
	sram_mem[103185] = 16'b0000000000000000;
	sram_mem[103186] = 16'b0000000000000000;
	sram_mem[103187] = 16'b0000000000000000;
	sram_mem[103188] = 16'b0000000000000000;
	sram_mem[103189] = 16'b0000000000000000;
	sram_mem[103190] = 16'b0000000000000000;
	sram_mem[103191] = 16'b0000000000000000;
	sram_mem[103192] = 16'b0000000000000000;
	sram_mem[103193] = 16'b0000000000000000;
	sram_mem[103194] = 16'b0000000000000000;
	sram_mem[103195] = 16'b0000000000000000;
	sram_mem[103196] = 16'b0000000000000000;
	sram_mem[103197] = 16'b0000000000000000;
	sram_mem[103198] = 16'b0000000000000000;
	sram_mem[103199] = 16'b0000000000000000;
	sram_mem[103200] = 16'b0000000000000000;
	sram_mem[103201] = 16'b0000000000000000;
	sram_mem[103202] = 16'b0000000000000000;
	sram_mem[103203] = 16'b0000000000000000;
	sram_mem[103204] = 16'b0000000000000000;
	sram_mem[103205] = 16'b0000000000000000;
	sram_mem[103206] = 16'b0000000000000000;
	sram_mem[103207] = 16'b0000000000000000;
	sram_mem[103208] = 16'b0000000000000000;
	sram_mem[103209] = 16'b0000000000000000;
	sram_mem[103210] = 16'b0000000000000000;
	sram_mem[103211] = 16'b0000000000000000;
	sram_mem[103212] = 16'b0000000000000000;
	sram_mem[103213] = 16'b0000000000000000;
	sram_mem[103214] = 16'b0000000000000000;
	sram_mem[103215] = 16'b0000000000000000;
	sram_mem[103216] = 16'b0000000000000000;
	sram_mem[103217] = 16'b0000000000000000;
	sram_mem[103218] = 16'b0000000000000000;
	sram_mem[103219] = 16'b0000000000000000;
	sram_mem[103220] = 16'b0000000000000000;
	sram_mem[103221] = 16'b0000000000000000;
	sram_mem[103222] = 16'b0000000000000000;
	sram_mem[103223] = 16'b0000000000000000;
	sram_mem[103224] = 16'b0000000000000000;
	sram_mem[103225] = 16'b0000000000000000;
	sram_mem[103226] = 16'b0000000000000000;
	sram_mem[103227] = 16'b0000000000000000;
	sram_mem[103228] = 16'b0000000000000000;
	sram_mem[103229] = 16'b0000000000000000;
	sram_mem[103230] = 16'b0000000000000000;
	sram_mem[103231] = 16'b0000000000000000;
	sram_mem[103232] = 16'b0000000000000000;
	sram_mem[103233] = 16'b0000000000000000;
	sram_mem[103234] = 16'b0000000000000000;
	sram_mem[103235] = 16'b0000000000000000;
	sram_mem[103236] = 16'b0000000000000000;
	sram_mem[103237] = 16'b0000000000000000;
	sram_mem[103238] = 16'b0000000000000000;
	sram_mem[103239] = 16'b0000000000000000;
	sram_mem[103240] = 16'b0000000000000000;
	sram_mem[103241] = 16'b0000000000000000;
	sram_mem[103242] = 16'b0000000000000000;
	sram_mem[103243] = 16'b0000000000000000;
	sram_mem[103244] = 16'b0000000000000000;
	sram_mem[103245] = 16'b0000000000000000;
	sram_mem[103246] = 16'b0000000000000000;
	sram_mem[103247] = 16'b0000000000000000;
	sram_mem[103248] = 16'b0000000000000000;
	sram_mem[103249] = 16'b0000000000000000;
	sram_mem[103250] = 16'b0000000000000000;
	sram_mem[103251] = 16'b0000000000000000;
	sram_mem[103252] = 16'b0000000000000000;
	sram_mem[103253] = 16'b0000000000000000;
	sram_mem[103254] = 16'b0000000000000000;
	sram_mem[103255] = 16'b0000000000000000;
	sram_mem[103256] = 16'b0000000000000000;
	sram_mem[103257] = 16'b0000000000000000;
	sram_mem[103258] = 16'b0000000000000000;
	sram_mem[103259] = 16'b0000000000000000;
	sram_mem[103260] = 16'b0000000000000000;
	sram_mem[103261] = 16'b0000000000000000;
	sram_mem[103262] = 16'b0000000000000000;
	sram_mem[103263] = 16'b0000000000000000;
	sram_mem[103264] = 16'b0000000000000000;
	sram_mem[103265] = 16'b0000000000000000;
	sram_mem[103266] = 16'b0000000000000000;
	sram_mem[103267] = 16'b0000000000000000;
	sram_mem[103268] = 16'b0000000000000000;
	sram_mem[103269] = 16'b0000000000000000;
	sram_mem[103270] = 16'b0000000000000000;
	sram_mem[103271] = 16'b0000000000000000;
	sram_mem[103272] = 16'b0000000000000000;
	sram_mem[103273] = 16'b0000000000000000;
	sram_mem[103274] = 16'b0000000000000000;
	sram_mem[103275] = 16'b0000000000000000;
	sram_mem[103276] = 16'b0000000000000000;
	sram_mem[103277] = 16'b0000000000000000;
	sram_mem[103278] = 16'b0000000000000000;
	sram_mem[103279] = 16'b0000000000000000;
	sram_mem[103280] = 16'b0000000000000000;
	sram_mem[103281] = 16'b0000000000000000;
	sram_mem[103282] = 16'b0000000000000000;
	sram_mem[103283] = 16'b0000000000000000;
	sram_mem[103284] = 16'b0000000000000000;
	sram_mem[103285] = 16'b0000000000000000;
	sram_mem[103286] = 16'b0000000000000000;
	sram_mem[103287] = 16'b0000000000000000;
	sram_mem[103288] = 16'b0000000000000000;
	sram_mem[103289] = 16'b0000000000000000;
	sram_mem[103290] = 16'b0000000000000000;
	sram_mem[103291] = 16'b0000000000000000;
	sram_mem[103292] = 16'b0000000000000000;
	sram_mem[103293] = 16'b0000000000000000;
	sram_mem[103294] = 16'b0000000000000000;
	sram_mem[103295] = 16'b0000000000000000;
	sram_mem[103296] = 16'b0000000000000000;
	sram_mem[103297] = 16'b0000000000000000;
	sram_mem[103298] = 16'b0000000000000000;
	sram_mem[103299] = 16'b0000000000000000;
	sram_mem[103300] = 16'b0000000000000000;
	sram_mem[103301] = 16'b0000000000000000;
	sram_mem[103302] = 16'b0000000000000000;
	sram_mem[103303] = 16'b0000000000000000;
	sram_mem[103304] = 16'b0000000000000000;
	sram_mem[103305] = 16'b0000000000000000;
	sram_mem[103306] = 16'b0000000000000000;
	sram_mem[103307] = 16'b0000000000000000;
	sram_mem[103308] = 16'b0000000000000000;
	sram_mem[103309] = 16'b0000000000000000;
	sram_mem[103310] = 16'b0000000000000000;
	sram_mem[103311] = 16'b0000000000000000;
	sram_mem[103312] = 16'b0000000000000000;
	sram_mem[103313] = 16'b0000000000000000;
	sram_mem[103314] = 16'b0000000000000000;
	sram_mem[103315] = 16'b0000000000000000;
	sram_mem[103316] = 16'b0000000000000000;
	sram_mem[103317] = 16'b0000000000000000;
	sram_mem[103318] = 16'b0000000000000000;
	sram_mem[103319] = 16'b0000000000000000;
	sram_mem[103320] = 16'b0000000000000000;
	sram_mem[103321] = 16'b0000000000000000;
	sram_mem[103322] = 16'b0000000000000000;
	sram_mem[103323] = 16'b0000000000000000;
	sram_mem[103324] = 16'b0000000000000000;
	sram_mem[103325] = 16'b0000000000000000;
	sram_mem[103326] = 16'b0000000000000000;
	sram_mem[103327] = 16'b0000000000000000;
	sram_mem[103328] = 16'b0000000000000000;
	sram_mem[103329] = 16'b0000000000000000;
	sram_mem[103330] = 16'b0000000000000000;
	sram_mem[103331] = 16'b0000000000000000;
	sram_mem[103332] = 16'b0000000000000000;
	sram_mem[103333] = 16'b0000000000000000;
	sram_mem[103334] = 16'b0000000000000000;
	sram_mem[103335] = 16'b0000000000000000;
	sram_mem[103336] = 16'b0000000000000000;
	sram_mem[103337] = 16'b0000000000000000;
	sram_mem[103338] = 16'b0000000000000000;
	sram_mem[103339] = 16'b0000000000000000;
	sram_mem[103340] = 16'b0000000000000000;
	sram_mem[103341] = 16'b0000000000000000;
	sram_mem[103342] = 16'b0000000000000000;
	sram_mem[103343] = 16'b0000000000000000;
	sram_mem[103344] = 16'b0000000000000000;
	sram_mem[103345] = 16'b0000000000000000;
	sram_mem[103346] = 16'b0000000000000000;
	sram_mem[103347] = 16'b0000000000000000;
	sram_mem[103348] = 16'b0000000000000000;
	sram_mem[103349] = 16'b0000000000000000;
	sram_mem[103350] = 16'b0000000000000000;
	sram_mem[103351] = 16'b0000000000000000;
	sram_mem[103352] = 16'b0000000000000000;
	sram_mem[103353] = 16'b0000000000000000;
	sram_mem[103354] = 16'b0000000000000000;
	sram_mem[103355] = 16'b0000000000000000;
	sram_mem[103356] = 16'b0000000000000000;
	sram_mem[103357] = 16'b0000000000000000;
	sram_mem[103358] = 16'b0000000000000000;
	sram_mem[103359] = 16'b0000000000000000;
	sram_mem[103360] = 16'b0000000000000000;
	sram_mem[103361] = 16'b0000000000000000;
	sram_mem[103362] = 16'b0000000000000000;
	sram_mem[103363] = 16'b0000000000000000;
	sram_mem[103364] = 16'b0000000000000000;
	sram_mem[103365] = 16'b0000000000000000;
	sram_mem[103366] = 16'b0000000000000000;
	sram_mem[103367] = 16'b0000000000000000;
	sram_mem[103368] = 16'b0000000000000000;
	sram_mem[103369] = 16'b0000000000000000;
	sram_mem[103370] = 16'b0000000000000000;
	sram_mem[103371] = 16'b0000000000000000;
	sram_mem[103372] = 16'b0000000000000000;
	sram_mem[103373] = 16'b0000000000000000;
	sram_mem[103374] = 16'b0000000000000000;
	sram_mem[103375] = 16'b0000000000000000;
	sram_mem[103376] = 16'b0000000000000000;
	sram_mem[103377] = 16'b0000000000000000;
	sram_mem[103378] = 16'b0000000000000000;
	sram_mem[103379] = 16'b0000000000000000;
	sram_mem[103380] = 16'b0000000000000000;
	sram_mem[103381] = 16'b0000000000000000;
	sram_mem[103382] = 16'b0000000000000000;
	sram_mem[103383] = 16'b0000000000000000;
	sram_mem[103384] = 16'b0000000000000000;
	sram_mem[103385] = 16'b0000000000000000;
	sram_mem[103386] = 16'b0000000000000000;
	sram_mem[103387] = 16'b0000000000000000;
	sram_mem[103388] = 16'b0000000000000000;
	sram_mem[103389] = 16'b0000000000000000;
	sram_mem[103390] = 16'b0000000000000000;
	sram_mem[103391] = 16'b0000000000000000;
	sram_mem[103392] = 16'b0000000000000000;
	sram_mem[103393] = 16'b0000000000000000;
	sram_mem[103394] = 16'b0000000000000000;
	sram_mem[103395] = 16'b0000000000000000;
	sram_mem[103396] = 16'b0000000000000000;
	sram_mem[103397] = 16'b0000000000000000;
	sram_mem[103398] = 16'b0000000000000000;
	sram_mem[103399] = 16'b0000000000000000;
	sram_mem[103400] = 16'b0000000000000000;
	sram_mem[103401] = 16'b0000000000000000;
	sram_mem[103402] = 16'b0000000000000000;
	sram_mem[103403] = 16'b0000000000000000;
	sram_mem[103404] = 16'b0000000000000000;
	sram_mem[103405] = 16'b0000000000000000;
	sram_mem[103406] = 16'b0000000000000000;
	sram_mem[103407] = 16'b0000000000000000;
	sram_mem[103408] = 16'b0000000000000000;
	sram_mem[103409] = 16'b0000000000000000;
	sram_mem[103410] = 16'b0000000000000000;
	sram_mem[103411] = 16'b0000000000000000;
	sram_mem[103412] = 16'b0000000000000000;
	sram_mem[103413] = 16'b0000000000000000;
	sram_mem[103414] = 16'b0000000000000000;
	sram_mem[103415] = 16'b0000000000000000;
	sram_mem[103416] = 16'b0000000000000000;
	sram_mem[103417] = 16'b0000000000000000;
	sram_mem[103418] = 16'b0000000000000000;
	sram_mem[103419] = 16'b0000000000000000;
	sram_mem[103420] = 16'b0000000000000000;
	sram_mem[103421] = 16'b0000000000000000;
	sram_mem[103422] = 16'b0000000000000000;
	sram_mem[103423] = 16'b0000000000000000;
	sram_mem[103424] = 16'b0000000000000000;
	sram_mem[103425] = 16'b0000000000000000;
	sram_mem[103426] = 16'b0000000000000000;
	sram_mem[103427] = 16'b0000000000000000;
	sram_mem[103428] = 16'b0000000000000000;
	sram_mem[103429] = 16'b0000000000000000;
	sram_mem[103430] = 16'b0000000000000000;
	sram_mem[103431] = 16'b0000000000000000;
	sram_mem[103432] = 16'b0000000000000000;
	sram_mem[103433] = 16'b0000000000000000;
	sram_mem[103434] = 16'b0000000000000000;
	sram_mem[103435] = 16'b0000000000000000;
	sram_mem[103436] = 16'b0000000000000000;
	sram_mem[103437] = 16'b0000000000000000;
	sram_mem[103438] = 16'b0000000000000000;
	sram_mem[103439] = 16'b0000000000000000;
	sram_mem[103440] = 16'b0000000000000000;
	sram_mem[103441] = 16'b0000000000000000;
	sram_mem[103442] = 16'b0000000000000000;
	sram_mem[103443] = 16'b0000000000000000;
	sram_mem[103444] = 16'b0000000000000000;
	sram_mem[103445] = 16'b0000000000000000;
	sram_mem[103446] = 16'b0000000000000000;
	sram_mem[103447] = 16'b0000000000000000;
	sram_mem[103448] = 16'b0000000000000000;
	sram_mem[103449] = 16'b0000000000000000;
	sram_mem[103450] = 16'b0000000000000000;
	sram_mem[103451] = 16'b0000000000000000;
	sram_mem[103452] = 16'b0000000000000000;
	sram_mem[103453] = 16'b0000000000000000;
	sram_mem[103454] = 16'b0000000000000000;
	sram_mem[103455] = 16'b0000000000000000;
	sram_mem[103456] = 16'b0000000000000000;
	sram_mem[103457] = 16'b0000000000000000;
	sram_mem[103458] = 16'b0000000000000000;
	sram_mem[103459] = 16'b0000000000000000;
	sram_mem[103460] = 16'b0000000000000000;
	sram_mem[103461] = 16'b0000000000000000;
	sram_mem[103462] = 16'b0000000000000000;
	sram_mem[103463] = 16'b0000000000000000;
	sram_mem[103464] = 16'b0000000000000000;
	sram_mem[103465] = 16'b0000000000000000;
	sram_mem[103466] = 16'b0000000000000000;
	sram_mem[103467] = 16'b0000000000000000;
	sram_mem[103468] = 16'b0000000000000000;
	sram_mem[103469] = 16'b0000000000000000;
	sram_mem[103470] = 16'b0000000000000000;
	sram_mem[103471] = 16'b0000000000000000;
	sram_mem[103472] = 16'b0000000000000000;
	sram_mem[103473] = 16'b0000000000000000;
	sram_mem[103474] = 16'b0000000000000000;
	sram_mem[103475] = 16'b0000000000000000;
	sram_mem[103476] = 16'b0000000000000000;
	sram_mem[103477] = 16'b0000000000000000;
	sram_mem[103478] = 16'b0000000000000000;
	sram_mem[103479] = 16'b0000000000000000;
	sram_mem[103480] = 16'b0000000000000000;
	sram_mem[103481] = 16'b0000000000000000;
	sram_mem[103482] = 16'b0000000000000000;
	sram_mem[103483] = 16'b0000000000000000;
	sram_mem[103484] = 16'b0000000000000000;
	sram_mem[103485] = 16'b0000000000000000;
	sram_mem[103486] = 16'b0000000000000000;
	sram_mem[103487] = 16'b0000000000000000;
	sram_mem[103488] = 16'b0000000000000000;
	sram_mem[103489] = 16'b0000000000000000;
	sram_mem[103490] = 16'b0000000000000000;
	sram_mem[103491] = 16'b0000000000000000;
	sram_mem[103492] = 16'b0000000000000000;
	sram_mem[103493] = 16'b0000000000000000;
	sram_mem[103494] = 16'b0000000000000000;
	sram_mem[103495] = 16'b0000000000000000;
	sram_mem[103496] = 16'b0000000000000000;
	sram_mem[103497] = 16'b0000000000000000;
	sram_mem[103498] = 16'b0000000000000000;
	sram_mem[103499] = 16'b0000000000000000;
	sram_mem[103500] = 16'b0000000000000000;
	sram_mem[103501] = 16'b0000000000000000;
	sram_mem[103502] = 16'b0000000000000000;
	sram_mem[103503] = 16'b0000000000000000;
	sram_mem[103504] = 16'b0000000000000000;
	sram_mem[103505] = 16'b0000000000000000;
	sram_mem[103506] = 16'b0000000000000000;
	sram_mem[103507] = 16'b0000000000000000;
	sram_mem[103508] = 16'b0000000000000000;
	sram_mem[103509] = 16'b0000000000000000;
	sram_mem[103510] = 16'b0000000000000000;
	sram_mem[103511] = 16'b0000000000000000;
	sram_mem[103512] = 16'b0000000000000000;
	sram_mem[103513] = 16'b0000000000000000;
	sram_mem[103514] = 16'b0000000000000000;
	sram_mem[103515] = 16'b0000000000000000;
	sram_mem[103516] = 16'b0000000000000000;
	sram_mem[103517] = 16'b0000000000000000;
	sram_mem[103518] = 16'b0000000000000000;
	sram_mem[103519] = 16'b0000000000000000;
	sram_mem[103520] = 16'b0000000000000000;
	sram_mem[103521] = 16'b0000000000000000;
	sram_mem[103522] = 16'b0000000000000000;
	sram_mem[103523] = 16'b0000000000000000;
	sram_mem[103524] = 16'b0000000000000000;
	sram_mem[103525] = 16'b0000000000000000;
	sram_mem[103526] = 16'b0000000000000000;
	sram_mem[103527] = 16'b0000000000000000;
	sram_mem[103528] = 16'b0000000000000000;
	sram_mem[103529] = 16'b0000000000000000;
	sram_mem[103530] = 16'b0000000000000000;
	sram_mem[103531] = 16'b0000000000000000;
	sram_mem[103532] = 16'b0000000000000000;
	sram_mem[103533] = 16'b0000000000000000;
	sram_mem[103534] = 16'b0000000000000000;
	sram_mem[103535] = 16'b0000000000000000;
	sram_mem[103536] = 16'b0000000000000000;
	sram_mem[103537] = 16'b0000000000000000;
	sram_mem[103538] = 16'b0000000000000000;
	sram_mem[103539] = 16'b0000000000000000;
	sram_mem[103540] = 16'b0000000000000000;
	sram_mem[103541] = 16'b0000000000000000;
	sram_mem[103542] = 16'b0000000000000000;
	sram_mem[103543] = 16'b0000000000000000;
	sram_mem[103544] = 16'b0000000000000000;
	sram_mem[103545] = 16'b0000000000000000;
	sram_mem[103546] = 16'b0000000000000000;
	sram_mem[103547] = 16'b0000000000000000;
	sram_mem[103548] = 16'b0000000000000000;
	sram_mem[103549] = 16'b0000000000000000;
	sram_mem[103550] = 16'b0000000000000000;
	sram_mem[103551] = 16'b0000000000000000;
	sram_mem[103552] = 16'b0000000000000000;
	sram_mem[103553] = 16'b0000000000000000;
	sram_mem[103554] = 16'b0000000000000000;
	sram_mem[103555] = 16'b0000000000000000;
	sram_mem[103556] = 16'b0000000000000000;
	sram_mem[103557] = 16'b0000000000000000;
	sram_mem[103558] = 16'b0000000000000000;
	sram_mem[103559] = 16'b0000000000000000;
	sram_mem[103560] = 16'b0000000000000000;
	sram_mem[103561] = 16'b0000000000000000;
	sram_mem[103562] = 16'b0000000000000000;
	sram_mem[103563] = 16'b0000000000000000;
	sram_mem[103564] = 16'b0000000000000000;
	sram_mem[103565] = 16'b0000000000000000;
	sram_mem[103566] = 16'b0000000000000000;
	sram_mem[103567] = 16'b0000000000000000;
	sram_mem[103568] = 16'b0000000000000000;
	sram_mem[103569] = 16'b0000000000000000;
	sram_mem[103570] = 16'b0000000000000000;
	sram_mem[103571] = 16'b0000000000000000;
	sram_mem[103572] = 16'b0000000000000000;
	sram_mem[103573] = 16'b0000000000000000;
	sram_mem[103574] = 16'b0000000000000000;
	sram_mem[103575] = 16'b0000000000000000;
	sram_mem[103576] = 16'b0000000000000000;
	sram_mem[103577] = 16'b0000000000000000;
	sram_mem[103578] = 16'b0000000000000000;
	sram_mem[103579] = 16'b0000000000000000;
	sram_mem[103580] = 16'b0000000000000000;
	sram_mem[103581] = 16'b0000000000000000;
	sram_mem[103582] = 16'b0000000000000000;
	sram_mem[103583] = 16'b0000000000000000;
	sram_mem[103584] = 16'b0000000000000000;
	sram_mem[103585] = 16'b0000000000000000;
	sram_mem[103586] = 16'b0000000000000000;
	sram_mem[103587] = 16'b0000000000000000;
	sram_mem[103588] = 16'b0000000000000000;
	sram_mem[103589] = 16'b0000000000000000;
	sram_mem[103590] = 16'b0000000000000000;
	sram_mem[103591] = 16'b0000000000000000;
	sram_mem[103592] = 16'b0000000000000000;
	sram_mem[103593] = 16'b0000000000000000;
	sram_mem[103594] = 16'b0000000000000000;
	sram_mem[103595] = 16'b0000000000000000;
	sram_mem[103596] = 16'b0000000000000000;
	sram_mem[103597] = 16'b0000000000000000;
	sram_mem[103598] = 16'b0000000000000000;
	sram_mem[103599] = 16'b0000000000000000;
	sram_mem[103600] = 16'b0000000000000000;
	sram_mem[103601] = 16'b0000000000000000;
	sram_mem[103602] = 16'b0000000000000000;
	sram_mem[103603] = 16'b0000000000000000;
	sram_mem[103604] = 16'b0000000000000000;
	sram_mem[103605] = 16'b0000000000000000;
	sram_mem[103606] = 16'b0000000000000000;
	sram_mem[103607] = 16'b0000000000000000;
	sram_mem[103608] = 16'b0000000000000000;
	sram_mem[103609] = 16'b0000000000000000;
	sram_mem[103610] = 16'b0000000000000000;
	sram_mem[103611] = 16'b0000000000000000;
	sram_mem[103612] = 16'b0000000000000000;
	sram_mem[103613] = 16'b0000000000000000;
	sram_mem[103614] = 16'b0000000000000000;
	sram_mem[103615] = 16'b0000000000000000;
	sram_mem[103616] = 16'b0000000000000000;
	sram_mem[103617] = 16'b0000000000000000;
	sram_mem[103618] = 16'b0000000000000000;
	sram_mem[103619] = 16'b0000000000000000;
	sram_mem[103620] = 16'b0000000000000000;
	sram_mem[103621] = 16'b0000000000000000;
	sram_mem[103622] = 16'b0000000000000000;
	sram_mem[103623] = 16'b0000000000000000;
	sram_mem[103624] = 16'b0000000000000000;
	sram_mem[103625] = 16'b0000000000000000;
	sram_mem[103626] = 16'b0000000000000000;
	sram_mem[103627] = 16'b0000000000000000;
	sram_mem[103628] = 16'b0000000000000000;
	sram_mem[103629] = 16'b0000000000000000;
	sram_mem[103630] = 16'b0000000000000000;
	sram_mem[103631] = 16'b0000000000000000;
	sram_mem[103632] = 16'b0000000000000000;
	sram_mem[103633] = 16'b0000000000000000;
	sram_mem[103634] = 16'b0000000000000000;
	sram_mem[103635] = 16'b0000000000000000;
	sram_mem[103636] = 16'b0000000000000000;
	sram_mem[103637] = 16'b0000000000000000;
	sram_mem[103638] = 16'b0000000000000000;
	sram_mem[103639] = 16'b0000000000000000;
	sram_mem[103640] = 16'b0000000000000000;
	sram_mem[103641] = 16'b0000000000000000;
	sram_mem[103642] = 16'b0000000000000000;
	sram_mem[103643] = 16'b0000000000000000;
	sram_mem[103644] = 16'b0000000000000000;
	sram_mem[103645] = 16'b0000000000000000;
	sram_mem[103646] = 16'b0000000000000000;
	sram_mem[103647] = 16'b0000000000000000;
	sram_mem[103648] = 16'b0000000000000000;
	sram_mem[103649] = 16'b0000000000000000;
	sram_mem[103650] = 16'b0000000000000000;
	sram_mem[103651] = 16'b0000000000000000;
	sram_mem[103652] = 16'b0000000000000000;
	sram_mem[103653] = 16'b0000000000000000;
	sram_mem[103654] = 16'b0000000000000000;
	sram_mem[103655] = 16'b0000000000000000;
	sram_mem[103656] = 16'b0000000000000000;
	sram_mem[103657] = 16'b0000000000000000;
	sram_mem[103658] = 16'b0000000000000000;
	sram_mem[103659] = 16'b0000000000000000;
	sram_mem[103660] = 16'b0000000000000000;
	sram_mem[103661] = 16'b0000000000000000;
	sram_mem[103662] = 16'b0000000000000000;
	sram_mem[103663] = 16'b0000000000000000;
	sram_mem[103664] = 16'b0000000000000000;
	sram_mem[103665] = 16'b0000000000000000;
	sram_mem[103666] = 16'b0000000000000000;
	sram_mem[103667] = 16'b0000000000000000;
	sram_mem[103668] = 16'b0000000000000000;
	sram_mem[103669] = 16'b0000000000000000;
	sram_mem[103670] = 16'b0000000000000000;
	sram_mem[103671] = 16'b0000000000000000;
	sram_mem[103672] = 16'b0000000000000000;
	sram_mem[103673] = 16'b0000000000000000;
	sram_mem[103674] = 16'b0000000000000000;
	sram_mem[103675] = 16'b0000000000000000;
	sram_mem[103676] = 16'b0000000000000000;
	sram_mem[103677] = 16'b0000000000000000;
	sram_mem[103678] = 16'b0000000000000000;
	sram_mem[103679] = 16'b0000000000000000;
	sram_mem[103680] = 16'b0000000000000000;
	sram_mem[103681] = 16'b0000000000000000;
	sram_mem[103682] = 16'b0000000000000000;
	sram_mem[103683] = 16'b0000000000000000;
	sram_mem[103684] = 16'b0000000000000000;
	sram_mem[103685] = 16'b0000000000000000;
	sram_mem[103686] = 16'b0000000000000000;
	sram_mem[103687] = 16'b0000000000000000;
	sram_mem[103688] = 16'b0000000000000000;
	sram_mem[103689] = 16'b0000000000000000;
	sram_mem[103690] = 16'b0000000000000000;
	sram_mem[103691] = 16'b0000000000000000;
	sram_mem[103692] = 16'b0000000000000000;
	sram_mem[103693] = 16'b0000000000000000;
	sram_mem[103694] = 16'b0000000000000000;
	sram_mem[103695] = 16'b0000000000000000;
	sram_mem[103696] = 16'b0000000000000000;
	sram_mem[103697] = 16'b0000000000000000;
	sram_mem[103698] = 16'b0000000000000000;
	sram_mem[103699] = 16'b0000000000000000;
	sram_mem[103700] = 16'b0000000000000000;
	sram_mem[103701] = 16'b0000000000000000;
	sram_mem[103702] = 16'b0000000000000000;
	sram_mem[103703] = 16'b0000000000000000;
	sram_mem[103704] = 16'b0000000000000000;
	sram_mem[103705] = 16'b0000000000000000;
	sram_mem[103706] = 16'b0000000000000000;
	sram_mem[103707] = 16'b0000000000000000;
	sram_mem[103708] = 16'b0000000000000000;
	sram_mem[103709] = 16'b0000000000000000;
	sram_mem[103710] = 16'b0000000000000000;
	sram_mem[103711] = 16'b0000000000000000;
	sram_mem[103712] = 16'b0000000000000000;
	sram_mem[103713] = 16'b0000000000000000;
	sram_mem[103714] = 16'b0000000000000000;
	sram_mem[103715] = 16'b0000000000000000;
	sram_mem[103716] = 16'b0000000000000000;
	sram_mem[103717] = 16'b0000000000000000;
	sram_mem[103718] = 16'b0000000000000000;
	sram_mem[103719] = 16'b0000000000000000;
	sram_mem[103720] = 16'b0000000000000000;
	sram_mem[103721] = 16'b0000000000000000;
	sram_mem[103722] = 16'b0000000000000000;
	sram_mem[103723] = 16'b0000000000000000;
	sram_mem[103724] = 16'b0000000000000000;
	sram_mem[103725] = 16'b0000000000000000;
	sram_mem[103726] = 16'b0000000000000000;
	sram_mem[103727] = 16'b0000000000000000;
	sram_mem[103728] = 16'b0000000000000000;
	sram_mem[103729] = 16'b0000000000000000;
	sram_mem[103730] = 16'b0000000000000000;
	sram_mem[103731] = 16'b0000000000000000;
	sram_mem[103732] = 16'b0000000000000000;
	sram_mem[103733] = 16'b0000000000000000;
	sram_mem[103734] = 16'b0000000000000000;
	sram_mem[103735] = 16'b0000000000000000;
	sram_mem[103736] = 16'b0000000000000000;
	sram_mem[103737] = 16'b0000000000000000;
	sram_mem[103738] = 16'b0000000000000000;
	sram_mem[103739] = 16'b0000000000000000;
	sram_mem[103740] = 16'b0000000000000000;
	sram_mem[103741] = 16'b0000000000000000;
	sram_mem[103742] = 16'b0000000000000000;
	sram_mem[103743] = 16'b0000000000000000;
	sram_mem[103744] = 16'b0000000000000000;
	sram_mem[103745] = 16'b0000000000000000;
	sram_mem[103746] = 16'b0000000000000000;
	sram_mem[103747] = 16'b0000000000000000;
	sram_mem[103748] = 16'b0000000000000000;
	sram_mem[103749] = 16'b0000000000000000;
	sram_mem[103750] = 16'b0000000000000000;
	sram_mem[103751] = 16'b0000000000000000;
	sram_mem[103752] = 16'b0000000000000000;
	sram_mem[103753] = 16'b0000000000000000;
	sram_mem[103754] = 16'b0000000000000000;
	sram_mem[103755] = 16'b0000000000000000;
	sram_mem[103756] = 16'b0000000000000000;
	sram_mem[103757] = 16'b0000000000000000;
	sram_mem[103758] = 16'b0000000000000000;
	sram_mem[103759] = 16'b0000000000000000;
	sram_mem[103760] = 16'b0000000000000000;
	sram_mem[103761] = 16'b0000000000000000;
	sram_mem[103762] = 16'b0000000000000000;
	sram_mem[103763] = 16'b0000000000000000;
	sram_mem[103764] = 16'b0000000000000000;
	sram_mem[103765] = 16'b0000000000000000;
	sram_mem[103766] = 16'b0000000000000000;
	sram_mem[103767] = 16'b0000000000000000;
	sram_mem[103768] = 16'b0000000000000000;
	sram_mem[103769] = 16'b0000000000000000;
	sram_mem[103770] = 16'b0000000000000000;
	sram_mem[103771] = 16'b0000000000000000;
	sram_mem[103772] = 16'b0000000000000000;
	sram_mem[103773] = 16'b0000000000000000;
	sram_mem[103774] = 16'b0000000000000000;
	sram_mem[103775] = 16'b0000000000000000;
	sram_mem[103776] = 16'b0000000000000000;
	sram_mem[103777] = 16'b0000000000000000;
	sram_mem[103778] = 16'b0000000000000000;
	sram_mem[103779] = 16'b0000000000000000;
	sram_mem[103780] = 16'b0000000000000000;
	sram_mem[103781] = 16'b0000000000000000;
	sram_mem[103782] = 16'b0000000000000000;
	sram_mem[103783] = 16'b0000000000000000;
	sram_mem[103784] = 16'b0000000000000000;
	sram_mem[103785] = 16'b0000000000000000;
	sram_mem[103786] = 16'b0000000000000000;
	sram_mem[103787] = 16'b0000000000000000;
	sram_mem[103788] = 16'b0000000000000000;
	sram_mem[103789] = 16'b0000000000000000;
	sram_mem[103790] = 16'b0000000000000000;
	sram_mem[103791] = 16'b0000000000000000;
	sram_mem[103792] = 16'b0000000000000000;
	sram_mem[103793] = 16'b0000000000000000;
	sram_mem[103794] = 16'b0000000000000000;
	sram_mem[103795] = 16'b0000000000000000;
	sram_mem[103796] = 16'b0000000000000000;
	sram_mem[103797] = 16'b0000000000000000;
	sram_mem[103798] = 16'b0000000000000000;
	sram_mem[103799] = 16'b0000000000000000;
	sram_mem[103800] = 16'b0000000000000000;
	sram_mem[103801] = 16'b0000000000000000;
	sram_mem[103802] = 16'b0000000000000000;
	sram_mem[103803] = 16'b0000000000000000;
	sram_mem[103804] = 16'b0000000000000000;
	sram_mem[103805] = 16'b0000000000000000;
	sram_mem[103806] = 16'b0000000000000000;
	sram_mem[103807] = 16'b0000000000000000;
	sram_mem[103808] = 16'b0000000000000000;
	sram_mem[103809] = 16'b0000000000000000;
	sram_mem[103810] = 16'b0000000000000000;
	sram_mem[103811] = 16'b0000000000000000;
	sram_mem[103812] = 16'b0000000000000000;
	sram_mem[103813] = 16'b0000000000000000;
	sram_mem[103814] = 16'b0000000000000000;
	sram_mem[103815] = 16'b0000000000000000;
	sram_mem[103816] = 16'b0000000000000000;
	sram_mem[103817] = 16'b0000000000000000;
	sram_mem[103818] = 16'b0000000000000000;
	sram_mem[103819] = 16'b0000000000000000;
	sram_mem[103820] = 16'b0000000000000000;
	sram_mem[103821] = 16'b0000000000000000;
	sram_mem[103822] = 16'b0000000000000000;
	sram_mem[103823] = 16'b0000000000000000;
	sram_mem[103824] = 16'b0000000000000000;
	sram_mem[103825] = 16'b0000000000000000;
	sram_mem[103826] = 16'b0000000000000000;
	sram_mem[103827] = 16'b0000000000000000;
	sram_mem[103828] = 16'b0000000000000000;
	sram_mem[103829] = 16'b0000000000000000;
	sram_mem[103830] = 16'b0000000000000000;
	sram_mem[103831] = 16'b0000000000000000;
	sram_mem[103832] = 16'b0000000000000000;
	sram_mem[103833] = 16'b0000000000000000;
	sram_mem[103834] = 16'b0000000000000000;
	sram_mem[103835] = 16'b0000000000000000;
	sram_mem[103836] = 16'b0000000000000000;
	sram_mem[103837] = 16'b0000000000000000;
	sram_mem[103838] = 16'b0000000000000000;
	sram_mem[103839] = 16'b0000000000000000;
	sram_mem[103840] = 16'b0000000000000000;
	sram_mem[103841] = 16'b0000000000000000;
	sram_mem[103842] = 16'b0000000000000000;
	sram_mem[103843] = 16'b0000000000000000;
	sram_mem[103844] = 16'b0000000000000000;
	sram_mem[103845] = 16'b0000000000000000;
	sram_mem[103846] = 16'b0000000000000000;
	sram_mem[103847] = 16'b0000000000000000;
	sram_mem[103848] = 16'b0000000000000000;
	sram_mem[103849] = 16'b0000000000000000;
	sram_mem[103850] = 16'b0000000000000000;
	sram_mem[103851] = 16'b0000000000000000;
	sram_mem[103852] = 16'b0000000000000000;
	sram_mem[103853] = 16'b0000000000000000;
	sram_mem[103854] = 16'b0000000000000000;
	sram_mem[103855] = 16'b0000000000000000;
	sram_mem[103856] = 16'b0000000000000000;
	sram_mem[103857] = 16'b0000000000000000;
	sram_mem[103858] = 16'b0000000000000000;
	sram_mem[103859] = 16'b0000000000000000;
	sram_mem[103860] = 16'b0000000000000000;
	sram_mem[103861] = 16'b0000000000000000;
	sram_mem[103862] = 16'b0000000000000000;
	sram_mem[103863] = 16'b0000000000000000;
	sram_mem[103864] = 16'b0000000000000000;
	sram_mem[103865] = 16'b0000000000000000;
	sram_mem[103866] = 16'b0000000000000000;
	sram_mem[103867] = 16'b0000000000000000;
	sram_mem[103868] = 16'b0000000000000000;
	sram_mem[103869] = 16'b0000000000000000;
	sram_mem[103870] = 16'b0000000000000000;
	sram_mem[103871] = 16'b0000000000000000;
	sram_mem[103872] = 16'b0000000000000000;
	sram_mem[103873] = 16'b0000000000000000;
	sram_mem[103874] = 16'b0000000000000000;
	sram_mem[103875] = 16'b0000000000000000;
	sram_mem[103876] = 16'b0000000000000000;
	sram_mem[103877] = 16'b0000000000000000;
	sram_mem[103878] = 16'b0000000000000000;
	sram_mem[103879] = 16'b0000000000000000;
	sram_mem[103880] = 16'b0000000000000000;
	sram_mem[103881] = 16'b0000000000000000;
	sram_mem[103882] = 16'b0000000000000000;
	sram_mem[103883] = 16'b0000000000000000;
	sram_mem[103884] = 16'b0000000000000000;
	sram_mem[103885] = 16'b0000000000000000;
	sram_mem[103886] = 16'b0000000000000000;
	sram_mem[103887] = 16'b0000000000000000;
	sram_mem[103888] = 16'b0000000000000000;
	sram_mem[103889] = 16'b0000000000000000;
	sram_mem[103890] = 16'b0000000000000000;
	sram_mem[103891] = 16'b0000000000000000;
	sram_mem[103892] = 16'b0000000000000000;
	sram_mem[103893] = 16'b0000000000000000;
	sram_mem[103894] = 16'b0000000000000000;
	sram_mem[103895] = 16'b0000000000000000;
	sram_mem[103896] = 16'b0000000000000000;
	sram_mem[103897] = 16'b0000000000000000;
	sram_mem[103898] = 16'b0000000000000000;
	sram_mem[103899] = 16'b0000000000000000;
	sram_mem[103900] = 16'b0000000000000000;
	sram_mem[103901] = 16'b0000000000000000;
	sram_mem[103902] = 16'b0000000000000000;
	sram_mem[103903] = 16'b0000000000000000;
	sram_mem[103904] = 16'b0000000000000000;
	sram_mem[103905] = 16'b0000000000000000;
	sram_mem[103906] = 16'b0000000000000000;
	sram_mem[103907] = 16'b0000000000000000;
	sram_mem[103908] = 16'b0000000000000000;
	sram_mem[103909] = 16'b0000000000000000;
	sram_mem[103910] = 16'b0000000000000000;
	sram_mem[103911] = 16'b0000000000000000;
	sram_mem[103912] = 16'b0000000000000000;
	sram_mem[103913] = 16'b0000000000000000;
	sram_mem[103914] = 16'b0000000000000000;
	sram_mem[103915] = 16'b0000000000000000;
	sram_mem[103916] = 16'b0000000000000000;
	sram_mem[103917] = 16'b0000000000000000;
	sram_mem[103918] = 16'b0000000000000000;
	sram_mem[103919] = 16'b0000000000000000;
	sram_mem[103920] = 16'b0000000000000000;
	sram_mem[103921] = 16'b0000000000000000;
	sram_mem[103922] = 16'b0000000000000000;
	sram_mem[103923] = 16'b0000000000000000;
	sram_mem[103924] = 16'b0000000000000000;
	sram_mem[103925] = 16'b0000000000000000;
	sram_mem[103926] = 16'b0000000000000000;
	sram_mem[103927] = 16'b0000000000000000;
	sram_mem[103928] = 16'b0000000000000000;
	sram_mem[103929] = 16'b0000000000000000;
	sram_mem[103930] = 16'b0000000000000000;
	sram_mem[103931] = 16'b0000000000000000;
	sram_mem[103932] = 16'b0000000000000000;
	sram_mem[103933] = 16'b0000000000000000;
	sram_mem[103934] = 16'b0000000000000000;
	sram_mem[103935] = 16'b0000000000000000;
	sram_mem[103936] = 16'b0000000000000000;
	sram_mem[103937] = 16'b0000000000000000;
	sram_mem[103938] = 16'b0000000000000000;
	sram_mem[103939] = 16'b0000000000000000;
	sram_mem[103940] = 16'b0000000000000000;
	sram_mem[103941] = 16'b0000000000000000;
	sram_mem[103942] = 16'b0000000000000000;
	sram_mem[103943] = 16'b0000000000000000;
	sram_mem[103944] = 16'b0000000000000000;
	sram_mem[103945] = 16'b0000000000000000;
	sram_mem[103946] = 16'b0000000000000000;
	sram_mem[103947] = 16'b0000000000000000;
	sram_mem[103948] = 16'b0000000000000000;
	sram_mem[103949] = 16'b0000000000000000;
	sram_mem[103950] = 16'b0000000000000000;
	sram_mem[103951] = 16'b0000000000000000;
	sram_mem[103952] = 16'b0000000000000000;
	sram_mem[103953] = 16'b0000000000000000;
	sram_mem[103954] = 16'b0000000000000000;
	sram_mem[103955] = 16'b0000000000000000;
	sram_mem[103956] = 16'b0000000000000000;
	sram_mem[103957] = 16'b0000000000000000;
	sram_mem[103958] = 16'b0000000000000000;
	sram_mem[103959] = 16'b0000000000000000;
	sram_mem[103960] = 16'b0000000000000000;
	sram_mem[103961] = 16'b0000000000000000;
	sram_mem[103962] = 16'b0000000000000000;
	sram_mem[103963] = 16'b0000000000000000;
	sram_mem[103964] = 16'b0000000000000000;
	sram_mem[103965] = 16'b0000000000000000;
	sram_mem[103966] = 16'b0000000000000000;
	sram_mem[103967] = 16'b0000000000000000;
	sram_mem[103968] = 16'b0000000000000000;
	sram_mem[103969] = 16'b0000000000000000;
	sram_mem[103970] = 16'b0000000000000000;
	sram_mem[103971] = 16'b0000000000000000;
	sram_mem[103972] = 16'b0000000000000000;
	sram_mem[103973] = 16'b0000000000000000;
	sram_mem[103974] = 16'b0000000000000000;
	sram_mem[103975] = 16'b0000000000000000;
	sram_mem[103976] = 16'b0000000000000000;
	sram_mem[103977] = 16'b0000000000000000;
	sram_mem[103978] = 16'b0000000000000000;
	sram_mem[103979] = 16'b0000000000000000;
	sram_mem[103980] = 16'b0000000000000000;
	sram_mem[103981] = 16'b0000000000000000;
	sram_mem[103982] = 16'b0000000000000000;
	sram_mem[103983] = 16'b0000000000000000;
	sram_mem[103984] = 16'b0000000000000000;
	sram_mem[103985] = 16'b0000000000000000;
	sram_mem[103986] = 16'b0000000000000000;
	sram_mem[103987] = 16'b0000000000000000;
	sram_mem[103988] = 16'b0000000000000000;
	sram_mem[103989] = 16'b0000000000000000;
	sram_mem[103990] = 16'b0000000000000000;
	sram_mem[103991] = 16'b0000000000000000;
	sram_mem[103992] = 16'b0000000000000000;
	sram_mem[103993] = 16'b0000000000000000;
	sram_mem[103994] = 16'b0000000000000000;
	sram_mem[103995] = 16'b0000000000000000;
	sram_mem[103996] = 16'b0000000000000000;
	sram_mem[103997] = 16'b0000000000000000;
	sram_mem[103998] = 16'b0000000000000000;
	sram_mem[103999] = 16'b0000000000000000;
	sram_mem[104000] = 16'b0000000000000000;
	sram_mem[104001] = 16'b0000000000000000;
	sram_mem[104002] = 16'b0000000000000000;
	sram_mem[104003] = 16'b0000000000000000;
	sram_mem[104004] = 16'b0000000000000000;
	sram_mem[104005] = 16'b0000000000000000;
	sram_mem[104006] = 16'b0000000000000000;
	sram_mem[104007] = 16'b0000000000000000;
	sram_mem[104008] = 16'b0000000000000000;
	sram_mem[104009] = 16'b0000000000000000;
	sram_mem[104010] = 16'b0000000000000000;
	sram_mem[104011] = 16'b0000000000000000;
	sram_mem[104012] = 16'b0000000000000000;
	sram_mem[104013] = 16'b0000000000000000;
	sram_mem[104014] = 16'b0000000000000000;
	sram_mem[104015] = 16'b0000000000000000;
	sram_mem[104016] = 16'b0000000000000000;
	sram_mem[104017] = 16'b0000000000000000;
	sram_mem[104018] = 16'b0000000000000000;
	sram_mem[104019] = 16'b0000000000000000;
	sram_mem[104020] = 16'b0000000000000000;
	sram_mem[104021] = 16'b0000000000000000;
	sram_mem[104022] = 16'b0000000000000000;
	sram_mem[104023] = 16'b0000000000000000;
	sram_mem[104024] = 16'b0000000000000000;
	sram_mem[104025] = 16'b0000000000000000;
	sram_mem[104026] = 16'b0000000000000000;
	sram_mem[104027] = 16'b0000000000000000;
	sram_mem[104028] = 16'b0000000000000000;
	sram_mem[104029] = 16'b0000000000000000;
	sram_mem[104030] = 16'b0000000000000000;
	sram_mem[104031] = 16'b0000000000000000;
	sram_mem[104032] = 16'b0000000000000000;
	sram_mem[104033] = 16'b0000000000000000;
	sram_mem[104034] = 16'b0000000000000000;
	sram_mem[104035] = 16'b0000000000000000;
	sram_mem[104036] = 16'b0000000000000000;
	sram_mem[104037] = 16'b0000000000000000;
	sram_mem[104038] = 16'b0000000000000000;
	sram_mem[104039] = 16'b0000000000000000;
	sram_mem[104040] = 16'b0000000000000000;
	sram_mem[104041] = 16'b0000000000000000;
	sram_mem[104042] = 16'b0000000000000000;
	sram_mem[104043] = 16'b0000000000000000;
	sram_mem[104044] = 16'b0000000000000000;
	sram_mem[104045] = 16'b0000000000000000;
	sram_mem[104046] = 16'b0000000000000000;
	sram_mem[104047] = 16'b0000000000000000;
	sram_mem[104048] = 16'b0000000000000000;
	sram_mem[104049] = 16'b0000000000000000;
	sram_mem[104050] = 16'b0000000000000000;
	sram_mem[104051] = 16'b0000000000000000;
	sram_mem[104052] = 16'b0000000000000000;
	sram_mem[104053] = 16'b0000000000000000;
	sram_mem[104054] = 16'b0000000000000000;
	sram_mem[104055] = 16'b0000000000000000;
	sram_mem[104056] = 16'b0000000000000000;
	sram_mem[104057] = 16'b0000000000000000;
	sram_mem[104058] = 16'b0000000000000000;
	sram_mem[104059] = 16'b0000000000000000;
	sram_mem[104060] = 16'b0000000000000000;
	sram_mem[104061] = 16'b0000000000000000;
	sram_mem[104062] = 16'b0000000000000000;
	sram_mem[104063] = 16'b0000000000000000;
	sram_mem[104064] = 16'b0000000000000000;
	sram_mem[104065] = 16'b0000000000000000;
	sram_mem[104066] = 16'b0000000000000000;
	sram_mem[104067] = 16'b0000000000000000;
	sram_mem[104068] = 16'b0000000000000000;
	sram_mem[104069] = 16'b0000000000000000;
	sram_mem[104070] = 16'b0000000000000000;
	sram_mem[104071] = 16'b0000000000000000;
	sram_mem[104072] = 16'b0000000000000000;
	sram_mem[104073] = 16'b0000000000000000;
	sram_mem[104074] = 16'b0000000000000000;
	sram_mem[104075] = 16'b0000000000000000;
	sram_mem[104076] = 16'b0000000000000000;
	sram_mem[104077] = 16'b0000000000000000;
	sram_mem[104078] = 16'b0000000000000000;
	sram_mem[104079] = 16'b0000000000000000;
	sram_mem[104080] = 16'b0000000000000000;
	sram_mem[104081] = 16'b0000000000000000;
	sram_mem[104082] = 16'b0000000000000000;
	sram_mem[104083] = 16'b0000000000000000;
	sram_mem[104084] = 16'b0000000000000000;
	sram_mem[104085] = 16'b0000000000000000;
	sram_mem[104086] = 16'b0000000000000000;
	sram_mem[104087] = 16'b0000000000000000;
	sram_mem[104088] = 16'b0000000000000000;
	sram_mem[104089] = 16'b0000000000000000;
	sram_mem[104090] = 16'b0000000000000000;
	sram_mem[104091] = 16'b0000000000000000;
	sram_mem[104092] = 16'b0000000000000000;
	sram_mem[104093] = 16'b0000000000000000;
	sram_mem[104094] = 16'b0000000000000000;
	sram_mem[104095] = 16'b0000000000000000;
	sram_mem[104096] = 16'b0000000000000000;
	sram_mem[104097] = 16'b0000000000000000;
	sram_mem[104098] = 16'b0000000000000000;
	sram_mem[104099] = 16'b0000000000000000;
	sram_mem[104100] = 16'b0000000000000000;
	sram_mem[104101] = 16'b0000000000000000;
	sram_mem[104102] = 16'b0000000000000000;
	sram_mem[104103] = 16'b0000000000000000;
	sram_mem[104104] = 16'b0000000000000000;
	sram_mem[104105] = 16'b0000000000000000;
	sram_mem[104106] = 16'b0000000000000000;
	sram_mem[104107] = 16'b0000000000000000;
	sram_mem[104108] = 16'b0000000000000000;
	sram_mem[104109] = 16'b0000000000000000;
	sram_mem[104110] = 16'b0000000000000000;
	sram_mem[104111] = 16'b0000000000000000;
	sram_mem[104112] = 16'b0000000000000000;
	sram_mem[104113] = 16'b0000000000000000;
	sram_mem[104114] = 16'b0000000000000000;
	sram_mem[104115] = 16'b0000000000000000;
	sram_mem[104116] = 16'b0000000000000000;
	sram_mem[104117] = 16'b0000000000000000;
	sram_mem[104118] = 16'b0000000000000000;
	sram_mem[104119] = 16'b0000000000000000;
	sram_mem[104120] = 16'b0000000000000000;
	sram_mem[104121] = 16'b0000000000000000;
	sram_mem[104122] = 16'b0000000000000000;
	sram_mem[104123] = 16'b0000000000000000;
	sram_mem[104124] = 16'b0000000000000000;
	sram_mem[104125] = 16'b0000000000000000;
	sram_mem[104126] = 16'b0000000000000000;
	sram_mem[104127] = 16'b0000000000000000;
	sram_mem[104128] = 16'b0000000000000000;
	sram_mem[104129] = 16'b0000000000000000;
	sram_mem[104130] = 16'b0000000000000000;
	sram_mem[104131] = 16'b0000000000000000;
	sram_mem[104132] = 16'b0000000000000000;
	sram_mem[104133] = 16'b0000000000000000;
	sram_mem[104134] = 16'b0000000000000000;
	sram_mem[104135] = 16'b0000000000000000;
	sram_mem[104136] = 16'b0000000000000000;
	sram_mem[104137] = 16'b0000000000000000;
	sram_mem[104138] = 16'b0000000000000000;
	sram_mem[104139] = 16'b0000000000000000;
	sram_mem[104140] = 16'b0000000000000000;
	sram_mem[104141] = 16'b0000000000000000;
	sram_mem[104142] = 16'b0000000000000000;
	sram_mem[104143] = 16'b0000000000000000;
	sram_mem[104144] = 16'b0000000000000000;
	sram_mem[104145] = 16'b0000000000000000;
	sram_mem[104146] = 16'b0000000000000000;
	sram_mem[104147] = 16'b0000000000000000;
	sram_mem[104148] = 16'b0000000000000000;
	sram_mem[104149] = 16'b0000000000000000;
	sram_mem[104150] = 16'b0000000000000000;
	sram_mem[104151] = 16'b0000000000000000;
	sram_mem[104152] = 16'b0000000000000000;
	sram_mem[104153] = 16'b0000000000000000;
	sram_mem[104154] = 16'b0000000000000000;
	sram_mem[104155] = 16'b0000000000000000;
	sram_mem[104156] = 16'b0000000000000000;
	sram_mem[104157] = 16'b0000000000000000;
	sram_mem[104158] = 16'b0000000000000000;
	sram_mem[104159] = 16'b0000000000000000;
	sram_mem[104160] = 16'b0000000000000000;
	sram_mem[104161] = 16'b0000000000000000;
	sram_mem[104162] = 16'b0000000000000000;
	sram_mem[104163] = 16'b0000000000000000;
	sram_mem[104164] = 16'b0000000000000000;
	sram_mem[104165] = 16'b0000000000000000;
	sram_mem[104166] = 16'b0000000000000000;
	sram_mem[104167] = 16'b0000000000000000;
	sram_mem[104168] = 16'b0000000000000000;
	sram_mem[104169] = 16'b0000000000000000;
	sram_mem[104170] = 16'b0000000000000000;
	sram_mem[104171] = 16'b0000000000000000;
	sram_mem[104172] = 16'b0000000000000000;
	sram_mem[104173] = 16'b0000000000000000;
	sram_mem[104174] = 16'b0000000000000000;
	sram_mem[104175] = 16'b0000000000000000;
	sram_mem[104176] = 16'b0000000000000000;
	sram_mem[104177] = 16'b0000000000000000;
	sram_mem[104178] = 16'b0000000000000000;
	sram_mem[104179] = 16'b0000000000000000;
	sram_mem[104180] = 16'b0000000000000000;
	sram_mem[104181] = 16'b0000000000000000;
	sram_mem[104182] = 16'b0000000000000000;
	sram_mem[104183] = 16'b0000000000000000;
	sram_mem[104184] = 16'b0000000000000000;
	sram_mem[104185] = 16'b0000000000000000;
	sram_mem[104186] = 16'b0000000000000000;
	sram_mem[104187] = 16'b0000000000000000;
	sram_mem[104188] = 16'b0000000000000000;
	sram_mem[104189] = 16'b0000000000000000;
	sram_mem[104190] = 16'b0000000000000000;
	sram_mem[104191] = 16'b0000000000000000;
	sram_mem[104192] = 16'b0000000000000000;
	sram_mem[104193] = 16'b0000000000000000;
	sram_mem[104194] = 16'b0000000000000000;
	sram_mem[104195] = 16'b0000000000000000;
	sram_mem[104196] = 16'b0000000000000000;
	sram_mem[104197] = 16'b0000000000000000;
	sram_mem[104198] = 16'b0000000000000000;
	sram_mem[104199] = 16'b0000000000000000;
	sram_mem[104200] = 16'b0000000000000000;
	sram_mem[104201] = 16'b0000000000000000;
	sram_mem[104202] = 16'b0000000000000000;
	sram_mem[104203] = 16'b0000000000000000;
	sram_mem[104204] = 16'b0000000000000000;
	sram_mem[104205] = 16'b0000000000000000;
	sram_mem[104206] = 16'b0000000000000000;
	sram_mem[104207] = 16'b0000000000000000;
	sram_mem[104208] = 16'b0000000000000000;
	sram_mem[104209] = 16'b0000000000000000;
	sram_mem[104210] = 16'b0000000000000000;
	sram_mem[104211] = 16'b0000000000000000;
	sram_mem[104212] = 16'b0000000000000000;
	sram_mem[104213] = 16'b0000000000000000;
	sram_mem[104214] = 16'b0000000000000000;
	sram_mem[104215] = 16'b0000000000000000;
	sram_mem[104216] = 16'b0000000000000000;
	sram_mem[104217] = 16'b0000000000000000;
	sram_mem[104218] = 16'b0000000000000000;
	sram_mem[104219] = 16'b0000000000000000;
	sram_mem[104220] = 16'b0000000000000000;
	sram_mem[104221] = 16'b0000000000000000;
	sram_mem[104222] = 16'b0000000000000000;
	sram_mem[104223] = 16'b0000000000000000;
	sram_mem[104224] = 16'b0000000000000000;
	sram_mem[104225] = 16'b0000000000000000;
	sram_mem[104226] = 16'b0000000000000000;
	sram_mem[104227] = 16'b0000000000000000;
	sram_mem[104228] = 16'b0000000000000000;
	sram_mem[104229] = 16'b0000000000000000;
	sram_mem[104230] = 16'b0000000000000000;
	sram_mem[104231] = 16'b0000000000000000;
	sram_mem[104232] = 16'b0000000000000000;
	sram_mem[104233] = 16'b0000000000000000;
	sram_mem[104234] = 16'b0000000000000000;
	sram_mem[104235] = 16'b0000000000000000;
	sram_mem[104236] = 16'b0000000000000000;
	sram_mem[104237] = 16'b0000000000000000;
	sram_mem[104238] = 16'b0000000000000000;
	sram_mem[104239] = 16'b0000000000000000;
	sram_mem[104240] = 16'b0000000000000000;
	sram_mem[104241] = 16'b0000000000000000;
	sram_mem[104242] = 16'b0000000000000000;
	sram_mem[104243] = 16'b0000000000000000;
	sram_mem[104244] = 16'b0000000000000000;
	sram_mem[104245] = 16'b0000000000000000;
	sram_mem[104246] = 16'b0000000000000000;
	sram_mem[104247] = 16'b0000000000000000;
	sram_mem[104248] = 16'b0000000000000000;
	sram_mem[104249] = 16'b0000000000000000;
	sram_mem[104250] = 16'b0000000000000000;
	sram_mem[104251] = 16'b0000000000000000;
	sram_mem[104252] = 16'b0000000000000000;
	sram_mem[104253] = 16'b0000000000000000;
	sram_mem[104254] = 16'b0000000000000000;
	sram_mem[104255] = 16'b0000000000000000;
	sram_mem[104256] = 16'b0000000000000000;
	sram_mem[104257] = 16'b0000000000000000;
	sram_mem[104258] = 16'b0000000000000000;
	sram_mem[104259] = 16'b0000000000000000;
	sram_mem[104260] = 16'b0000000000000000;
	sram_mem[104261] = 16'b0000000000000000;
	sram_mem[104262] = 16'b0000000000000000;
	sram_mem[104263] = 16'b0000000000000000;
	sram_mem[104264] = 16'b0000000000000000;
	sram_mem[104265] = 16'b0000000000000000;
	sram_mem[104266] = 16'b0000000000000000;
	sram_mem[104267] = 16'b0000000000000000;
	sram_mem[104268] = 16'b0000000000000000;
	sram_mem[104269] = 16'b0000000000000000;
	sram_mem[104270] = 16'b0000000000000000;
	sram_mem[104271] = 16'b0000000000000000;
	sram_mem[104272] = 16'b0000000000000000;
	sram_mem[104273] = 16'b0000000000000000;
	sram_mem[104274] = 16'b0000000000000000;
	sram_mem[104275] = 16'b0000000000000000;
	sram_mem[104276] = 16'b0000000000000000;
	sram_mem[104277] = 16'b0000000000000000;
	sram_mem[104278] = 16'b0000000000000000;
	sram_mem[104279] = 16'b0000000000000000;
	sram_mem[104280] = 16'b0000000000000000;
	sram_mem[104281] = 16'b0000000000000000;
	sram_mem[104282] = 16'b0000000000000000;
	sram_mem[104283] = 16'b0000000000000000;
	sram_mem[104284] = 16'b0000000000000000;
	sram_mem[104285] = 16'b0000000000000000;
	sram_mem[104286] = 16'b0000000000000000;
	sram_mem[104287] = 16'b0000000000000000;
	sram_mem[104288] = 16'b0000000000000000;
	sram_mem[104289] = 16'b0000000000000000;
	sram_mem[104290] = 16'b0000000000000000;
	sram_mem[104291] = 16'b0000000000000000;
	sram_mem[104292] = 16'b0000000000000000;
	sram_mem[104293] = 16'b0000000000000000;
	sram_mem[104294] = 16'b0000000000000000;
	sram_mem[104295] = 16'b0000000000000000;
	sram_mem[104296] = 16'b0000000000000000;
	sram_mem[104297] = 16'b0000000000000000;
	sram_mem[104298] = 16'b0000000000000000;
	sram_mem[104299] = 16'b0000000000000000;
	sram_mem[104300] = 16'b0000000000000000;
	sram_mem[104301] = 16'b0000000000000000;
	sram_mem[104302] = 16'b0000000000000000;
	sram_mem[104303] = 16'b0000000000000000;
	sram_mem[104304] = 16'b0000000000000000;
	sram_mem[104305] = 16'b0000000000000000;
	sram_mem[104306] = 16'b0000000000000000;
	sram_mem[104307] = 16'b0000000000000000;
	sram_mem[104308] = 16'b0000000000000000;
	sram_mem[104309] = 16'b0000000000000000;
	sram_mem[104310] = 16'b0000000000000000;
	sram_mem[104311] = 16'b0000000000000000;
	sram_mem[104312] = 16'b0000000000000000;
	sram_mem[104313] = 16'b0000000000000000;
	sram_mem[104314] = 16'b0000000000000000;
	sram_mem[104315] = 16'b0000000000000000;
	sram_mem[104316] = 16'b0000000000000000;
	sram_mem[104317] = 16'b0000000000000000;
	sram_mem[104318] = 16'b0000000000000000;
	sram_mem[104319] = 16'b0000000000000000;
	sram_mem[104320] = 16'b0000000000000000;
	sram_mem[104321] = 16'b0000000000000000;
	sram_mem[104322] = 16'b0000000000000000;
	sram_mem[104323] = 16'b0000000000000000;
	sram_mem[104324] = 16'b0000000000000000;
	sram_mem[104325] = 16'b0000000000000000;
	sram_mem[104326] = 16'b0000000000000000;
	sram_mem[104327] = 16'b0000000000000000;
	sram_mem[104328] = 16'b0000000000000000;
	sram_mem[104329] = 16'b0000000000000000;
	sram_mem[104330] = 16'b0000000000000000;
	sram_mem[104331] = 16'b0000000000000000;
	sram_mem[104332] = 16'b0000000000000000;
	sram_mem[104333] = 16'b0000000000000000;
	sram_mem[104334] = 16'b0000000000000000;
	sram_mem[104335] = 16'b0000000000000000;
	sram_mem[104336] = 16'b0000000000000000;
	sram_mem[104337] = 16'b0000000000000000;
	sram_mem[104338] = 16'b0000000000000000;
	sram_mem[104339] = 16'b0000000000000000;
	sram_mem[104340] = 16'b0000000000000000;
	sram_mem[104341] = 16'b0000000000000000;
	sram_mem[104342] = 16'b0000000000000000;
	sram_mem[104343] = 16'b0000000000000000;
	sram_mem[104344] = 16'b0000000000000000;
	sram_mem[104345] = 16'b0000000000000000;
	sram_mem[104346] = 16'b0000000000000000;
	sram_mem[104347] = 16'b0000000000000000;
	sram_mem[104348] = 16'b0000000000000000;
	sram_mem[104349] = 16'b0000000000000000;
	sram_mem[104350] = 16'b0000000000000000;
	sram_mem[104351] = 16'b0000000000000000;
	sram_mem[104352] = 16'b0000000000000000;
	sram_mem[104353] = 16'b0000000000000000;
	sram_mem[104354] = 16'b0000000000000000;
	sram_mem[104355] = 16'b0000000000000000;
	sram_mem[104356] = 16'b0000000000000000;
	sram_mem[104357] = 16'b0000000000000000;
	sram_mem[104358] = 16'b0000000000000000;
	sram_mem[104359] = 16'b0000000000000000;
	sram_mem[104360] = 16'b0000000000000000;
	sram_mem[104361] = 16'b0000000000000000;
	sram_mem[104362] = 16'b0000000000000000;
	sram_mem[104363] = 16'b0000000000000000;
	sram_mem[104364] = 16'b0000000000000000;
	sram_mem[104365] = 16'b0000000000000000;
	sram_mem[104366] = 16'b0000000000000000;
	sram_mem[104367] = 16'b0000000000000000;
	sram_mem[104368] = 16'b0000000000000000;
	sram_mem[104369] = 16'b0000000000000000;
	sram_mem[104370] = 16'b0000000000000000;
	sram_mem[104371] = 16'b0000000000000000;
	sram_mem[104372] = 16'b0000000000000000;
	sram_mem[104373] = 16'b0000000000000000;
	sram_mem[104374] = 16'b0000000000000000;
	sram_mem[104375] = 16'b0000000000000000;
	sram_mem[104376] = 16'b0000000000000000;
	sram_mem[104377] = 16'b0000000000000000;
	sram_mem[104378] = 16'b0000000000000000;
	sram_mem[104379] = 16'b0000000000000000;
	sram_mem[104380] = 16'b0000000000000000;
	sram_mem[104381] = 16'b0000000000000000;
	sram_mem[104382] = 16'b0000000000000000;
	sram_mem[104383] = 16'b0000000000000000;
	sram_mem[104384] = 16'b0000000000000000;
	sram_mem[104385] = 16'b0000000000000000;
	sram_mem[104386] = 16'b0000000000000000;
	sram_mem[104387] = 16'b0000000000000000;
	sram_mem[104388] = 16'b0000000000000000;
	sram_mem[104389] = 16'b0000000000000000;
	sram_mem[104390] = 16'b0000000000000000;
	sram_mem[104391] = 16'b0000000000000000;
	sram_mem[104392] = 16'b0000000000000000;
	sram_mem[104393] = 16'b0000000000000000;
	sram_mem[104394] = 16'b0000000000000000;
	sram_mem[104395] = 16'b0000000000000000;
	sram_mem[104396] = 16'b0000000000000000;
	sram_mem[104397] = 16'b0000000000000000;
	sram_mem[104398] = 16'b0000000000000000;
	sram_mem[104399] = 16'b0000000000000000;
	sram_mem[104400] = 16'b0000000000000000;
	sram_mem[104401] = 16'b0000000000000000;
	sram_mem[104402] = 16'b0000000000000000;
	sram_mem[104403] = 16'b0000000000000000;
	sram_mem[104404] = 16'b0000000000000000;
	sram_mem[104405] = 16'b0000000000000000;
	sram_mem[104406] = 16'b0000000000000000;
	sram_mem[104407] = 16'b0000000000000000;
	sram_mem[104408] = 16'b0000000000000000;
	sram_mem[104409] = 16'b0000000000000000;
	sram_mem[104410] = 16'b0000000000000000;
	sram_mem[104411] = 16'b0000000000000000;
	sram_mem[104412] = 16'b0000000000000000;
	sram_mem[104413] = 16'b0000000000000000;
	sram_mem[104414] = 16'b0000000000000000;
	sram_mem[104415] = 16'b0000000000000000;
	sram_mem[104416] = 16'b0000000000000000;
	sram_mem[104417] = 16'b0000000000000000;
	sram_mem[104418] = 16'b0000000000000000;
	sram_mem[104419] = 16'b0000000000000000;
	sram_mem[104420] = 16'b0000000000000000;
	sram_mem[104421] = 16'b0000000000000000;
	sram_mem[104422] = 16'b0000000000000000;
	sram_mem[104423] = 16'b0000000000000000;
	sram_mem[104424] = 16'b0000000000000000;
	sram_mem[104425] = 16'b0000000000000000;
	sram_mem[104426] = 16'b0000000000000000;
	sram_mem[104427] = 16'b0000000000000000;
	sram_mem[104428] = 16'b0000000000000000;
	sram_mem[104429] = 16'b0000000000000000;
	sram_mem[104430] = 16'b0000000000000000;
	sram_mem[104431] = 16'b0000000000000000;
	sram_mem[104432] = 16'b0000000000000000;
	sram_mem[104433] = 16'b0000000000000000;
	sram_mem[104434] = 16'b0000000000000000;
	sram_mem[104435] = 16'b0000000000000000;
	sram_mem[104436] = 16'b0000000000000000;
	sram_mem[104437] = 16'b0000000000000000;
	sram_mem[104438] = 16'b0000000000000000;
	sram_mem[104439] = 16'b0000000000000000;
	sram_mem[104440] = 16'b0000000000000000;
	sram_mem[104441] = 16'b0000000000000000;
	sram_mem[104442] = 16'b0000000000000000;
	sram_mem[104443] = 16'b0000000000000000;
	sram_mem[104444] = 16'b0000000000000000;
	sram_mem[104445] = 16'b0000000000000000;
	sram_mem[104446] = 16'b0000000000000000;
	sram_mem[104447] = 16'b0000000000000000;
	sram_mem[104448] = 16'b0000000000000000;
	sram_mem[104449] = 16'b0000000000000000;
	sram_mem[104450] = 16'b0000000000000000;
	sram_mem[104451] = 16'b0000000000000000;
	sram_mem[104452] = 16'b0000000000000000;
	sram_mem[104453] = 16'b0000000000000000;
	sram_mem[104454] = 16'b0000000000000000;
	sram_mem[104455] = 16'b0000000000000000;
	sram_mem[104456] = 16'b0000000000000000;
	sram_mem[104457] = 16'b0000000000000000;
	sram_mem[104458] = 16'b0000000000000000;
	sram_mem[104459] = 16'b0000000000000000;
	sram_mem[104460] = 16'b0000000000000000;
	sram_mem[104461] = 16'b0000000000000000;
	sram_mem[104462] = 16'b0000000000000000;
	sram_mem[104463] = 16'b0000000000000000;
	sram_mem[104464] = 16'b0000000000000000;
	sram_mem[104465] = 16'b0000000000000000;
	sram_mem[104466] = 16'b0000000000000000;
	sram_mem[104467] = 16'b0000000000000000;
	sram_mem[104468] = 16'b0000000000000000;
	sram_mem[104469] = 16'b0000000000000000;
	sram_mem[104470] = 16'b0000000000000000;
	sram_mem[104471] = 16'b0000000000000000;
	sram_mem[104472] = 16'b0000000000000000;
	sram_mem[104473] = 16'b0000000000000000;
	sram_mem[104474] = 16'b0000000000000000;
	sram_mem[104475] = 16'b0000000000000000;
	sram_mem[104476] = 16'b0000000000000000;
	sram_mem[104477] = 16'b0000000000000000;
	sram_mem[104478] = 16'b0000000000000000;
	sram_mem[104479] = 16'b0000000000000000;
	sram_mem[104480] = 16'b0000000000000000;
	sram_mem[104481] = 16'b0000000000000000;
	sram_mem[104482] = 16'b0000000000000000;
	sram_mem[104483] = 16'b0000000000000000;
	sram_mem[104484] = 16'b0000000000000000;
	sram_mem[104485] = 16'b0000000000000000;
	sram_mem[104486] = 16'b0000000000000000;
	sram_mem[104487] = 16'b0000000000000000;
	sram_mem[104488] = 16'b0000000000000000;
	sram_mem[104489] = 16'b0000000000000000;
	sram_mem[104490] = 16'b0000000000000000;
	sram_mem[104491] = 16'b0000000000000000;
	sram_mem[104492] = 16'b0000000000000000;
	sram_mem[104493] = 16'b0000000000000000;
	sram_mem[104494] = 16'b0000000000000000;
	sram_mem[104495] = 16'b0000000000000000;
	sram_mem[104496] = 16'b0000000000000000;
	sram_mem[104497] = 16'b0000000000000000;
	sram_mem[104498] = 16'b0000000000000000;
	sram_mem[104499] = 16'b0000000000000000;
	sram_mem[104500] = 16'b0000000000000000;
	sram_mem[104501] = 16'b0000000000000000;
	sram_mem[104502] = 16'b0000000000000000;
	sram_mem[104503] = 16'b0000000000000000;
	sram_mem[104504] = 16'b0000000000000000;
	sram_mem[104505] = 16'b0000000000000000;
	sram_mem[104506] = 16'b0000000000000000;
	sram_mem[104507] = 16'b0000000000000000;
	sram_mem[104508] = 16'b0000000000000000;
	sram_mem[104509] = 16'b0000000000000000;
	sram_mem[104510] = 16'b0000000000000000;
	sram_mem[104511] = 16'b0000000000000000;
	sram_mem[104512] = 16'b0000000000000000;
	sram_mem[104513] = 16'b0000000000000000;
	sram_mem[104514] = 16'b0000000000000000;
	sram_mem[104515] = 16'b0000000000000000;
	sram_mem[104516] = 16'b0000000000000000;
	sram_mem[104517] = 16'b0000000000000000;
	sram_mem[104518] = 16'b0000000000000000;
	sram_mem[104519] = 16'b0000000000000000;
	sram_mem[104520] = 16'b0000000000000000;
	sram_mem[104521] = 16'b0000000000000000;
	sram_mem[104522] = 16'b0000000000000000;
	sram_mem[104523] = 16'b0000000000000000;
	sram_mem[104524] = 16'b0000000000000000;
	sram_mem[104525] = 16'b0000000000000000;
	sram_mem[104526] = 16'b0000000000000000;
	sram_mem[104527] = 16'b0000000000000000;
	sram_mem[104528] = 16'b0000000000000000;
	sram_mem[104529] = 16'b0000000000000000;
	sram_mem[104530] = 16'b0000000000000000;
	sram_mem[104531] = 16'b0000000000000000;
	sram_mem[104532] = 16'b0000000000000000;
	sram_mem[104533] = 16'b0000000000000000;
	sram_mem[104534] = 16'b0000000000000000;
	sram_mem[104535] = 16'b0000000000000000;
	sram_mem[104536] = 16'b0000000000000000;
	sram_mem[104537] = 16'b0000000000000000;
	sram_mem[104538] = 16'b0000000000000000;
	sram_mem[104539] = 16'b0000000000000000;
	sram_mem[104540] = 16'b0000000000000000;
	sram_mem[104541] = 16'b0000000000000000;
	sram_mem[104542] = 16'b0000000000000000;
	sram_mem[104543] = 16'b0000000000000000;
	sram_mem[104544] = 16'b0000000000000000;
	sram_mem[104545] = 16'b0000000000000000;
	sram_mem[104546] = 16'b0000000000000000;
	sram_mem[104547] = 16'b0000000000000000;
	sram_mem[104548] = 16'b0000000000000000;
	sram_mem[104549] = 16'b0000000000000000;
	sram_mem[104550] = 16'b0000000000000000;
	sram_mem[104551] = 16'b0000000000000000;
	sram_mem[104552] = 16'b0000000000000000;
	sram_mem[104553] = 16'b0000000000000000;
	sram_mem[104554] = 16'b0000000000000000;
	sram_mem[104555] = 16'b0000000000000000;
	sram_mem[104556] = 16'b0000000000000000;
	sram_mem[104557] = 16'b0000000000000000;
	sram_mem[104558] = 16'b0000000000000000;
	sram_mem[104559] = 16'b0000000000000000;
	sram_mem[104560] = 16'b0000000000000000;
	sram_mem[104561] = 16'b0000000000000000;
	sram_mem[104562] = 16'b0000000000000000;
	sram_mem[104563] = 16'b0000000000000000;
	sram_mem[104564] = 16'b0000000000000000;
	sram_mem[104565] = 16'b0000000000000000;
	sram_mem[104566] = 16'b0000000000000000;
	sram_mem[104567] = 16'b0000000000000000;
	sram_mem[104568] = 16'b0000000000000000;
	sram_mem[104569] = 16'b0000000000000000;
	sram_mem[104570] = 16'b0000000000000000;
	sram_mem[104571] = 16'b0000000000000000;
	sram_mem[104572] = 16'b0000000000000000;
	sram_mem[104573] = 16'b0000000000000000;
	sram_mem[104574] = 16'b0000000000000000;
	sram_mem[104575] = 16'b0000000000000000;
	sram_mem[104576] = 16'b0000000000000000;
	sram_mem[104577] = 16'b0000000000000000;
	sram_mem[104578] = 16'b0000000000000000;
	sram_mem[104579] = 16'b0000000000000000;
	sram_mem[104580] = 16'b0000000000000000;
	sram_mem[104581] = 16'b0000000000000000;
	sram_mem[104582] = 16'b0000000000000000;
	sram_mem[104583] = 16'b0000000000000000;
	sram_mem[104584] = 16'b0000000000000000;
	sram_mem[104585] = 16'b0000000000000000;
	sram_mem[104586] = 16'b0000000000000000;
	sram_mem[104587] = 16'b0000000000000000;
	sram_mem[104588] = 16'b0000000000000000;
	sram_mem[104589] = 16'b0000000000000000;
	sram_mem[104590] = 16'b0000000000000000;
	sram_mem[104591] = 16'b0000000000000000;
	sram_mem[104592] = 16'b0000000000000000;
	sram_mem[104593] = 16'b0000000000000000;
	sram_mem[104594] = 16'b0000000000000000;
	sram_mem[104595] = 16'b0000000000000000;
	sram_mem[104596] = 16'b0000000000000000;
	sram_mem[104597] = 16'b0000000000000000;
	sram_mem[104598] = 16'b0000000000000000;
	sram_mem[104599] = 16'b0000000000000000;
	sram_mem[104600] = 16'b0000000000000000;
	sram_mem[104601] = 16'b0000000000000000;
	sram_mem[104602] = 16'b0000000000000000;
	sram_mem[104603] = 16'b0000000000000000;
	sram_mem[104604] = 16'b0000000000000000;
	sram_mem[104605] = 16'b0000000000000000;
	sram_mem[104606] = 16'b0000000000000000;
	sram_mem[104607] = 16'b0000000000000000;
	sram_mem[104608] = 16'b0000000000000000;
	sram_mem[104609] = 16'b0000000000000000;
	sram_mem[104610] = 16'b0000000000000000;
	sram_mem[104611] = 16'b0000000000000000;
	sram_mem[104612] = 16'b0000000000000000;
	sram_mem[104613] = 16'b0000000000000000;
	sram_mem[104614] = 16'b0000000000000000;
	sram_mem[104615] = 16'b0000000000000000;
	sram_mem[104616] = 16'b0000000000000000;
	sram_mem[104617] = 16'b0000000000000000;
	sram_mem[104618] = 16'b0000000000000000;
	sram_mem[104619] = 16'b0000000000000000;
	sram_mem[104620] = 16'b0000000000000000;
	sram_mem[104621] = 16'b0000000000000000;
	sram_mem[104622] = 16'b0000000000000000;
	sram_mem[104623] = 16'b0000000000000000;
	sram_mem[104624] = 16'b0000000000000000;
	sram_mem[104625] = 16'b0000000000000000;
	sram_mem[104626] = 16'b0000000000000000;
	sram_mem[104627] = 16'b0000000000000000;
	sram_mem[104628] = 16'b0000000000000000;
	sram_mem[104629] = 16'b0000000000000000;
	sram_mem[104630] = 16'b0000000000000000;
	sram_mem[104631] = 16'b0000000000000000;
	sram_mem[104632] = 16'b0000000000000000;
	sram_mem[104633] = 16'b0000000000000000;
	sram_mem[104634] = 16'b0000000000000000;
	sram_mem[104635] = 16'b0000000000000000;
	sram_mem[104636] = 16'b0000000000000000;
	sram_mem[104637] = 16'b0000000000000000;
	sram_mem[104638] = 16'b0000000000000000;
	sram_mem[104639] = 16'b0000000000000000;
	sram_mem[104640] = 16'b0000000000000000;
	sram_mem[104641] = 16'b0000000000000000;
	sram_mem[104642] = 16'b0000000000000000;
	sram_mem[104643] = 16'b0000000000000000;
	sram_mem[104644] = 16'b0000000000000000;
	sram_mem[104645] = 16'b0000000000000000;
	sram_mem[104646] = 16'b0000000000000000;
	sram_mem[104647] = 16'b0000000000000000;
	sram_mem[104648] = 16'b0000000000000000;
	sram_mem[104649] = 16'b0000000000000000;
	sram_mem[104650] = 16'b0000000000000000;
	sram_mem[104651] = 16'b0000000000000000;
	sram_mem[104652] = 16'b0000000000000000;
	sram_mem[104653] = 16'b0000000000000000;
	sram_mem[104654] = 16'b0000000000000000;
	sram_mem[104655] = 16'b0000000000000000;
	sram_mem[104656] = 16'b0000000000000000;
	sram_mem[104657] = 16'b0000000000000000;
	sram_mem[104658] = 16'b0000000000000000;
	sram_mem[104659] = 16'b0000000000000000;
	sram_mem[104660] = 16'b0000000000000000;
	sram_mem[104661] = 16'b0000000000000000;
	sram_mem[104662] = 16'b0000000000000000;
	sram_mem[104663] = 16'b0000000000000000;
	sram_mem[104664] = 16'b0000000000000000;
	sram_mem[104665] = 16'b0000000000000000;
	sram_mem[104666] = 16'b0000000000000000;
	sram_mem[104667] = 16'b0000000000000000;
	sram_mem[104668] = 16'b0000000000000000;
	sram_mem[104669] = 16'b0000000000000000;
	sram_mem[104670] = 16'b0000000000000000;
	sram_mem[104671] = 16'b0000000000000000;
	sram_mem[104672] = 16'b0000000000000000;
	sram_mem[104673] = 16'b0000000000000000;
	sram_mem[104674] = 16'b0000000000000000;
	sram_mem[104675] = 16'b0000000000000000;
	sram_mem[104676] = 16'b0000000000000000;
	sram_mem[104677] = 16'b0000000000000000;
	sram_mem[104678] = 16'b0000000000000000;
	sram_mem[104679] = 16'b0000000000000000;
	sram_mem[104680] = 16'b0000000000000000;
	sram_mem[104681] = 16'b0000000000000000;
	sram_mem[104682] = 16'b0000000000000000;
	sram_mem[104683] = 16'b0000000000000000;
	sram_mem[104684] = 16'b0000000000000000;
	sram_mem[104685] = 16'b0000000000000000;
	sram_mem[104686] = 16'b0000000000000000;
	sram_mem[104687] = 16'b0000000000000000;
	sram_mem[104688] = 16'b0000000000000000;
	sram_mem[104689] = 16'b0000000000000000;
	sram_mem[104690] = 16'b0000000000000000;
	sram_mem[104691] = 16'b0000000000000000;
	sram_mem[104692] = 16'b0000000000000000;
	sram_mem[104693] = 16'b0000000000000000;
	sram_mem[104694] = 16'b0000000000000000;
	sram_mem[104695] = 16'b0000000000000000;
	sram_mem[104696] = 16'b0000000000000000;
	sram_mem[104697] = 16'b0000000000000000;
	sram_mem[104698] = 16'b0000000000000000;
	sram_mem[104699] = 16'b0000000000000000;
	sram_mem[104700] = 16'b0000000000000000;
	sram_mem[104701] = 16'b0000000000000000;
	sram_mem[104702] = 16'b0000000000000000;
	sram_mem[104703] = 16'b0000000000000000;
	sram_mem[104704] = 16'b0000000000000000;
	sram_mem[104705] = 16'b0000000000000000;
	sram_mem[104706] = 16'b0000000000000000;
	sram_mem[104707] = 16'b0000000000000000;
	sram_mem[104708] = 16'b0000000000000000;
	sram_mem[104709] = 16'b0000000000000000;
	sram_mem[104710] = 16'b0000000000000000;
	sram_mem[104711] = 16'b0000000000000000;
	sram_mem[104712] = 16'b0000000000000000;
	sram_mem[104713] = 16'b0000000000000000;
	sram_mem[104714] = 16'b0000000000000000;
	sram_mem[104715] = 16'b0000000000000000;
	sram_mem[104716] = 16'b0000000000000000;
	sram_mem[104717] = 16'b0000000000000000;
	sram_mem[104718] = 16'b0000000000000000;
	sram_mem[104719] = 16'b0000000000000000;
	sram_mem[104720] = 16'b0000000000000000;
	sram_mem[104721] = 16'b0000000000000000;
	sram_mem[104722] = 16'b0000000000000000;
	sram_mem[104723] = 16'b0000000000000000;
	sram_mem[104724] = 16'b0000000000000000;
	sram_mem[104725] = 16'b0000000000000000;
	sram_mem[104726] = 16'b0000000000000000;
	sram_mem[104727] = 16'b0000000000000000;
	sram_mem[104728] = 16'b0000000000000000;
	sram_mem[104729] = 16'b0000000000000000;
	sram_mem[104730] = 16'b0000000000000000;
	sram_mem[104731] = 16'b0000000000000000;
	sram_mem[104732] = 16'b0000000000000000;
	sram_mem[104733] = 16'b0000000000000000;
	sram_mem[104734] = 16'b0000000000000000;
	sram_mem[104735] = 16'b0000000000000000;
	sram_mem[104736] = 16'b0000000000000000;
	sram_mem[104737] = 16'b0000000000000000;
	sram_mem[104738] = 16'b0000000000000000;
	sram_mem[104739] = 16'b0000000000000000;
	sram_mem[104740] = 16'b0000000000000000;
	sram_mem[104741] = 16'b0000000000000000;
	sram_mem[104742] = 16'b0000000000000000;
	sram_mem[104743] = 16'b0000000000000000;
	sram_mem[104744] = 16'b0000000000000000;
	sram_mem[104745] = 16'b0000000000000000;
	sram_mem[104746] = 16'b0000000000000000;
	sram_mem[104747] = 16'b0000000000000000;
	sram_mem[104748] = 16'b0000000000000000;
	sram_mem[104749] = 16'b0000000000000000;
	sram_mem[104750] = 16'b0000000000000000;
	sram_mem[104751] = 16'b0000000000000000;
	sram_mem[104752] = 16'b0000000000000000;
	sram_mem[104753] = 16'b0000000000000000;
	sram_mem[104754] = 16'b0000000000000000;
	sram_mem[104755] = 16'b0000000000000000;
	sram_mem[104756] = 16'b0000000000000000;
	sram_mem[104757] = 16'b0000000000000000;
	sram_mem[104758] = 16'b0000000000000000;
	sram_mem[104759] = 16'b0000000000000000;
	sram_mem[104760] = 16'b0000000000000000;
	sram_mem[104761] = 16'b0000000000000000;
	sram_mem[104762] = 16'b0000000000000000;
	sram_mem[104763] = 16'b0000000000000000;
	sram_mem[104764] = 16'b0000000000000000;
	sram_mem[104765] = 16'b0000000000000000;
	sram_mem[104766] = 16'b0000000000000000;
	sram_mem[104767] = 16'b0000000000000000;
	sram_mem[104768] = 16'b0000000000000000;
	sram_mem[104769] = 16'b0000000000000000;
	sram_mem[104770] = 16'b0000000000000000;
	sram_mem[104771] = 16'b0000000000000000;
	sram_mem[104772] = 16'b0000000000000000;
	sram_mem[104773] = 16'b0000000000000000;
	sram_mem[104774] = 16'b0000000000000000;
	sram_mem[104775] = 16'b0000000000000000;
	sram_mem[104776] = 16'b0000000000000000;
	sram_mem[104777] = 16'b0000000000000000;
	sram_mem[104778] = 16'b0000000000000000;
	sram_mem[104779] = 16'b0000000000000000;
	sram_mem[104780] = 16'b0000000000000000;
	sram_mem[104781] = 16'b0000000000000000;
	sram_mem[104782] = 16'b0000000000000000;
	sram_mem[104783] = 16'b0000000000000000;
	sram_mem[104784] = 16'b0000000000000000;
	sram_mem[104785] = 16'b0000000000000000;
	sram_mem[104786] = 16'b0000000000000000;
	sram_mem[104787] = 16'b0000000000000000;
	sram_mem[104788] = 16'b0000000000000000;
	sram_mem[104789] = 16'b0000000000000000;
	sram_mem[104790] = 16'b0000000000000000;
	sram_mem[104791] = 16'b0000000000000000;
	sram_mem[104792] = 16'b0000000000000000;
	sram_mem[104793] = 16'b0000000000000000;
	sram_mem[104794] = 16'b0000000000000000;
	sram_mem[104795] = 16'b0000000000000000;
	sram_mem[104796] = 16'b0000000000000000;
	sram_mem[104797] = 16'b0000000000000000;
	sram_mem[104798] = 16'b0000000000000000;
	sram_mem[104799] = 16'b0000000000000000;
	sram_mem[104800] = 16'b0000000000000000;
	sram_mem[104801] = 16'b0000000000000000;
	sram_mem[104802] = 16'b0000000000000000;
	sram_mem[104803] = 16'b0000000000000000;
	sram_mem[104804] = 16'b0000000000000000;
	sram_mem[104805] = 16'b0000000000000000;
	sram_mem[104806] = 16'b0000000000000000;
	sram_mem[104807] = 16'b0000000000000000;
	sram_mem[104808] = 16'b0000000000000000;
	sram_mem[104809] = 16'b0000000000000000;
	sram_mem[104810] = 16'b0000000000000000;
	sram_mem[104811] = 16'b0000000000000000;
	sram_mem[104812] = 16'b0000000000000000;
	sram_mem[104813] = 16'b0000000000000000;
	sram_mem[104814] = 16'b0000000000000000;
	sram_mem[104815] = 16'b0000000000000000;
	sram_mem[104816] = 16'b0000000000000000;
	sram_mem[104817] = 16'b0000000000000000;
	sram_mem[104818] = 16'b0000000000000000;
	sram_mem[104819] = 16'b0000000000000000;
	sram_mem[104820] = 16'b0000000000000000;
	sram_mem[104821] = 16'b0000000000000000;
	sram_mem[104822] = 16'b0000000000000000;
	sram_mem[104823] = 16'b0000000000000000;
	sram_mem[104824] = 16'b0000000000000000;
	sram_mem[104825] = 16'b0000000000000000;
	sram_mem[104826] = 16'b0000000000000000;
	sram_mem[104827] = 16'b0000000000000000;
	sram_mem[104828] = 16'b0000000000000000;
	sram_mem[104829] = 16'b0000000000000000;
	sram_mem[104830] = 16'b0000000000000000;
	sram_mem[104831] = 16'b0000000000000000;
	sram_mem[104832] = 16'b0000000000000000;
	sram_mem[104833] = 16'b0000000000000000;
	sram_mem[104834] = 16'b0000000000000000;
	sram_mem[104835] = 16'b0000000000000000;
	sram_mem[104836] = 16'b0000000000000000;
	sram_mem[104837] = 16'b0000000000000000;
	sram_mem[104838] = 16'b0000000000000000;
	sram_mem[104839] = 16'b0000000000000000;
	sram_mem[104840] = 16'b0000000000000000;
	sram_mem[104841] = 16'b0000000000000000;
	sram_mem[104842] = 16'b0000000000000000;
	sram_mem[104843] = 16'b0000000000000000;
	sram_mem[104844] = 16'b0000000000000000;
	sram_mem[104845] = 16'b0000000000000000;
	sram_mem[104846] = 16'b0000000000000000;
	sram_mem[104847] = 16'b0000000000000000;
	sram_mem[104848] = 16'b0000000000000000;
	sram_mem[104849] = 16'b0000000000000000;
	sram_mem[104850] = 16'b0000000000000000;
	sram_mem[104851] = 16'b0000000000000000;
	sram_mem[104852] = 16'b0000000000000000;
	sram_mem[104853] = 16'b0000000000000000;
	sram_mem[104854] = 16'b0000000000000000;
	sram_mem[104855] = 16'b0000000000000000;
	sram_mem[104856] = 16'b0000000000000000;
	sram_mem[104857] = 16'b0000000000000000;
	sram_mem[104858] = 16'b0000000000000000;
	sram_mem[104859] = 16'b0000000000000000;
	sram_mem[104860] = 16'b0000000000000000;
	sram_mem[104861] = 16'b0000000000000000;
	sram_mem[104862] = 16'b0000000000000000;
	sram_mem[104863] = 16'b0000000000000000;
	sram_mem[104864] = 16'b0000000000000000;
	sram_mem[104865] = 16'b0000000000000000;
	sram_mem[104866] = 16'b0000000000000000;
	sram_mem[104867] = 16'b0000000000000000;
	sram_mem[104868] = 16'b0000000000000000;
	sram_mem[104869] = 16'b0000000000000000;
	sram_mem[104870] = 16'b0000000000000000;
	sram_mem[104871] = 16'b0000000000000000;
	sram_mem[104872] = 16'b0000000000000000;
	sram_mem[104873] = 16'b0000000000000000;
	sram_mem[104874] = 16'b0000000000000000;
	sram_mem[104875] = 16'b0000000000000000;
	sram_mem[104876] = 16'b0000000000000000;
	sram_mem[104877] = 16'b0000000000000000;
	sram_mem[104878] = 16'b0000000000000000;
	sram_mem[104879] = 16'b0000000000000000;
	sram_mem[104880] = 16'b0000000000000000;
	sram_mem[104881] = 16'b0000000000000000;
	sram_mem[104882] = 16'b0000000000000000;
	sram_mem[104883] = 16'b0000000000000000;
	sram_mem[104884] = 16'b0000000000000000;
	sram_mem[104885] = 16'b0000000000000000;
	sram_mem[104886] = 16'b0000000000000000;
	sram_mem[104887] = 16'b0000000000000000;
	sram_mem[104888] = 16'b0000000000000000;
	sram_mem[104889] = 16'b0000000000000000;
	sram_mem[104890] = 16'b0000000000000000;
	sram_mem[104891] = 16'b0000000000000000;
	sram_mem[104892] = 16'b0000000000000000;
	sram_mem[104893] = 16'b0000000000000000;
	sram_mem[104894] = 16'b0000000000000000;
	sram_mem[104895] = 16'b0000000000000000;
	sram_mem[104896] = 16'b0000000000000000;
	sram_mem[104897] = 16'b0000000000000000;
	sram_mem[104898] = 16'b0000000000000000;
	sram_mem[104899] = 16'b0000000000000000;
	sram_mem[104900] = 16'b0000000000000000;
	sram_mem[104901] = 16'b0000000000000000;
	sram_mem[104902] = 16'b0000000000000000;
	sram_mem[104903] = 16'b0000000000000000;
	sram_mem[104904] = 16'b0000000000000000;
	sram_mem[104905] = 16'b0000000000000000;
	sram_mem[104906] = 16'b0000000000000000;
	sram_mem[104907] = 16'b0000000000000000;
	sram_mem[104908] = 16'b0000000000000000;
	sram_mem[104909] = 16'b0000000000000000;
	sram_mem[104910] = 16'b0000000000000000;
	sram_mem[104911] = 16'b0000000000000000;
	sram_mem[104912] = 16'b0000000000000000;
	sram_mem[104913] = 16'b0000000000000000;
	sram_mem[104914] = 16'b0000000000000000;
	sram_mem[104915] = 16'b0000000000000000;
	sram_mem[104916] = 16'b0000000000000000;
	sram_mem[104917] = 16'b0000000000000000;
	sram_mem[104918] = 16'b0000000000000000;
	sram_mem[104919] = 16'b0000000000000000;
	sram_mem[104920] = 16'b0000000000000000;
	sram_mem[104921] = 16'b0000000000000000;
	sram_mem[104922] = 16'b0000000000000000;
	sram_mem[104923] = 16'b0000000000000000;
	sram_mem[104924] = 16'b0000000000000000;
	sram_mem[104925] = 16'b0000000000000000;
	sram_mem[104926] = 16'b0000000000000000;
	sram_mem[104927] = 16'b0000000000000000;
	sram_mem[104928] = 16'b0000000000000000;
	sram_mem[104929] = 16'b0000000000000000;
	sram_mem[104930] = 16'b0000000000000000;
	sram_mem[104931] = 16'b0000000000000000;
	sram_mem[104932] = 16'b0000000000000000;
	sram_mem[104933] = 16'b0000000000000000;
	sram_mem[104934] = 16'b0000000000000000;
	sram_mem[104935] = 16'b0000000000000000;
	sram_mem[104936] = 16'b0000000000000000;
	sram_mem[104937] = 16'b0000000000000000;
	sram_mem[104938] = 16'b0000000000000000;
	sram_mem[104939] = 16'b0000000000000000;
	sram_mem[104940] = 16'b0000000000000000;
	sram_mem[104941] = 16'b0000000000000000;
	sram_mem[104942] = 16'b0000000000000000;
	sram_mem[104943] = 16'b0000000000000000;
	sram_mem[104944] = 16'b0000000000000000;
	sram_mem[104945] = 16'b0000000000000000;
	sram_mem[104946] = 16'b0000000000000000;
	sram_mem[104947] = 16'b0000000000000000;
	sram_mem[104948] = 16'b0000000000000000;
	sram_mem[104949] = 16'b0000000000000000;
	sram_mem[104950] = 16'b0000000000000000;
	sram_mem[104951] = 16'b0000000000000000;
	sram_mem[104952] = 16'b0000000000000000;
	sram_mem[104953] = 16'b0000000000000000;
	sram_mem[104954] = 16'b0000000000000000;
	sram_mem[104955] = 16'b0000000000000000;
	sram_mem[104956] = 16'b0000000000000000;
	sram_mem[104957] = 16'b0000000000000000;
	sram_mem[104958] = 16'b0000000000000000;
	sram_mem[104959] = 16'b0000000000000000;
	sram_mem[104960] = 16'b0000000000000000;
	sram_mem[104961] = 16'b0000000000000000;
	sram_mem[104962] = 16'b0000000000000000;
	sram_mem[104963] = 16'b0000000000000000;
	sram_mem[104964] = 16'b0000000000000000;
	sram_mem[104965] = 16'b0000000000000000;
	sram_mem[104966] = 16'b0000000000000000;
	sram_mem[104967] = 16'b0000000000000000;
	sram_mem[104968] = 16'b0000000000000000;
	sram_mem[104969] = 16'b0000000000000000;
	sram_mem[104970] = 16'b0000000000000000;
	sram_mem[104971] = 16'b0000000000000000;
	sram_mem[104972] = 16'b0000000000000000;
	sram_mem[104973] = 16'b0000000000000000;
	sram_mem[104974] = 16'b0000000000000000;
	sram_mem[104975] = 16'b0000000000000000;
	sram_mem[104976] = 16'b0000000000000000;
	sram_mem[104977] = 16'b0000000000000000;
	sram_mem[104978] = 16'b0000000000000000;
	sram_mem[104979] = 16'b0000000000000000;
	sram_mem[104980] = 16'b0000000000000000;
	sram_mem[104981] = 16'b0000000000000000;
	sram_mem[104982] = 16'b0000000000000000;
	sram_mem[104983] = 16'b0000000000000000;
	sram_mem[104984] = 16'b0000000000000000;
	sram_mem[104985] = 16'b0000000000000000;
	sram_mem[104986] = 16'b0000000000000000;
	sram_mem[104987] = 16'b0000000000000000;
	sram_mem[104988] = 16'b0000000000000000;
	sram_mem[104989] = 16'b0000000000000000;
	sram_mem[104990] = 16'b0000000000000000;
	sram_mem[104991] = 16'b0000000000000000;
	sram_mem[104992] = 16'b0000000000000000;
	sram_mem[104993] = 16'b0000000000000000;
	sram_mem[104994] = 16'b0000000000000000;
	sram_mem[104995] = 16'b0000000000000000;
	sram_mem[104996] = 16'b0000000000000000;
	sram_mem[104997] = 16'b0000000000000000;
	sram_mem[104998] = 16'b0000000000000000;
	sram_mem[104999] = 16'b0000000000000000;
	sram_mem[105000] = 16'b0000000000000000;
	sram_mem[105001] = 16'b0000000000000000;
	sram_mem[105002] = 16'b0000000000000000;
	sram_mem[105003] = 16'b0000000000000000;
	sram_mem[105004] = 16'b0000000000000000;
	sram_mem[105005] = 16'b0000000000000000;
	sram_mem[105006] = 16'b0000000000000000;
	sram_mem[105007] = 16'b0000000000000000;
	sram_mem[105008] = 16'b0000000000000000;
	sram_mem[105009] = 16'b0000000000000000;
	sram_mem[105010] = 16'b0000000000000000;
	sram_mem[105011] = 16'b0000000000000000;
	sram_mem[105012] = 16'b0000000000000000;
	sram_mem[105013] = 16'b0000000000000000;
	sram_mem[105014] = 16'b0000000000000000;
	sram_mem[105015] = 16'b0000000000000000;
	sram_mem[105016] = 16'b0000000000000000;
	sram_mem[105017] = 16'b0000000000000000;
	sram_mem[105018] = 16'b0000000000000000;
	sram_mem[105019] = 16'b0000000000000000;
	sram_mem[105020] = 16'b0000000000000000;
	sram_mem[105021] = 16'b0000000000000000;
	sram_mem[105022] = 16'b0000000000000000;
	sram_mem[105023] = 16'b0000000000000000;
	sram_mem[105024] = 16'b0000000000000000;
	sram_mem[105025] = 16'b0000000000000000;
	sram_mem[105026] = 16'b0000000000000000;
	sram_mem[105027] = 16'b0000000000000000;
	sram_mem[105028] = 16'b0000000000000000;
	sram_mem[105029] = 16'b0000000000000000;
	sram_mem[105030] = 16'b0000000000000000;
	sram_mem[105031] = 16'b0000000000000000;
	sram_mem[105032] = 16'b0000000000000000;
	sram_mem[105033] = 16'b0000000000000000;
	sram_mem[105034] = 16'b0000000000000000;
	sram_mem[105035] = 16'b0000000000000000;
	sram_mem[105036] = 16'b0000000000000000;
	sram_mem[105037] = 16'b0000000000000000;
	sram_mem[105038] = 16'b0000000000000000;
	sram_mem[105039] = 16'b0000000000000000;
	sram_mem[105040] = 16'b0000000000000000;
	sram_mem[105041] = 16'b0000000000000000;
	sram_mem[105042] = 16'b0000000000000000;
	sram_mem[105043] = 16'b0000000000000000;
	sram_mem[105044] = 16'b0000000000000000;
	sram_mem[105045] = 16'b0000000000000000;
	sram_mem[105046] = 16'b0000000000000000;
	sram_mem[105047] = 16'b0000000000000000;
	sram_mem[105048] = 16'b0000000000000000;
	sram_mem[105049] = 16'b0000000000000000;
	sram_mem[105050] = 16'b0000000000000000;
	sram_mem[105051] = 16'b0000000000000000;
	sram_mem[105052] = 16'b0000000000000000;
	sram_mem[105053] = 16'b0000000000000000;
	sram_mem[105054] = 16'b0000000000000000;
	sram_mem[105055] = 16'b0000000000000000;
	sram_mem[105056] = 16'b0000000000000000;
	sram_mem[105057] = 16'b0000000000000000;
	sram_mem[105058] = 16'b0000000000000000;
	sram_mem[105059] = 16'b0000000000000000;
	sram_mem[105060] = 16'b0000000000000000;
	sram_mem[105061] = 16'b0000000000000000;
	sram_mem[105062] = 16'b0000000000000000;
	sram_mem[105063] = 16'b0000000000000000;
	sram_mem[105064] = 16'b0000000000000000;
	sram_mem[105065] = 16'b0000000000000000;
	sram_mem[105066] = 16'b0000000000000000;
	sram_mem[105067] = 16'b0000000000000000;
	sram_mem[105068] = 16'b0000000000000000;
	sram_mem[105069] = 16'b0000000000000000;
	sram_mem[105070] = 16'b0000000000000000;
	sram_mem[105071] = 16'b0000000000000000;
	sram_mem[105072] = 16'b0000000000000000;
	sram_mem[105073] = 16'b0000000000000000;
	sram_mem[105074] = 16'b0000000000000000;
	sram_mem[105075] = 16'b0000000000000000;
	sram_mem[105076] = 16'b0000000000000000;
	sram_mem[105077] = 16'b0000000000000000;
	sram_mem[105078] = 16'b0000000000000000;
	sram_mem[105079] = 16'b0000000000000000;
	sram_mem[105080] = 16'b0000000000000000;
	sram_mem[105081] = 16'b0000000000000000;
	sram_mem[105082] = 16'b0000000000000000;
	sram_mem[105083] = 16'b0000000000000000;
	sram_mem[105084] = 16'b0000000000000000;
	sram_mem[105085] = 16'b0000000000000000;
	sram_mem[105086] = 16'b0000000000000000;
	sram_mem[105087] = 16'b0000000000000000;
	sram_mem[105088] = 16'b0000000000000000;
	sram_mem[105089] = 16'b0000000000000000;
	sram_mem[105090] = 16'b0000000000000000;
	sram_mem[105091] = 16'b0000000000000000;
	sram_mem[105092] = 16'b0000000000000000;
	sram_mem[105093] = 16'b0000000000000000;
	sram_mem[105094] = 16'b0000000000000000;
	sram_mem[105095] = 16'b0000000000000000;
	sram_mem[105096] = 16'b0000000000000000;
	sram_mem[105097] = 16'b0000000000000000;
	sram_mem[105098] = 16'b0000000000000000;
	sram_mem[105099] = 16'b0000000000000000;
	sram_mem[105100] = 16'b0000000000000000;
	sram_mem[105101] = 16'b0000000000000000;
	sram_mem[105102] = 16'b0000000000000000;
	sram_mem[105103] = 16'b0000000000000000;
	sram_mem[105104] = 16'b0000000000000000;
	sram_mem[105105] = 16'b0000000000000000;
	sram_mem[105106] = 16'b0000000000000000;
	sram_mem[105107] = 16'b0000000000000000;
	sram_mem[105108] = 16'b0000000000000000;
	sram_mem[105109] = 16'b0000000000000000;
	sram_mem[105110] = 16'b0000000000000000;
	sram_mem[105111] = 16'b0000000000000000;
	sram_mem[105112] = 16'b0000000000000000;
	sram_mem[105113] = 16'b0000000000000000;
	sram_mem[105114] = 16'b0000000000000000;
	sram_mem[105115] = 16'b0000000000000000;
	sram_mem[105116] = 16'b0000000000000000;
	sram_mem[105117] = 16'b0000000000000000;
	sram_mem[105118] = 16'b0000000000000000;
	sram_mem[105119] = 16'b0000000000000000;
	sram_mem[105120] = 16'b0000000000000000;
	sram_mem[105121] = 16'b0000000000000000;
	sram_mem[105122] = 16'b0000000000000000;
	sram_mem[105123] = 16'b0000000000000000;
	sram_mem[105124] = 16'b0000000000000000;
	sram_mem[105125] = 16'b0000000000000000;
	sram_mem[105126] = 16'b0000000000000000;
	sram_mem[105127] = 16'b0000000000000000;
	sram_mem[105128] = 16'b0000000000000000;
	sram_mem[105129] = 16'b0000000000000000;
	sram_mem[105130] = 16'b0000000000000000;
	sram_mem[105131] = 16'b0000000000000000;
	sram_mem[105132] = 16'b0000000000000000;
	sram_mem[105133] = 16'b0000000000000000;
	sram_mem[105134] = 16'b0000000000000000;
	sram_mem[105135] = 16'b0000000000000000;
	sram_mem[105136] = 16'b0000000000000000;
	sram_mem[105137] = 16'b0000000000000000;
	sram_mem[105138] = 16'b0000000000000000;
	sram_mem[105139] = 16'b0000000000000000;
	sram_mem[105140] = 16'b0000000000000000;
	sram_mem[105141] = 16'b0000000000000000;
	sram_mem[105142] = 16'b0000000000000000;
	sram_mem[105143] = 16'b0000000000000000;
	sram_mem[105144] = 16'b0000000000000000;
	sram_mem[105145] = 16'b0000000000000000;
	sram_mem[105146] = 16'b0000000000000000;
	sram_mem[105147] = 16'b0000000000000000;
	sram_mem[105148] = 16'b0000000000000000;
	sram_mem[105149] = 16'b0000000000000000;
	sram_mem[105150] = 16'b0000000000000000;
	sram_mem[105151] = 16'b0000000000000000;
	sram_mem[105152] = 16'b0000000000000000;
	sram_mem[105153] = 16'b0000000000000000;
	sram_mem[105154] = 16'b0000000000000000;
	sram_mem[105155] = 16'b0000000000000000;
	sram_mem[105156] = 16'b0000000000000000;
	sram_mem[105157] = 16'b0000000000000000;
	sram_mem[105158] = 16'b0000000000000000;
	sram_mem[105159] = 16'b0000000000000000;
	sram_mem[105160] = 16'b0000000000000000;
	sram_mem[105161] = 16'b0000000000000000;
	sram_mem[105162] = 16'b0000000000000000;
	sram_mem[105163] = 16'b0000000000000000;
	sram_mem[105164] = 16'b0000000000000000;
	sram_mem[105165] = 16'b0000000000000000;
	sram_mem[105166] = 16'b0000000000000000;
	sram_mem[105167] = 16'b0000000000000000;
	sram_mem[105168] = 16'b0000000000000000;
	sram_mem[105169] = 16'b0000000000000000;
	sram_mem[105170] = 16'b0000000000000000;
	sram_mem[105171] = 16'b0000000000000000;
	sram_mem[105172] = 16'b0000000000000000;
	sram_mem[105173] = 16'b0000000000000000;
	sram_mem[105174] = 16'b0000000000000000;
	sram_mem[105175] = 16'b0000000000000000;
	sram_mem[105176] = 16'b0000000000000000;
	sram_mem[105177] = 16'b0000000000000000;
	sram_mem[105178] = 16'b0000000000000000;
	sram_mem[105179] = 16'b0000000000000000;
	sram_mem[105180] = 16'b0000000000000000;
	sram_mem[105181] = 16'b0000000000000000;
	sram_mem[105182] = 16'b0000000000000000;
	sram_mem[105183] = 16'b0000000000000000;
	sram_mem[105184] = 16'b0000000000000000;
	sram_mem[105185] = 16'b0000000000000000;
	sram_mem[105186] = 16'b0000000000000000;
	sram_mem[105187] = 16'b0000000000000000;
	sram_mem[105188] = 16'b0000000000000000;
	sram_mem[105189] = 16'b0000000000000000;
	sram_mem[105190] = 16'b0000000000000000;
	sram_mem[105191] = 16'b0000000000000000;
	sram_mem[105192] = 16'b0000000000000000;
	sram_mem[105193] = 16'b0000000000000000;
	sram_mem[105194] = 16'b0000000000000000;
	sram_mem[105195] = 16'b0000000000000000;
	sram_mem[105196] = 16'b0000000000000000;
	sram_mem[105197] = 16'b0000000000000000;
	sram_mem[105198] = 16'b0000000000000000;
	sram_mem[105199] = 16'b0000000000000000;
	sram_mem[105200] = 16'b0000000000000000;
	sram_mem[105201] = 16'b0000000000000000;
	sram_mem[105202] = 16'b0000000000000000;
	sram_mem[105203] = 16'b0000000000000000;
	sram_mem[105204] = 16'b0000000000000000;
	sram_mem[105205] = 16'b0000000000000000;
	sram_mem[105206] = 16'b0000000000000000;
	sram_mem[105207] = 16'b0000000000000000;
	sram_mem[105208] = 16'b0000000000000000;
	sram_mem[105209] = 16'b0000000000000000;
	sram_mem[105210] = 16'b0000000000000000;
	sram_mem[105211] = 16'b0000000000000000;
	sram_mem[105212] = 16'b0000000000000000;
	sram_mem[105213] = 16'b0000000000000000;
	sram_mem[105214] = 16'b0000000000000000;
	sram_mem[105215] = 16'b0000000000000000;
	sram_mem[105216] = 16'b0000000000000000;
	sram_mem[105217] = 16'b0000000000000000;
	sram_mem[105218] = 16'b0000000000000000;
	sram_mem[105219] = 16'b0000000000000000;
	sram_mem[105220] = 16'b0000000000000000;
	sram_mem[105221] = 16'b0000000000000000;
	sram_mem[105222] = 16'b0000000000000000;
	sram_mem[105223] = 16'b0000000000000000;
	sram_mem[105224] = 16'b0000000000000000;
	sram_mem[105225] = 16'b0000000000000000;
	sram_mem[105226] = 16'b0000000000000000;
	sram_mem[105227] = 16'b0000000000000000;
	sram_mem[105228] = 16'b0000000000000000;
	sram_mem[105229] = 16'b0000000000000000;
	sram_mem[105230] = 16'b0000000000000000;
	sram_mem[105231] = 16'b0000000000000000;
	sram_mem[105232] = 16'b0000000000000000;
	sram_mem[105233] = 16'b0000000000000000;
	sram_mem[105234] = 16'b0000000000000000;
	sram_mem[105235] = 16'b0000000000000000;
	sram_mem[105236] = 16'b0000000000000000;
	sram_mem[105237] = 16'b0000000000000000;
	sram_mem[105238] = 16'b0000000000000000;
	sram_mem[105239] = 16'b0000000000000000;
	sram_mem[105240] = 16'b0000000000000000;
	sram_mem[105241] = 16'b0000000000000000;
	sram_mem[105242] = 16'b0000000000000000;
	sram_mem[105243] = 16'b0000000000000000;
	sram_mem[105244] = 16'b0000000000000000;
	sram_mem[105245] = 16'b0000000000000000;
	sram_mem[105246] = 16'b0000000000000000;
	sram_mem[105247] = 16'b0000000000000000;
	sram_mem[105248] = 16'b0000000000000000;
	sram_mem[105249] = 16'b0000000000000000;
	sram_mem[105250] = 16'b0000000000000000;
	sram_mem[105251] = 16'b0000000000000000;
	sram_mem[105252] = 16'b0000000000000000;
	sram_mem[105253] = 16'b0000000000000000;
	sram_mem[105254] = 16'b0000000000000000;
	sram_mem[105255] = 16'b0000000000000000;
	sram_mem[105256] = 16'b0000000000000000;
	sram_mem[105257] = 16'b0000000000000000;
	sram_mem[105258] = 16'b0000000000000000;
	sram_mem[105259] = 16'b0000000000000000;
	sram_mem[105260] = 16'b0000000000000000;
	sram_mem[105261] = 16'b0000000000000000;
	sram_mem[105262] = 16'b0000000000000000;
	sram_mem[105263] = 16'b0000000000000000;
	sram_mem[105264] = 16'b0000000000000000;
	sram_mem[105265] = 16'b0000000000000000;
	sram_mem[105266] = 16'b0000000000000000;
	sram_mem[105267] = 16'b0000000000000000;
	sram_mem[105268] = 16'b0000000000000000;
	sram_mem[105269] = 16'b0000000000000000;
	sram_mem[105270] = 16'b0000000000000000;
	sram_mem[105271] = 16'b0000000000000000;
	sram_mem[105272] = 16'b0000000000000000;
	sram_mem[105273] = 16'b0000000000000000;
	sram_mem[105274] = 16'b0000000000000000;
	sram_mem[105275] = 16'b0000000000000000;
	sram_mem[105276] = 16'b0000000000000000;
	sram_mem[105277] = 16'b0000000000000000;
	sram_mem[105278] = 16'b0000000000000000;
	sram_mem[105279] = 16'b0000000000000000;
	sram_mem[105280] = 16'b0000000000000000;
	sram_mem[105281] = 16'b0000000000000000;
	sram_mem[105282] = 16'b0000000000000000;
	sram_mem[105283] = 16'b0000000000000000;
	sram_mem[105284] = 16'b0000000000000000;
	sram_mem[105285] = 16'b0000000000000000;
	sram_mem[105286] = 16'b0000000000000000;
	sram_mem[105287] = 16'b0000000000000000;
	sram_mem[105288] = 16'b0000000000000000;
	sram_mem[105289] = 16'b0000000000000000;
	sram_mem[105290] = 16'b0000000000000000;
	sram_mem[105291] = 16'b0000000000000000;
	sram_mem[105292] = 16'b0000000000000000;
	sram_mem[105293] = 16'b0000000000000000;
	sram_mem[105294] = 16'b0000000000000000;
	sram_mem[105295] = 16'b0000000000000000;
	sram_mem[105296] = 16'b0000000000000000;
	sram_mem[105297] = 16'b0000000000000000;
	sram_mem[105298] = 16'b0000000000000000;
	sram_mem[105299] = 16'b0000000000000000;
	sram_mem[105300] = 16'b0000000000000000;
	sram_mem[105301] = 16'b0000000000000000;
	sram_mem[105302] = 16'b0000000000000000;
	sram_mem[105303] = 16'b0000000000000000;
	sram_mem[105304] = 16'b0000000000000000;
	sram_mem[105305] = 16'b0000000000000000;
	sram_mem[105306] = 16'b0000000000000000;
	sram_mem[105307] = 16'b0000000000000000;
	sram_mem[105308] = 16'b0000000000000000;
	sram_mem[105309] = 16'b0000000000000000;
	sram_mem[105310] = 16'b0000000000000000;
	sram_mem[105311] = 16'b0000000000000000;
	sram_mem[105312] = 16'b0000000000000000;
	sram_mem[105313] = 16'b0000000000000000;
	sram_mem[105314] = 16'b0000000000000000;
	sram_mem[105315] = 16'b0000000000000000;
	sram_mem[105316] = 16'b0000000000000000;
	sram_mem[105317] = 16'b0000000000000000;
	sram_mem[105318] = 16'b0000000000000000;
	sram_mem[105319] = 16'b0000000000000000;
	sram_mem[105320] = 16'b0000000000000000;
	sram_mem[105321] = 16'b0000000000000000;
	sram_mem[105322] = 16'b0000000000000000;
	sram_mem[105323] = 16'b0000000000000000;
	sram_mem[105324] = 16'b0000000000000000;
	sram_mem[105325] = 16'b0000000000000000;
	sram_mem[105326] = 16'b0000000000000000;
	sram_mem[105327] = 16'b0000000000000000;
	sram_mem[105328] = 16'b0000000000000000;
	sram_mem[105329] = 16'b0000000000000000;
	sram_mem[105330] = 16'b0000000000000000;
	sram_mem[105331] = 16'b0000000000000000;
	sram_mem[105332] = 16'b0000000000000000;
	sram_mem[105333] = 16'b0000000000000000;
	sram_mem[105334] = 16'b0000000000000000;
	sram_mem[105335] = 16'b0000000000000000;
	sram_mem[105336] = 16'b0000000000000000;
	sram_mem[105337] = 16'b0000000000000000;
	sram_mem[105338] = 16'b0000000000000000;
	sram_mem[105339] = 16'b0000000000000000;
	sram_mem[105340] = 16'b0000000000000000;
	sram_mem[105341] = 16'b0000000000000000;
	sram_mem[105342] = 16'b0000000000000000;
	sram_mem[105343] = 16'b0000000000000000;
	sram_mem[105344] = 16'b0000000000000000;
	sram_mem[105345] = 16'b0000000000000000;
	sram_mem[105346] = 16'b0000000000000000;
	sram_mem[105347] = 16'b0000000000000000;
	sram_mem[105348] = 16'b0000000000000000;
	sram_mem[105349] = 16'b0000000000000000;
	sram_mem[105350] = 16'b0000000000000000;
	sram_mem[105351] = 16'b0000000000000000;
	sram_mem[105352] = 16'b0000000000000000;
	sram_mem[105353] = 16'b0000000000000000;
	sram_mem[105354] = 16'b0000000000000000;
	sram_mem[105355] = 16'b0000000000000000;
	sram_mem[105356] = 16'b0000000000000000;
	sram_mem[105357] = 16'b0000000000000000;
	sram_mem[105358] = 16'b0000000000000000;
	sram_mem[105359] = 16'b0000000000000000;
	sram_mem[105360] = 16'b0000000000000000;
	sram_mem[105361] = 16'b0000000000000000;
	sram_mem[105362] = 16'b0000000000000000;
	sram_mem[105363] = 16'b0000000000000000;
	sram_mem[105364] = 16'b0000000000000000;
	sram_mem[105365] = 16'b0000000000000000;
	sram_mem[105366] = 16'b0000000000000000;
	sram_mem[105367] = 16'b0000000000000000;
	sram_mem[105368] = 16'b0000000000000000;
	sram_mem[105369] = 16'b0000000000000000;
	sram_mem[105370] = 16'b0000000000000000;
	sram_mem[105371] = 16'b0000000000000000;
	sram_mem[105372] = 16'b0000000000000000;
	sram_mem[105373] = 16'b0000000000000000;
	sram_mem[105374] = 16'b0000000000000000;
	sram_mem[105375] = 16'b0000000000000000;
	sram_mem[105376] = 16'b0000000000000000;
	sram_mem[105377] = 16'b0000000000000000;
	sram_mem[105378] = 16'b0000000000000000;
	sram_mem[105379] = 16'b0000000000000000;
	sram_mem[105380] = 16'b0000000000000000;
	sram_mem[105381] = 16'b0000000000000000;
	sram_mem[105382] = 16'b0000000000000000;
	sram_mem[105383] = 16'b0000000000000000;
	sram_mem[105384] = 16'b0000000000000000;
	sram_mem[105385] = 16'b0000000000000000;
	sram_mem[105386] = 16'b0000000000000000;
	sram_mem[105387] = 16'b0000000000000000;
	sram_mem[105388] = 16'b0000000000000000;
	sram_mem[105389] = 16'b0000000000000000;
	sram_mem[105390] = 16'b0000000000000000;
	sram_mem[105391] = 16'b0000000000000000;
	sram_mem[105392] = 16'b0000000000000000;
	sram_mem[105393] = 16'b0000000000000000;
	sram_mem[105394] = 16'b0000000000000000;
	sram_mem[105395] = 16'b0000000000000000;
	sram_mem[105396] = 16'b0000000000000000;
	sram_mem[105397] = 16'b0000000000000000;
	sram_mem[105398] = 16'b0000000000000000;
	sram_mem[105399] = 16'b0000000000000000;
	sram_mem[105400] = 16'b0000000000000000;
	sram_mem[105401] = 16'b0000000000000000;
	sram_mem[105402] = 16'b0000000000000000;
	sram_mem[105403] = 16'b0000000000000000;
	sram_mem[105404] = 16'b0000000000000000;
	sram_mem[105405] = 16'b0000000000000000;
	sram_mem[105406] = 16'b0000000000000000;
	sram_mem[105407] = 16'b0000000000000000;
	sram_mem[105408] = 16'b0000000000000000;
	sram_mem[105409] = 16'b0000000000000000;
	sram_mem[105410] = 16'b0000000000000000;
	sram_mem[105411] = 16'b0000000000000000;
	sram_mem[105412] = 16'b0000000000000000;
	sram_mem[105413] = 16'b0000000000000000;
	sram_mem[105414] = 16'b0000000000000000;
	sram_mem[105415] = 16'b0000000000000000;
	sram_mem[105416] = 16'b0000000000000000;
	sram_mem[105417] = 16'b0000000000000000;
	sram_mem[105418] = 16'b0000000000000000;
	sram_mem[105419] = 16'b0000000000000000;
	sram_mem[105420] = 16'b0000000000000000;
	sram_mem[105421] = 16'b0000000000000000;
	sram_mem[105422] = 16'b0000000000000000;
	sram_mem[105423] = 16'b0000000000000000;
	sram_mem[105424] = 16'b0000000000000000;
	sram_mem[105425] = 16'b0000000000000000;
	sram_mem[105426] = 16'b0000000000000000;
	sram_mem[105427] = 16'b0000000000000000;
	sram_mem[105428] = 16'b0000000000000000;
	sram_mem[105429] = 16'b0000000000000000;
	sram_mem[105430] = 16'b0000000000000000;
	sram_mem[105431] = 16'b0000000000000000;
	sram_mem[105432] = 16'b0000000000000000;
	sram_mem[105433] = 16'b0000000000000000;
	sram_mem[105434] = 16'b0000000000000000;
	sram_mem[105435] = 16'b0000000000000000;
	sram_mem[105436] = 16'b0000000000000000;
	sram_mem[105437] = 16'b0000000000000000;
	sram_mem[105438] = 16'b0000000000000000;
	sram_mem[105439] = 16'b0000000000000000;
	sram_mem[105440] = 16'b0000000000000000;
	sram_mem[105441] = 16'b0000000000000000;
	sram_mem[105442] = 16'b0000000000000000;
	sram_mem[105443] = 16'b0000000000000000;
	sram_mem[105444] = 16'b0000000000000000;
	sram_mem[105445] = 16'b0000000000000000;
	sram_mem[105446] = 16'b0000000000000000;
	sram_mem[105447] = 16'b0000000000000000;
	sram_mem[105448] = 16'b0000000000000000;
	sram_mem[105449] = 16'b0000000000000000;
	sram_mem[105450] = 16'b0000000000000000;
	sram_mem[105451] = 16'b0000000000000000;
	sram_mem[105452] = 16'b0000000000000000;
	sram_mem[105453] = 16'b0000000000000000;
	sram_mem[105454] = 16'b0000000000000000;
	sram_mem[105455] = 16'b0000000000000000;
	sram_mem[105456] = 16'b0000000000000000;
	sram_mem[105457] = 16'b0000000000000000;
	sram_mem[105458] = 16'b0000000000000000;
	sram_mem[105459] = 16'b0000000000000000;
	sram_mem[105460] = 16'b0000000000000000;
	sram_mem[105461] = 16'b0000000000000000;
	sram_mem[105462] = 16'b0000000000000000;
	sram_mem[105463] = 16'b0000000000000000;
	sram_mem[105464] = 16'b0000000000000000;
	sram_mem[105465] = 16'b0000000000000000;
	sram_mem[105466] = 16'b0000000000000000;
	sram_mem[105467] = 16'b0000000000000000;
	sram_mem[105468] = 16'b0000000000000000;
	sram_mem[105469] = 16'b0000000000000000;
	sram_mem[105470] = 16'b0000000000000000;
	sram_mem[105471] = 16'b0000000000000000;
	sram_mem[105472] = 16'b0000000000000000;
	sram_mem[105473] = 16'b0000000000000000;
	sram_mem[105474] = 16'b0000000000000000;
	sram_mem[105475] = 16'b0000000000000000;
	sram_mem[105476] = 16'b0000000000000000;
	sram_mem[105477] = 16'b0000000000000000;
	sram_mem[105478] = 16'b0000000000000000;
	sram_mem[105479] = 16'b0000000000000000;
	sram_mem[105480] = 16'b0000000000000000;
	sram_mem[105481] = 16'b0000000000000000;
	sram_mem[105482] = 16'b0000000000000000;
	sram_mem[105483] = 16'b0000000000000000;
	sram_mem[105484] = 16'b0000000000000000;
	sram_mem[105485] = 16'b0000000000000000;
	sram_mem[105486] = 16'b0000000000000000;
	sram_mem[105487] = 16'b0000000000000000;
	sram_mem[105488] = 16'b0000000000000000;
	sram_mem[105489] = 16'b0000000000000000;
	sram_mem[105490] = 16'b0000000000000000;
	sram_mem[105491] = 16'b0000000000000000;
	sram_mem[105492] = 16'b0000000000000000;
	sram_mem[105493] = 16'b0000000000000000;
	sram_mem[105494] = 16'b0000000000000000;
	sram_mem[105495] = 16'b0000000000000000;
	sram_mem[105496] = 16'b0000000000000000;
	sram_mem[105497] = 16'b0000000000000000;
	sram_mem[105498] = 16'b0000000000000000;
	sram_mem[105499] = 16'b0000000000000000;
	sram_mem[105500] = 16'b0000000000000000;
	sram_mem[105501] = 16'b0000000000000000;
	sram_mem[105502] = 16'b0000000000000000;
	sram_mem[105503] = 16'b0000000000000000;
	sram_mem[105504] = 16'b0000000000000000;
	sram_mem[105505] = 16'b0000000000000000;
	sram_mem[105506] = 16'b0000000000000000;
	sram_mem[105507] = 16'b0000000000000000;
	sram_mem[105508] = 16'b0000000000000000;
	sram_mem[105509] = 16'b0000000000000000;
	sram_mem[105510] = 16'b0000000000000000;
	sram_mem[105511] = 16'b0000000000000000;
	sram_mem[105512] = 16'b0000000000000000;
	sram_mem[105513] = 16'b0000000000000000;
	sram_mem[105514] = 16'b0000000000000000;
	sram_mem[105515] = 16'b0000000000000000;
	sram_mem[105516] = 16'b0000000000000000;
	sram_mem[105517] = 16'b0000000000000000;
	sram_mem[105518] = 16'b0000000000000000;
	sram_mem[105519] = 16'b0000000000000000;
	sram_mem[105520] = 16'b0000000000000000;
	sram_mem[105521] = 16'b0000000000000000;
	sram_mem[105522] = 16'b0000000000000000;
	sram_mem[105523] = 16'b0000000000000000;
	sram_mem[105524] = 16'b0000000000000000;
	sram_mem[105525] = 16'b0000000000000000;
	sram_mem[105526] = 16'b0000000000000000;
	sram_mem[105527] = 16'b0000000000000000;
	sram_mem[105528] = 16'b0000000000000000;
	sram_mem[105529] = 16'b0000000000000000;
	sram_mem[105530] = 16'b0000000000000000;
	sram_mem[105531] = 16'b0000000000000000;
	sram_mem[105532] = 16'b0000000000000000;
	sram_mem[105533] = 16'b0000000000000000;
	sram_mem[105534] = 16'b0000000000000000;
	sram_mem[105535] = 16'b0000000000000000;
	sram_mem[105536] = 16'b0000000000000000;
	sram_mem[105537] = 16'b0000000000000000;
	sram_mem[105538] = 16'b0000000000000000;
	sram_mem[105539] = 16'b0000000000000000;
	sram_mem[105540] = 16'b0000000000000000;
	sram_mem[105541] = 16'b0000000000000000;
	sram_mem[105542] = 16'b0000000000000000;
	sram_mem[105543] = 16'b0000000000000000;
	sram_mem[105544] = 16'b0000000000000000;
	sram_mem[105545] = 16'b0000000000000000;
	sram_mem[105546] = 16'b0000000000000000;
	sram_mem[105547] = 16'b0000000000000000;
	sram_mem[105548] = 16'b0000000000000000;
	sram_mem[105549] = 16'b0000000000000000;
	sram_mem[105550] = 16'b0000000000000000;
	sram_mem[105551] = 16'b0000000000000000;
	sram_mem[105552] = 16'b0000000000000000;
	sram_mem[105553] = 16'b0000000000000000;
	sram_mem[105554] = 16'b0000000000000000;
	sram_mem[105555] = 16'b0000000000000000;
	sram_mem[105556] = 16'b0000000000000000;
	sram_mem[105557] = 16'b0000000000000000;
	sram_mem[105558] = 16'b0000000000000000;
	sram_mem[105559] = 16'b0000000000000000;
	sram_mem[105560] = 16'b0000000000000000;
	sram_mem[105561] = 16'b0000000000000000;
	sram_mem[105562] = 16'b0000000000000000;
	sram_mem[105563] = 16'b0000000000000000;
	sram_mem[105564] = 16'b0000000000000000;
	sram_mem[105565] = 16'b0000000000000000;
	sram_mem[105566] = 16'b0000000000000000;
	sram_mem[105567] = 16'b0000000000000000;
	sram_mem[105568] = 16'b0000000000000000;
	sram_mem[105569] = 16'b0000000000000000;
	sram_mem[105570] = 16'b0000000000000000;
	sram_mem[105571] = 16'b0000000000000000;
	sram_mem[105572] = 16'b0000000000000000;
	sram_mem[105573] = 16'b0000000000000000;
	sram_mem[105574] = 16'b0000000000000000;
	sram_mem[105575] = 16'b0000000000000000;
	sram_mem[105576] = 16'b0000000000000000;
	sram_mem[105577] = 16'b0000000000000000;
	sram_mem[105578] = 16'b0000000000000000;
	sram_mem[105579] = 16'b0000000000000000;
	sram_mem[105580] = 16'b0000000000000000;
	sram_mem[105581] = 16'b0000000000000000;
	sram_mem[105582] = 16'b0000000000000000;
	sram_mem[105583] = 16'b0000000000000000;
	sram_mem[105584] = 16'b0000000000000000;
	sram_mem[105585] = 16'b0000000000000000;
	sram_mem[105586] = 16'b0000000000000000;
	sram_mem[105587] = 16'b0000000000000000;
	sram_mem[105588] = 16'b0000000000000000;
	sram_mem[105589] = 16'b0000000000000000;
	sram_mem[105590] = 16'b0000000000000000;
	sram_mem[105591] = 16'b0000000000000000;
	sram_mem[105592] = 16'b0000000000000000;
	sram_mem[105593] = 16'b0000000000000000;
	sram_mem[105594] = 16'b0000000000000000;
	sram_mem[105595] = 16'b0000000000000000;
	sram_mem[105596] = 16'b0000000000000000;
	sram_mem[105597] = 16'b0000000000000000;
	sram_mem[105598] = 16'b0000000000000000;
	sram_mem[105599] = 16'b0000000000000000;
	sram_mem[105600] = 16'b0000000000000000;
	sram_mem[105601] = 16'b0000000000000000;
	sram_mem[105602] = 16'b0000000000000000;
	sram_mem[105603] = 16'b0000000000000000;
	sram_mem[105604] = 16'b0000000000000000;
	sram_mem[105605] = 16'b0000000000000000;
	sram_mem[105606] = 16'b0000000000000000;
	sram_mem[105607] = 16'b0000000000000000;
	sram_mem[105608] = 16'b0000000000000000;
	sram_mem[105609] = 16'b0000000000000000;
	sram_mem[105610] = 16'b0000000000000000;
	sram_mem[105611] = 16'b0000000000000000;
	sram_mem[105612] = 16'b0000000000000000;
	sram_mem[105613] = 16'b0000000000000000;
	sram_mem[105614] = 16'b0000000000000000;
	sram_mem[105615] = 16'b0000000000000000;
	sram_mem[105616] = 16'b0000000000000000;
	sram_mem[105617] = 16'b0000000000000000;
	sram_mem[105618] = 16'b0000000000000000;
	sram_mem[105619] = 16'b0000000000000000;
	sram_mem[105620] = 16'b0000000000000000;
	sram_mem[105621] = 16'b0000000000000000;
	sram_mem[105622] = 16'b0000000000000000;
	sram_mem[105623] = 16'b0000000000000000;
	sram_mem[105624] = 16'b0000000000000000;
	sram_mem[105625] = 16'b0000000000000000;
	sram_mem[105626] = 16'b0000000000000000;
	sram_mem[105627] = 16'b0000000000000000;
	sram_mem[105628] = 16'b0000000000000000;
	sram_mem[105629] = 16'b0000000000000000;
	sram_mem[105630] = 16'b0000000000000000;
	sram_mem[105631] = 16'b0000000000000000;
	sram_mem[105632] = 16'b0000000000000000;
	sram_mem[105633] = 16'b0000000000000000;
	sram_mem[105634] = 16'b0000000000000000;
	sram_mem[105635] = 16'b0000000000000000;
	sram_mem[105636] = 16'b0000000000000000;
	sram_mem[105637] = 16'b0000000000000000;
	sram_mem[105638] = 16'b0000000000000000;
	sram_mem[105639] = 16'b0000000000000000;
	sram_mem[105640] = 16'b0000000000000000;
	sram_mem[105641] = 16'b0000000000000000;
	sram_mem[105642] = 16'b0000000000000000;
	sram_mem[105643] = 16'b0000000000000000;
	sram_mem[105644] = 16'b0000000000000000;
	sram_mem[105645] = 16'b0000000000000000;
	sram_mem[105646] = 16'b0000000000000000;
	sram_mem[105647] = 16'b0000000000000000;
	sram_mem[105648] = 16'b0000000000000000;
	sram_mem[105649] = 16'b0000000000000000;
	sram_mem[105650] = 16'b0000000000000000;
	sram_mem[105651] = 16'b0000000000000000;
	sram_mem[105652] = 16'b0000000000000000;
	sram_mem[105653] = 16'b0000000000000000;
	sram_mem[105654] = 16'b0000000000000000;
	sram_mem[105655] = 16'b0000000000000000;
	sram_mem[105656] = 16'b0000000000000000;
	sram_mem[105657] = 16'b0000000000000000;
	sram_mem[105658] = 16'b0000000000000000;
	sram_mem[105659] = 16'b0000000000000000;
	sram_mem[105660] = 16'b0000000000000000;
	sram_mem[105661] = 16'b0000000000000000;
	sram_mem[105662] = 16'b0000000000000000;
	sram_mem[105663] = 16'b0000000000000000;
	sram_mem[105664] = 16'b0000000000000000;
	sram_mem[105665] = 16'b0000000000000000;
	sram_mem[105666] = 16'b0000000000000000;
	sram_mem[105667] = 16'b0000000000000000;
	sram_mem[105668] = 16'b0000000000000000;
	sram_mem[105669] = 16'b0000000000000000;
	sram_mem[105670] = 16'b0000000000000000;
	sram_mem[105671] = 16'b0000000000000000;
	sram_mem[105672] = 16'b0000000000000000;
	sram_mem[105673] = 16'b0000000000000000;
	sram_mem[105674] = 16'b0000000000000000;
	sram_mem[105675] = 16'b0000000000000000;
	sram_mem[105676] = 16'b0000000000000000;
	sram_mem[105677] = 16'b0000000000000000;
	sram_mem[105678] = 16'b0000000000000000;
	sram_mem[105679] = 16'b0000000000000000;
	sram_mem[105680] = 16'b0000000000000000;
	sram_mem[105681] = 16'b0000000000000000;
	sram_mem[105682] = 16'b0000000000000000;
	sram_mem[105683] = 16'b0000000000000000;
	sram_mem[105684] = 16'b0000000000000000;
	sram_mem[105685] = 16'b0000000000000000;
	sram_mem[105686] = 16'b0000000000000000;
	sram_mem[105687] = 16'b0000000000000000;
	sram_mem[105688] = 16'b0000000000000000;
	sram_mem[105689] = 16'b0000000000000000;
	sram_mem[105690] = 16'b0000000000000000;
	sram_mem[105691] = 16'b0000000000000000;
	sram_mem[105692] = 16'b0000000000000000;
	sram_mem[105693] = 16'b0000000000000000;
	sram_mem[105694] = 16'b0000000000000000;
	sram_mem[105695] = 16'b0000000000000000;
	sram_mem[105696] = 16'b0000000000000000;
	sram_mem[105697] = 16'b0000000000000000;
	sram_mem[105698] = 16'b0000000000000000;
	sram_mem[105699] = 16'b0000000000000000;
	sram_mem[105700] = 16'b0000000000000000;
	sram_mem[105701] = 16'b0000000000000000;
	sram_mem[105702] = 16'b0000000000000000;
	sram_mem[105703] = 16'b0000000000000000;
	sram_mem[105704] = 16'b0000000000000000;
	sram_mem[105705] = 16'b0000000000000000;
	sram_mem[105706] = 16'b0000000000000000;
	sram_mem[105707] = 16'b0000000000000000;
	sram_mem[105708] = 16'b0000000000000000;
	sram_mem[105709] = 16'b0000000000000000;
	sram_mem[105710] = 16'b0000000000000000;
	sram_mem[105711] = 16'b0000000000000000;
	sram_mem[105712] = 16'b0000000000000000;
	sram_mem[105713] = 16'b0000000000000000;
	sram_mem[105714] = 16'b0000000000000000;
	sram_mem[105715] = 16'b0000000000000000;
	sram_mem[105716] = 16'b0000000000000000;
	sram_mem[105717] = 16'b0000000000000000;
	sram_mem[105718] = 16'b0000000000000000;
	sram_mem[105719] = 16'b0000000000000000;
	sram_mem[105720] = 16'b0000000000000000;
	sram_mem[105721] = 16'b0000000000000000;
	sram_mem[105722] = 16'b0000000000000000;
	sram_mem[105723] = 16'b0000000000000000;
	sram_mem[105724] = 16'b0000000000000000;
	sram_mem[105725] = 16'b0000000000000000;
	sram_mem[105726] = 16'b0000000000000000;
	sram_mem[105727] = 16'b0000000000000000;
	sram_mem[105728] = 16'b0000000000000000;
	sram_mem[105729] = 16'b0000000000000000;
	sram_mem[105730] = 16'b0000000000000000;
	sram_mem[105731] = 16'b0000000000000000;
	sram_mem[105732] = 16'b0000000000000000;
	sram_mem[105733] = 16'b0000000000000000;
	sram_mem[105734] = 16'b0000000000000000;
	sram_mem[105735] = 16'b0000000000000000;
	sram_mem[105736] = 16'b0000000000000000;
	sram_mem[105737] = 16'b0000000000000000;
	sram_mem[105738] = 16'b0000000000000000;
	sram_mem[105739] = 16'b0000000000000000;
	sram_mem[105740] = 16'b0000000000000000;
	sram_mem[105741] = 16'b0000000000000000;
	sram_mem[105742] = 16'b0000000000000000;
	sram_mem[105743] = 16'b0000000000000000;
	sram_mem[105744] = 16'b0000000000000000;
	sram_mem[105745] = 16'b0000000000000000;
	sram_mem[105746] = 16'b0000000000000000;
	sram_mem[105747] = 16'b0000000000000000;
	sram_mem[105748] = 16'b0000000000000000;
	sram_mem[105749] = 16'b0000000000000000;
	sram_mem[105750] = 16'b0000000000000000;
	sram_mem[105751] = 16'b0000000000000000;
	sram_mem[105752] = 16'b0000000000000000;
	sram_mem[105753] = 16'b0000000000000000;
	sram_mem[105754] = 16'b0000000000000000;
	sram_mem[105755] = 16'b0000000000000000;
	sram_mem[105756] = 16'b0000000000000000;
	sram_mem[105757] = 16'b0000000000000000;
	sram_mem[105758] = 16'b0000000000000000;
	sram_mem[105759] = 16'b0000000000000000;
	sram_mem[105760] = 16'b0000000000000000;
	sram_mem[105761] = 16'b0000000000000000;
	sram_mem[105762] = 16'b0000000000000000;
	sram_mem[105763] = 16'b0000000000000000;
	sram_mem[105764] = 16'b0000000000000000;
	sram_mem[105765] = 16'b0000000000000000;
	sram_mem[105766] = 16'b0000000000000000;
	sram_mem[105767] = 16'b0000000000000000;
	sram_mem[105768] = 16'b0000000000000000;
	sram_mem[105769] = 16'b0000000000000000;
	sram_mem[105770] = 16'b0000000000000000;
	sram_mem[105771] = 16'b0000000000000000;
	sram_mem[105772] = 16'b0000000000000000;
	sram_mem[105773] = 16'b0000000000000000;
	sram_mem[105774] = 16'b0000000000000000;
	sram_mem[105775] = 16'b0000000000000000;
	sram_mem[105776] = 16'b0000000000000000;
	sram_mem[105777] = 16'b0000000000000000;
	sram_mem[105778] = 16'b0000000000000000;
	sram_mem[105779] = 16'b0000000000000000;
	sram_mem[105780] = 16'b0000000000000000;
	sram_mem[105781] = 16'b0000000000000000;
	sram_mem[105782] = 16'b0000000000000000;
	sram_mem[105783] = 16'b0000000000000000;
	sram_mem[105784] = 16'b0000000000000000;
	sram_mem[105785] = 16'b0000000000000000;
	sram_mem[105786] = 16'b0000000000000000;
	sram_mem[105787] = 16'b0000000000000000;
	sram_mem[105788] = 16'b0000000000000000;
	sram_mem[105789] = 16'b0000000000000000;
	sram_mem[105790] = 16'b0000000000000000;
	sram_mem[105791] = 16'b0000000000000000;
	sram_mem[105792] = 16'b0000000000000000;
	sram_mem[105793] = 16'b0000000000000000;
	sram_mem[105794] = 16'b0000000000000000;
	sram_mem[105795] = 16'b0000000000000000;
	sram_mem[105796] = 16'b0000000000000000;
	sram_mem[105797] = 16'b0000000000000000;
	sram_mem[105798] = 16'b0000000000000000;
	sram_mem[105799] = 16'b0000000000000000;
	sram_mem[105800] = 16'b0000000000000000;
	sram_mem[105801] = 16'b0000000000000000;
	sram_mem[105802] = 16'b0000000000000000;
	sram_mem[105803] = 16'b0000000000000000;
	sram_mem[105804] = 16'b0000000000000000;
	sram_mem[105805] = 16'b0000000000000000;
	sram_mem[105806] = 16'b0000000000000000;
	sram_mem[105807] = 16'b0000000000000000;
	sram_mem[105808] = 16'b0000000000000000;
	sram_mem[105809] = 16'b0000000000000000;
	sram_mem[105810] = 16'b0000000000000000;
	sram_mem[105811] = 16'b0000000000000000;
	sram_mem[105812] = 16'b0000000000000000;
	sram_mem[105813] = 16'b0000000000000000;
	sram_mem[105814] = 16'b0000000000000000;
	sram_mem[105815] = 16'b0000000000000000;
	sram_mem[105816] = 16'b0000000000000000;
	sram_mem[105817] = 16'b0000000000000000;
	sram_mem[105818] = 16'b0000000000000000;
	sram_mem[105819] = 16'b0000000000000000;
	sram_mem[105820] = 16'b0000000000000000;
	sram_mem[105821] = 16'b0000000000000000;
	sram_mem[105822] = 16'b0000000000000000;
	sram_mem[105823] = 16'b0000000000000000;
	sram_mem[105824] = 16'b0000000000000000;
	sram_mem[105825] = 16'b0000000000000000;
	sram_mem[105826] = 16'b0000000000000000;
	sram_mem[105827] = 16'b0000000000000000;
	sram_mem[105828] = 16'b0000000000000000;
	sram_mem[105829] = 16'b0000000000000000;
	sram_mem[105830] = 16'b0000000000000000;
	sram_mem[105831] = 16'b0000000000000000;
	sram_mem[105832] = 16'b0000000000000000;
	sram_mem[105833] = 16'b0000000000000000;
	sram_mem[105834] = 16'b0000000000000000;
	sram_mem[105835] = 16'b0000000000000000;
	sram_mem[105836] = 16'b0000000000000000;
	sram_mem[105837] = 16'b0000000000000000;
	sram_mem[105838] = 16'b0000000000000000;
	sram_mem[105839] = 16'b0000000000000000;
	sram_mem[105840] = 16'b0000000000000000;
	sram_mem[105841] = 16'b0000000000000000;
	sram_mem[105842] = 16'b0000000000000000;
	sram_mem[105843] = 16'b0000000000000000;
	sram_mem[105844] = 16'b0000000000000000;
	sram_mem[105845] = 16'b0000000000000000;
	sram_mem[105846] = 16'b0000000000000000;
	sram_mem[105847] = 16'b0000000000000000;
	sram_mem[105848] = 16'b0000000000000000;
	sram_mem[105849] = 16'b0000000000000000;
	sram_mem[105850] = 16'b0000000000000000;
	sram_mem[105851] = 16'b0000000000000000;
	sram_mem[105852] = 16'b0000000000000000;
	sram_mem[105853] = 16'b0000000000000000;
	sram_mem[105854] = 16'b0000000000000000;
	sram_mem[105855] = 16'b0000000000000000;
	sram_mem[105856] = 16'b0000000000000000;
	sram_mem[105857] = 16'b0000000000000000;
	sram_mem[105858] = 16'b0000000000000000;
	sram_mem[105859] = 16'b0000000000000000;
	sram_mem[105860] = 16'b0000000000000000;
	sram_mem[105861] = 16'b0000000000000000;
	sram_mem[105862] = 16'b0000000000000000;
	sram_mem[105863] = 16'b0000000000000000;
	sram_mem[105864] = 16'b0000000000000000;
	sram_mem[105865] = 16'b0000000000000000;
	sram_mem[105866] = 16'b0000000000000000;
	sram_mem[105867] = 16'b0000000000000000;
	sram_mem[105868] = 16'b0000000000000000;
	sram_mem[105869] = 16'b0000000000000000;
	sram_mem[105870] = 16'b0000000000000000;
	sram_mem[105871] = 16'b0000000000000000;
	sram_mem[105872] = 16'b0000000000000000;
	sram_mem[105873] = 16'b0000000000000000;
	sram_mem[105874] = 16'b0000000000000000;
	sram_mem[105875] = 16'b0000000000000000;
	sram_mem[105876] = 16'b0000000000000000;
	sram_mem[105877] = 16'b0000000000000000;
	sram_mem[105878] = 16'b0000000000000000;
	sram_mem[105879] = 16'b0000000000000000;
	sram_mem[105880] = 16'b0000000000000000;
	sram_mem[105881] = 16'b0000000000000000;
	sram_mem[105882] = 16'b0000000000000000;
	sram_mem[105883] = 16'b0000000000000000;
	sram_mem[105884] = 16'b0000000000000000;
	sram_mem[105885] = 16'b0000000000000000;
	sram_mem[105886] = 16'b0000000000000000;
	sram_mem[105887] = 16'b0000000000000000;
	sram_mem[105888] = 16'b0000000000000000;
	sram_mem[105889] = 16'b0000000000000000;
	sram_mem[105890] = 16'b0000000000000000;
	sram_mem[105891] = 16'b0000000000000000;
	sram_mem[105892] = 16'b0000000000000000;
	sram_mem[105893] = 16'b0000000000000000;
	sram_mem[105894] = 16'b0000000000000000;
	sram_mem[105895] = 16'b0000000000000000;
	sram_mem[105896] = 16'b0000000000000000;
	sram_mem[105897] = 16'b0000000000000000;
	sram_mem[105898] = 16'b0000000000000000;
	sram_mem[105899] = 16'b0000000000000000;
	sram_mem[105900] = 16'b0000000000000000;
	sram_mem[105901] = 16'b0000000000000000;
	sram_mem[105902] = 16'b0000000000000000;
	sram_mem[105903] = 16'b0000000000000000;
	sram_mem[105904] = 16'b0000000000000000;
	sram_mem[105905] = 16'b0000000000000000;
	sram_mem[105906] = 16'b0000000000000000;
	sram_mem[105907] = 16'b0000000000000000;
	sram_mem[105908] = 16'b0000000000000000;
	sram_mem[105909] = 16'b0000000000000000;
	sram_mem[105910] = 16'b0000000000000000;
	sram_mem[105911] = 16'b0000000000000000;
	sram_mem[105912] = 16'b0000000000000000;
	sram_mem[105913] = 16'b0000000000000000;
	sram_mem[105914] = 16'b0000000000000000;
	sram_mem[105915] = 16'b0000000000000000;
	sram_mem[105916] = 16'b0000000000000000;
	sram_mem[105917] = 16'b0000000000000000;
	sram_mem[105918] = 16'b0000000000000000;
	sram_mem[105919] = 16'b0000000000000000;
	sram_mem[105920] = 16'b0000000000000000;
	sram_mem[105921] = 16'b0000000000000000;
	sram_mem[105922] = 16'b0000000000000000;
	sram_mem[105923] = 16'b0000000000000000;
	sram_mem[105924] = 16'b0000000000000000;
	sram_mem[105925] = 16'b0000000000000000;
	sram_mem[105926] = 16'b0000000000000000;
	sram_mem[105927] = 16'b0000000000000000;
	sram_mem[105928] = 16'b0000000000000000;
	sram_mem[105929] = 16'b0000000000000000;
	sram_mem[105930] = 16'b0000000000000000;
	sram_mem[105931] = 16'b0000000000000000;
	sram_mem[105932] = 16'b0000000000000000;
	sram_mem[105933] = 16'b0000000000000000;
	sram_mem[105934] = 16'b0000000000000000;
	sram_mem[105935] = 16'b0000000000000000;
	sram_mem[105936] = 16'b0000000000000000;
	sram_mem[105937] = 16'b0000000000000000;
	sram_mem[105938] = 16'b0000000000000000;
	sram_mem[105939] = 16'b0000000000000000;
	sram_mem[105940] = 16'b0000000000000000;
	sram_mem[105941] = 16'b0000000000000000;
	sram_mem[105942] = 16'b0000000000000000;
	sram_mem[105943] = 16'b0000000000000000;
	sram_mem[105944] = 16'b0000000000000000;
	sram_mem[105945] = 16'b0000000000000000;
	sram_mem[105946] = 16'b0000000000000000;
	sram_mem[105947] = 16'b0000000000000000;
	sram_mem[105948] = 16'b0000000000000000;
	sram_mem[105949] = 16'b0000000000000000;
	sram_mem[105950] = 16'b0000000000000000;
	sram_mem[105951] = 16'b0000000000000000;
	sram_mem[105952] = 16'b0000000000000000;
	sram_mem[105953] = 16'b0000000000000000;
	sram_mem[105954] = 16'b0000000000000000;
	sram_mem[105955] = 16'b0000000000000000;
	sram_mem[105956] = 16'b0000000000000000;
	sram_mem[105957] = 16'b0000000000000000;
	sram_mem[105958] = 16'b0000000000000000;
	sram_mem[105959] = 16'b0000000000000000;
	sram_mem[105960] = 16'b0000000000000000;
	sram_mem[105961] = 16'b0000000000000000;
	sram_mem[105962] = 16'b0000000000000000;
	sram_mem[105963] = 16'b0000000000000000;
	sram_mem[105964] = 16'b0000000000000000;
	sram_mem[105965] = 16'b0000000000000000;
	sram_mem[105966] = 16'b0000000000000000;
	sram_mem[105967] = 16'b0000000000000000;
	sram_mem[105968] = 16'b0000000000000000;
	sram_mem[105969] = 16'b0000000000000000;
	sram_mem[105970] = 16'b0000000000000000;
	sram_mem[105971] = 16'b0000000000000000;
	sram_mem[105972] = 16'b0000000000000000;
	sram_mem[105973] = 16'b0000000000000000;
	sram_mem[105974] = 16'b0000000000000000;
	sram_mem[105975] = 16'b0000000000000000;
	sram_mem[105976] = 16'b0000000000000000;
	sram_mem[105977] = 16'b0000000000000000;
	sram_mem[105978] = 16'b0000000000000000;
	sram_mem[105979] = 16'b0000000000000000;
	sram_mem[105980] = 16'b0000000000000000;
	sram_mem[105981] = 16'b0000000000000000;
	sram_mem[105982] = 16'b0000000000000000;
	sram_mem[105983] = 16'b0000000000000000;
	sram_mem[105984] = 16'b0000000000000000;
	sram_mem[105985] = 16'b0000000000000000;
	sram_mem[105986] = 16'b0000000000000000;
	sram_mem[105987] = 16'b0000000000000000;
	sram_mem[105988] = 16'b0000000000000000;
	sram_mem[105989] = 16'b0000000000000000;
	sram_mem[105990] = 16'b0000000000000000;
	sram_mem[105991] = 16'b0000000000000000;
	sram_mem[105992] = 16'b0000000000000000;
	sram_mem[105993] = 16'b0000000000000000;
	sram_mem[105994] = 16'b0000000000000000;
	sram_mem[105995] = 16'b0000000000000000;
	sram_mem[105996] = 16'b0000000000000000;
	sram_mem[105997] = 16'b0000000000000000;
	sram_mem[105998] = 16'b0000000000000000;
	sram_mem[105999] = 16'b0000000000000000;
	sram_mem[106000] = 16'b0000000000000000;
	sram_mem[106001] = 16'b0000000000000000;
	sram_mem[106002] = 16'b0000000000000000;
	sram_mem[106003] = 16'b0000000000000000;
	sram_mem[106004] = 16'b0000000000000000;
	sram_mem[106005] = 16'b0000000000000000;
	sram_mem[106006] = 16'b0000000000000000;
	sram_mem[106007] = 16'b0000000000000000;
	sram_mem[106008] = 16'b0000000000000000;
	sram_mem[106009] = 16'b0000000000000000;
	sram_mem[106010] = 16'b0000000000000000;
	sram_mem[106011] = 16'b0000000000000000;
	sram_mem[106012] = 16'b0000000000000000;
	sram_mem[106013] = 16'b0000000000000000;
	sram_mem[106014] = 16'b0000000000000000;
	sram_mem[106015] = 16'b0000000000000000;
	sram_mem[106016] = 16'b0000000000000000;
	sram_mem[106017] = 16'b0000000000000000;
	sram_mem[106018] = 16'b0000000000000000;
	sram_mem[106019] = 16'b0000000000000000;
	sram_mem[106020] = 16'b0000000000000000;
	sram_mem[106021] = 16'b0000000000000000;
	sram_mem[106022] = 16'b0000000000000000;
	sram_mem[106023] = 16'b0000000000000000;
	sram_mem[106024] = 16'b0000000000000000;
	sram_mem[106025] = 16'b0000000000000000;
	sram_mem[106026] = 16'b0000000000000000;
	sram_mem[106027] = 16'b0000000000000000;
	sram_mem[106028] = 16'b0000000000000000;
	sram_mem[106029] = 16'b0000000000000000;
	sram_mem[106030] = 16'b0000000000000000;
	sram_mem[106031] = 16'b0000000000000000;
	sram_mem[106032] = 16'b0000000000000000;
	sram_mem[106033] = 16'b0000000000000000;
	sram_mem[106034] = 16'b0000000000000000;
	sram_mem[106035] = 16'b0000000000000000;
	sram_mem[106036] = 16'b0000000000000000;
	sram_mem[106037] = 16'b0000000000000000;
	sram_mem[106038] = 16'b0000000000000000;
	sram_mem[106039] = 16'b0000000000000000;
	sram_mem[106040] = 16'b0000000000000000;
	sram_mem[106041] = 16'b0000000000000000;
	sram_mem[106042] = 16'b0000000000000000;
	sram_mem[106043] = 16'b0000000000000000;
	sram_mem[106044] = 16'b0000000000000000;
	sram_mem[106045] = 16'b0000000000000000;
	sram_mem[106046] = 16'b0000000000000000;
	sram_mem[106047] = 16'b0000000000000000;
	sram_mem[106048] = 16'b0000000000000000;
	sram_mem[106049] = 16'b0000000000000000;
	sram_mem[106050] = 16'b0000000000000000;
	sram_mem[106051] = 16'b0000000000000000;
	sram_mem[106052] = 16'b0000000000000000;
	sram_mem[106053] = 16'b0000000000000000;
	sram_mem[106054] = 16'b0000000000000000;
	sram_mem[106055] = 16'b0000000000000000;
	sram_mem[106056] = 16'b0000000000000000;
	sram_mem[106057] = 16'b0000000000000000;
	sram_mem[106058] = 16'b0000000000000000;
	sram_mem[106059] = 16'b0000000000000000;
	sram_mem[106060] = 16'b0000000000000000;
	sram_mem[106061] = 16'b0000000000000000;
	sram_mem[106062] = 16'b0000000000000000;
	sram_mem[106063] = 16'b0000000000000000;
	sram_mem[106064] = 16'b0000000000000000;
	sram_mem[106065] = 16'b0000000000000000;
	sram_mem[106066] = 16'b0000000000000000;
	sram_mem[106067] = 16'b0000000000000000;
	sram_mem[106068] = 16'b0000000000000000;
	sram_mem[106069] = 16'b0000000000000000;
	sram_mem[106070] = 16'b0000000000000000;
	sram_mem[106071] = 16'b0000000000000000;
	sram_mem[106072] = 16'b0000000000000000;
	sram_mem[106073] = 16'b0000000000000000;
	sram_mem[106074] = 16'b0000000000000000;
	sram_mem[106075] = 16'b0000000000000000;
	sram_mem[106076] = 16'b0000000000000000;
	sram_mem[106077] = 16'b0000000000000000;
	sram_mem[106078] = 16'b0000000000000000;
	sram_mem[106079] = 16'b0000000000000000;
	sram_mem[106080] = 16'b0000000000000000;
	sram_mem[106081] = 16'b0000000000000000;
	sram_mem[106082] = 16'b0000000000000000;
	sram_mem[106083] = 16'b0000000000000000;
	sram_mem[106084] = 16'b0000000000000000;
	sram_mem[106085] = 16'b0000000000000000;
	sram_mem[106086] = 16'b0000000000000000;
	sram_mem[106087] = 16'b0000000000000000;
	sram_mem[106088] = 16'b0000000000000000;
	sram_mem[106089] = 16'b0000000000000000;
	sram_mem[106090] = 16'b0000000000000000;
	sram_mem[106091] = 16'b0000000000000000;
	sram_mem[106092] = 16'b0000000000000000;
	sram_mem[106093] = 16'b0000000000000000;
	sram_mem[106094] = 16'b0000000000000000;
	sram_mem[106095] = 16'b0000000000000000;
	sram_mem[106096] = 16'b0000000000000000;
	sram_mem[106097] = 16'b0000000000000000;
	sram_mem[106098] = 16'b0000000000000000;
	sram_mem[106099] = 16'b0000000000000000;
	sram_mem[106100] = 16'b0000000000000000;
	sram_mem[106101] = 16'b0000000000000000;
	sram_mem[106102] = 16'b0000000000000000;
	sram_mem[106103] = 16'b0000000000000000;
	sram_mem[106104] = 16'b0000000000000000;
	sram_mem[106105] = 16'b0000000000000000;
	sram_mem[106106] = 16'b0000000000000000;
	sram_mem[106107] = 16'b0000000000000000;
	sram_mem[106108] = 16'b0000000000000000;
	sram_mem[106109] = 16'b0000000000000000;
	sram_mem[106110] = 16'b0000000000000000;
	sram_mem[106111] = 16'b0000000000000000;
	sram_mem[106112] = 16'b0000000000000000;
	sram_mem[106113] = 16'b0000000000000000;
	sram_mem[106114] = 16'b0000000000000000;
	sram_mem[106115] = 16'b0000000000000000;
	sram_mem[106116] = 16'b0000000000000000;
	sram_mem[106117] = 16'b0000000000000000;
	sram_mem[106118] = 16'b0000000000000000;
	sram_mem[106119] = 16'b0000000000000000;
	sram_mem[106120] = 16'b0000000000000000;
	sram_mem[106121] = 16'b0000000000000000;
	sram_mem[106122] = 16'b0000000000000000;
	sram_mem[106123] = 16'b0000000000000000;
	sram_mem[106124] = 16'b0000000000000000;
	sram_mem[106125] = 16'b0000000000000000;
	sram_mem[106126] = 16'b0000000000000000;
	sram_mem[106127] = 16'b0000000000000000;
	sram_mem[106128] = 16'b0000000000000000;
	sram_mem[106129] = 16'b0000000000000000;
	sram_mem[106130] = 16'b0000000000000000;
	sram_mem[106131] = 16'b0000000000000000;
	sram_mem[106132] = 16'b0000000000000000;
	sram_mem[106133] = 16'b0000000000000000;
	sram_mem[106134] = 16'b0000000000000000;
	sram_mem[106135] = 16'b0000000000000000;
	sram_mem[106136] = 16'b0000000000000000;
	sram_mem[106137] = 16'b0000000000000000;
	sram_mem[106138] = 16'b0000000000000000;
	sram_mem[106139] = 16'b0000000000000000;
	sram_mem[106140] = 16'b0000000000000000;
	sram_mem[106141] = 16'b0000000000000000;
	sram_mem[106142] = 16'b0000000000000000;
	sram_mem[106143] = 16'b0000000000000000;
	sram_mem[106144] = 16'b0000000000000000;
	sram_mem[106145] = 16'b0000000000000000;
	sram_mem[106146] = 16'b0000000000000000;
	sram_mem[106147] = 16'b0000000000000000;
	sram_mem[106148] = 16'b0000000000000000;
	sram_mem[106149] = 16'b0000000000000000;
	sram_mem[106150] = 16'b0000000000000000;
	sram_mem[106151] = 16'b0000000000000000;
	sram_mem[106152] = 16'b0000000000000000;
	sram_mem[106153] = 16'b0000000000000000;
	sram_mem[106154] = 16'b0000000000000000;
	sram_mem[106155] = 16'b0000000000000000;
	sram_mem[106156] = 16'b0000000000000000;
	sram_mem[106157] = 16'b0000000000000000;
	sram_mem[106158] = 16'b0000000000000000;
	sram_mem[106159] = 16'b0000000000000000;
	sram_mem[106160] = 16'b0000000000000000;
	sram_mem[106161] = 16'b0000000000000000;
	sram_mem[106162] = 16'b0000000000000000;
	sram_mem[106163] = 16'b0000000000000000;
	sram_mem[106164] = 16'b0000000000000000;
	sram_mem[106165] = 16'b0000000000000000;
	sram_mem[106166] = 16'b0000000000000000;
	sram_mem[106167] = 16'b0000000000000000;
	sram_mem[106168] = 16'b0000000000000000;
	sram_mem[106169] = 16'b0000000000000000;
	sram_mem[106170] = 16'b0000000000000000;
	sram_mem[106171] = 16'b0000000000000000;
	sram_mem[106172] = 16'b0000000000000000;
	sram_mem[106173] = 16'b0000000000000000;
	sram_mem[106174] = 16'b0000000000000000;
	sram_mem[106175] = 16'b0000000000000000;
	sram_mem[106176] = 16'b0000000000000000;
	sram_mem[106177] = 16'b0000000000000000;
	sram_mem[106178] = 16'b0000000000000000;
	sram_mem[106179] = 16'b0000000000000000;
	sram_mem[106180] = 16'b0000000000000000;
	sram_mem[106181] = 16'b0000000000000000;
	sram_mem[106182] = 16'b0000000000000000;
	sram_mem[106183] = 16'b0000000000000000;
	sram_mem[106184] = 16'b0000000000000000;
	sram_mem[106185] = 16'b0000000000000000;
	sram_mem[106186] = 16'b0000000000000000;
	sram_mem[106187] = 16'b0000000000000000;
	sram_mem[106188] = 16'b0000000000000000;
	sram_mem[106189] = 16'b0000000000000000;
	sram_mem[106190] = 16'b0000000000000000;
	sram_mem[106191] = 16'b0000000000000000;
	sram_mem[106192] = 16'b0000000000000000;
	sram_mem[106193] = 16'b0000000000000000;
	sram_mem[106194] = 16'b0000000000000000;
	sram_mem[106195] = 16'b0000000000000000;
	sram_mem[106196] = 16'b0000000000000000;
	sram_mem[106197] = 16'b0000000000000000;
	sram_mem[106198] = 16'b0000000000000000;
	sram_mem[106199] = 16'b0000000000000000;
	sram_mem[106200] = 16'b0000000000000000;
	sram_mem[106201] = 16'b0000000000000000;
	sram_mem[106202] = 16'b0000000000000000;
	sram_mem[106203] = 16'b0000000000000000;
	sram_mem[106204] = 16'b0000000000000000;
	sram_mem[106205] = 16'b0000000000000000;
	sram_mem[106206] = 16'b0000000000000000;
	sram_mem[106207] = 16'b0000000000000000;
	sram_mem[106208] = 16'b0000000000000000;
	sram_mem[106209] = 16'b0000000000000000;
	sram_mem[106210] = 16'b0000000000000000;
	sram_mem[106211] = 16'b0000000000000000;
	sram_mem[106212] = 16'b0000000000000000;
	sram_mem[106213] = 16'b0000000000000000;
	sram_mem[106214] = 16'b0000000000000000;
	sram_mem[106215] = 16'b0000000000000000;
	sram_mem[106216] = 16'b0000000000000000;
	sram_mem[106217] = 16'b0000000000000000;
	sram_mem[106218] = 16'b0000000000000000;
	sram_mem[106219] = 16'b0000000000000000;
	sram_mem[106220] = 16'b0000000000000000;
	sram_mem[106221] = 16'b0000000000000000;
	sram_mem[106222] = 16'b0000000000000000;
	sram_mem[106223] = 16'b0000000000000000;
	sram_mem[106224] = 16'b0000000000000000;
	sram_mem[106225] = 16'b0000000000000000;
	sram_mem[106226] = 16'b0000000000000000;
	sram_mem[106227] = 16'b0000000000000000;
	sram_mem[106228] = 16'b0000000000000000;
	sram_mem[106229] = 16'b0000000000000000;
	sram_mem[106230] = 16'b0000000000000000;
	sram_mem[106231] = 16'b0000000000000000;
	sram_mem[106232] = 16'b0000000000000000;
	sram_mem[106233] = 16'b0000000000000000;
	sram_mem[106234] = 16'b0000000000000000;
	sram_mem[106235] = 16'b0000000000000000;
	sram_mem[106236] = 16'b0000000000000000;
	sram_mem[106237] = 16'b0000000000000000;
	sram_mem[106238] = 16'b0000000000000000;
	sram_mem[106239] = 16'b0000000000000000;
	sram_mem[106240] = 16'b0000000000000000;
	sram_mem[106241] = 16'b0000000000000000;
	sram_mem[106242] = 16'b0000000000000000;
	sram_mem[106243] = 16'b0000000000000000;
	sram_mem[106244] = 16'b0000000000000000;
	sram_mem[106245] = 16'b0000000000000000;
	sram_mem[106246] = 16'b0000000000000000;
	sram_mem[106247] = 16'b0000000000000000;
	sram_mem[106248] = 16'b0000000000000000;
	sram_mem[106249] = 16'b0000000000000000;
	sram_mem[106250] = 16'b0000000000000000;
	sram_mem[106251] = 16'b0000000000000000;
	sram_mem[106252] = 16'b0000000000000000;
	sram_mem[106253] = 16'b0000000000000000;
	sram_mem[106254] = 16'b0000000000000000;
	sram_mem[106255] = 16'b0000000000000000;
	sram_mem[106256] = 16'b0000000000000000;
	sram_mem[106257] = 16'b0000000000000000;
	sram_mem[106258] = 16'b0000000000000000;
	sram_mem[106259] = 16'b0000000000000000;
	sram_mem[106260] = 16'b0000000000000000;
	sram_mem[106261] = 16'b0000000000000000;
	sram_mem[106262] = 16'b0000000000000000;
	sram_mem[106263] = 16'b0000000000000000;
	sram_mem[106264] = 16'b0000000000000000;
	sram_mem[106265] = 16'b0000000000000000;
	sram_mem[106266] = 16'b0000000000000000;
	sram_mem[106267] = 16'b0000000000000000;
	sram_mem[106268] = 16'b0000000000000000;
	sram_mem[106269] = 16'b0000000000000000;
	sram_mem[106270] = 16'b0000000000000000;
	sram_mem[106271] = 16'b0000000000000000;
	sram_mem[106272] = 16'b0000000000000000;
	sram_mem[106273] = 16'b0000000000000000;
	sram_mem[106274] = 16'b0000000000000000;
	sram_mem[106275] = 16'b0000000000000000;
	sram_mem[106276] = 16'b0000000000000000;
	sram_mem[106277] = 16'b0000000000000000;
	sram_mem[106278] = 16'b0000000000000000;
	sram_mem[106279] = 16'b0000000000000000;
	sram_mem[106280] = 16'b0000000000000000;
	sram_mem[106281] = 16'b0000000000000000;
	sram_mem[106282] = 16'b0000000000000000;
	sram_mem[106283] = 16'b0000000000000000;
	sram_mem[106284] = 16'b0000000000000000;
	sram_mem[106285] = 16'b0000000000000000;
	sram_mem[106286] = 16'b0000000000000000;
	sram_mem[106287] = 16'b0000000000000000;
	sram_mem[106288] = 16'b0000000000000000;
	sram_mem[106289] = 16'b0000000000000000;
	sram_mem[106290] = 16'b0000000000000000;
	sram_mem[106291] = 16'b0000000000000000;
	sram_mem[106292] = 16'b0000000000000000;
	sram_mem[106293] = 16'b0000000000000000;
	sram_mem[106294] = 16'b0000000000000000;
	sram_mem[106295] = 16'b0000000000000000;
	sram_mem[106296] = 16'b0000000000000000;
	sram_mem[106297] = 16'b0000000000000000;
	sram_mem[106298] = 16'b0000000000000000;
	sram_mem[106299] = 16'b0000000000000000;
	sram_mem[106300] = 16'b0000000000000000;
	sram_mem[106301] = 16'b0000000000000000;
	sram_mem[106302] = 16'b0000000000000000;
	sram_mem[106303] = 16'b0000000000000000;
	sram_mem[106304] = 16'b0000000000000000;
	sram_mem[106305] = 16'b0000000000000000;
	sram_mem[106306] = 16'b0000000000000000;
	sram_mem[106307] = 16'b0000000000000000;
	sram_mem[106308] = 16'b0000000000000000;
	sram_mem[106309] = 16'b0000000000000000;
	sram_mem[106310] = 16'b0000000000000000;
	sram_mem[106311] = 16'b0000000000000000;
	sram_mem[106312] = 16'b0000000000000000;
	sram_mem[106313] = 16'b0000000000000000;
	sram_mem[106314] = 16'b0000000000000000;
	sram_mem[106315] = 16'b0000000000000000;
	sram_mem[106316] = 16'b0000000000000000;
	sram_mem[106317] = 16'b0000000000000000;
	sram_mem[106318] = 16'b0000000000000000;
	sram_mem[106319] = 16'b0000000000000000;
	sram_mem[106320] = 16'b0000000000000000;
	sram_mem[106321] = 16'b0000000000000000;
	sram_mem[106322] = 16'b0000000000000000;
	sram_mem[106323] = 16'b0000000000000000;
	sram_mem[106324] = 16'b0000000000000000;
	sram_mem[106325] = 16'b0000000000000000;
	sram_mem[106326] = 16'b0000000000000000;
	sram_mem[106327] = 16'b0000000000000000;
	sram_mem[106328] = 16'b0000000000000000;
	sram_mem[106329] = 16'b0000000000000000;
	sram_mem[106330] = 16'b0000000000000000;
	sram_mem[106331] = 16'b0000000000000000;
	sram_mem[106332] = 16'b0000000000000000;
	sram_mem[106333] = 16'b0000000000000000;
	sram_mem[106334] = 16'b0000000000000000;
	sram_mem[106335] = 16'b0000000000000000;
	sram_mem[106336] = 16'b0000000000000000;
	sram_mem[106337] = 16'b0000000000000000;
	sram_mem[106338] = 16'b0000000000000000;
	sram_mem[106339] = 16'b0000000000000000;
	sram_mem[106340] = 16'b0000000000000000;
	sram_mem[106341] = 16'b0000000000000000;
	sram_mem[106342] = 16'b0000000000000000;
	sram_mem[106343] = 16'b0000000000000000;
	sram_mem[106344] = 16'b0000000000000000;
	sram_mem[106345] = 16'b0000000000000000;
	sram_mem[106346] = 16'b0000000000000000;
	sram_mem[106347] = 16'b0000000000000000;
	sram_mem[106348] = 16'b0000000000000000;
	sram_mem[106349] = 16'b0000000000000000;
	sram_mem[106350] = 16'b0000000000000000;
	sram_mem[106351] = 16'b0000000000000000;
	sram_mem[106352] = 16'b0000000000000000;
	sram_mem[106353] = 16'b0000000000000000;
	sram_mem[106354] = 16'b0000000000000000;
	sram_mem[106355] = 16'b0000000000000000;
	sram_mem[106356] = 16'b0000000000000000;
	sram_mem[106357] = 16'b0000000000000000;
	sram_mem[106358] = 16'b0000000000000000;
	sram_mem[106359] = 16'b0000000000000000;
	sram_mem[106360] = 16'b0000000000000000;
	sram_mem[106361] = 16'b0000000000000000;
	sram_mem[106362] = 16'b0000000000000000;
	sram_mem[106363] = 16'b0000000000000000;
	sram_mem[106364] = 16'b0000000000000000;
	sram_mem[106365] = 16'b0000000000000000;
	sram_mem[106366] = 16'b0000000000000000;
	sram_mem[106367] = 16'b0000000000000000;
	sram_mem[106368] = 16'b0000000000000000;
	sram_mem[106369] = 16'b0000000000000000;
	sram_mem[106370] = 16'b0000000000000000;
	sram_mem[106371] = 16'b0000000000000000;
	sram_mem[106372] = 16'b0000000000000000;
	sram_mem[106373] = 16'b0000000000000000;
	sram_mem[106374] = 16'b0000000000000000;
	sram_mem[106375] = 16'b0000000000000000;
	sram_mem[106376] = 16'b0000000000000000;
	sram_mem[106377] = 16'b0000000000000000;
	sram_mem[106378] = 16'b0000000000000000;
	sram_mem[106379] = 16'b0000000000000000;
	sram_mem[106380] = 16'b0000000000000000;
	sram_mem[106381] = 16'b0000000000000000;
	sram_mem[106382] = 16'b0000000000000000;
	sram_mem[106383] = 16'b0000000000000000;
	sram_mem[106384] = 16'b0000000000000000;
	sram_mem[106385] = 16'b0000000000000000;
	sram_mem[106386] = 16'b0000000000000000;
	sram_mem[106387] = 16'b0000000000000000;
	sram_mem[106388] = 16'b0000000000000000;
	sram_mem[106389] = 16'b0000000000000000;
	sram_mem[106390] = 16'b0000000000000000;
	sram_mem[106391] = 16'b0000000000000000;
	sram_mem[106392] = 16'b0000000000000000;
	sram_mem[106393] = 16'b0000000000000000;
	sram_mem[106394] = 16'b0000000000000000;
	sram_mem[106395] = 16'b0000000000000000;
	sram_mem[106396] = 16'b0000000000000000;
	sram_mem[106397] = 16'b0000000000000000;
	sram_mem[106398] = 16'b0000000000000000;
	sram_mem[106399] = 16'b0000000000000000;
	sram_mem[106400] = 16'b0000000000000000;
	sram_mem[106401] = 16'b0000000000000000;
	sram_mem[106402] = 16'b0000000000000000;
	sram_mem[106403] = 16'b0000000000000000;
	sram_mem[106404] = 16'b0000000000000000;
	sram_mem[106405] = 16'b0000000000000000;
	sram_mem[106406] = 16'b0000000000000000;
	sram_mem[106407] = 16'b0000000000000000;
	sram_mem[106408] = 16'b0000000000000000;
	sram_mem[106409] = 16'b0000000000000000;
	sram_mem[106410] = 16'b0000000000000000;
	sram_mem[106411] = 16'b0000000000000000;
	sram_mem[106412] = 16'b0000000000000000;
	sram_mem[106413] = 16'b0000000000000000;
	sram_mem[106414] = 16'b0000000000000000;
	sram_mem[106415] = 16'b0000000000000000;
	sram_mem[106416] = 16'b0000000000000000;
	sram_mem[106417] = 16'b0000000000000000;
	sram_mem[106418] = 16'b0000000000000000;
	sram_mem[106419] = 16'b0000000000000000;
	sram_mem[106420] = 16'b0000000000000000;
	sram_mem[106421] = 16'b0000000000000000;
	sram_mem[106422] = 16'b0000000000000000;
	sram_mem[106423] = 16'b0000000000000000;
	sram_mem[106424] = 16'b0000000000000000;
	sram_mem[106425] = 16'b0000000000000000;
	sram_mem[106426] = 16'b0000000000000000;
	sram_mem[106427] = 16'b0000000000000000;
	sram_mem[106428] = 16'b0000000000000000;
	sram_mem[106429] = 16'b0000000000000000;
	sram_mem[106430] = 16'b0000000000000000;
	sram_mem[106431] = 16'b0000000000000000;
	sram_mem[106432] = 16'b0000000000000000;
	sram_mem[106433] = 16'b0000000000000000;
	sram_mem[106434] = 16'b0000000000000000;
	sram_mem[106435] = 16'b0000000000000000;
	sram_mem[106436] = 16'b0000000000000000;
	sram_mem[106437] = 16'b0000000000000000;
	sram_mem[106438] = 16'b0000000000000000;
	sram_mem[106439] = 16'b0000000000000000;
	sram_mem[106440] = 16'b0000000000000000;
	sram_mem[106441] = 16'b0000000000000000;
	sram_mem[106442] = 16'b0000000000000000;
	sram_mem[106443] = 16'b0000000000000000;
	sram_mem[106444] = 16'b0000000000000000;
	sram_mem[106445] = 16'b0000000000000000;
	sram_mem[106446] = 16'b0000000000000000;
	sram_mem[106447] = 16'b0000000000000000;
	sram_mem[106448] = 16'b0000000000000000;
	sram_mem[106449] = 16'b0000000000000000;
	sram_mem[106450] = 16'b0000000000000000;
	sram_mem[106451] = 16'b0000000000000000;
	sram_mem[106452] = 16'b0000000000000000;
	sram_mem[106453] = 16'b0000000000000000;
	sram_mem[106454] = 16'b0000000000000000;
	sram_mem[106455] = 16'b0000000000000000;
	sram_mem[106456] = 16'b0000000000000000;
	sram_mem[106457] = 16'b0000000000000000;
	sram_mem[106458] = 16'b0000000000000000;
	sram_mem[106459] = 16'b0000000000000000;
	sram_mem[106460] = 16'b0000000000000000;
	sram_mem[106461] = 16'b0000000000000000;
	sram_mem[106462] = 16'b0000000000000000;
	sram_mem[106463] = 16'b0000000000000000;
	sram_mem[106464] = 16'b0000000000000000;
	sram_mem[106465] = 16'b0000000000000000;
	sram_mem[106466] = 16'b0000000000000000;
	sram_mem[106467] = 16'b0000000000000000;
	sram_mem[106468] = 16'b0000000000000000;
	sram_mem[106469] = 16'b0000000000000000;
	sram_mem[106470] = 16'b0000000000000000;
	sram_mem[106471] = 16'b0000000000000000;
	sram_mem[106472] = 16'b0000000000000000;
	sram_mem[106473] = 16'b0000000000000000;
	sram_mem[106474] = 16'b0000000000000000;
	sram_mem[106475] = 16'b0000000000000000;
	sram_mem[106476] = 16'b0000000000000000;
	sram_mem[106477] = 16'b0000000000000000;
	sram_mem[106478] = 16'b0000000000000000;
	sram_mem[106479] = 16'b0000000000000000;
	sram_mem[106480] = 16'b0000000000000000;
	sram_mem[106481] = 16'b0000000000000000;
	sram_mem[106482] = 16'b0000000000000000;
	sram_mem[106483] = 16'b0000000000000000;
	sram_mem[106484] = 16'b0000000000000000;
	sram_mem[106485] = 16'b0000000000000000;
	sram_mem[106486] = 16'b0000000000000000;
	sram_mem[106487] = 16'b0000000000000000;
	sram_mem[106488] = 16'b0000000000000000;
	sram_mem[106489] = 16'b0000000000000000;
	sram_mem[106490] = 16'b0000000000000000;
	sram_mem[106491] = 16'b0000000000000000;
	sram_mem[106492] = 16'b0000000000000000;
	sram_mem[106493] = 16'b0000000000000000;
	sram_mem[106494] = 16'b0000000000000000;
	sram_mem[106495] = 16'b0000000000000000;
	sram_mem[106496] = 16'b0000000000000000;
	sram_mem[106497] = 16'b0000000000000000;
	sram_mem[106498] = 16'b0000000000000000;
	sram_mem[106499] = 16'b0000000000000000;
	sram_mem[106500] = 16'b0000000000000000;
	sram_mem[106501] = 16'b0000000000000000;
	sram_mem[106502] = 16'b0000000000000000;
	sram_mem[106503] = 16'b0000000000000000;
	sram_mem[106504] = 16'b0000000000000000;
	sram_mem[106505] = 16'b0000000000000000;
	sram_mem[106506] = 16'b0000000000000000;
	sram_mem[106507] = 16'b0000000000000000;
	sram_mem[106508] = 16'b0000000000000000;
	sram_mem[106509] = 16'b0000000000000000;
	sram_mem[106510] = 16'b0000000000000000;
	sram_mem[106511] = 16'b0000000000000000;
	sram_mem[106512] = 16'b0000000000000000;
	sram_mem[106513] = 16'b0000000000000000;
	sram_mem[106514] = 16'b0000000000000000;
	sram_mem[106515] = 16'b0000000000000000;
	sram_mem[106516] = 16'b0000000000000000;
	sram_mem[106517] = 16'b0000000000000000;
	sram_mem[106518] = 16'b0000000000000000;
	sram_mem[106519] = 16'b0000000000000000;
	sram_mem[106520] = 16'b0000000000000000;
	sram_mem[106521] = 16'b0000000000000000;
	sram_mem[106522] = 16'b0000000000000000;
	sram_mem[106523] = 16'b0000000000000000;
	sram_mem[106524] = 16'b0000000000000000;
	sram_mem[106525] = 16'b0000000000000000;
	sram_mem[106526] = 16'b0000000000000000;
	sram_mem[106527] = 16'b0000000000000000;
	sram_mem[106528] = 16'b0000000000000000;
	sram_mem[106529] = 16'b0000000000000000;
	sram_mem[106530] = 16'b0000000000000000;
	sram_mem[106531] = 16'b0000000000000000;
	sram_mem[106532] = 16'b0000000000000000;
	sram_mem[106533] = 16'b0000000000000000;
	sram_mem[106534] = 16'b0000000000000000;
	sram_mem[106535] = 16'b0000000000000000;
	sram_mem[106536] = 16'b0000000000000000;
	sram_mem[106537] = 16'b0000000000000000;
	sram_mem[106538] = 16'b0000000000000000;
	sram_mem[106539] = 16'b0000000000000000;
	sram_mem[106540] = 16'b0000000000000000;
	sram_mem[106541] = 16'b0000000000000000;
	sram_mem[106542] = 16'b0000000000000000;
	sram_mem[106543] = 16'b0000000000000000;
	sram_mem[106544] = 16'b0000000000000000;
	sram_mem[106545] = 16'b0000000000000000;
	sram_mem[106546] = 16'b0000000000000000;
	sram_mem[106547] = 16'b0000000000000000;
	sram_mem[106548] = 16'b0000000000000000;
	sram_mem[106549] = 16'b0000000000000000;
	sram_mem[106550] = 16'b0000000000000000;
	sram_mem[106551] = 16'b0000000000000000;
	sram_mem[106552] = 16'b0000000000000000;
	sram_mem[106553] = 16'b0000000000000000;
	sram_mem[106554] = 16'b0000000000000000;
	sram_mem[106555] = 16'b0000000000000000;
	sram_mem[106556] = 16'b0000000000000000;
	sram_mem[106557] = 16'b0000000000000000;
	sram_mem[106558] = 16'b0000000000000000;
	sram_mem[106559] = 16'b0000000000000000;
	sram_mem[106560] = 16'b0000000000000000;
	sram_mem[106561] = 16'b0000000000000000;
	sram_mem[106562] = 16'b0000000000000000;
	sram_mem[106563] = 16'b0000000000000000;
	sram_mem[106564] = 16'b0000000000000000;
	sram_mem[106565] = 16'b0000000000000000;
	sram_mem[106566] = 16'b0000000000000000;
	sram_mem[106567] = 16'b0000000000000000;
	sram_mem[106568] = 16'b0000000000000000;
	sram_mem[106569] = 16'b0000000000000000;
	sram_mem[106570] = 16'b0000000000000000;
	sram_mem[106571] = 16'b0000000000000000;
	sram_mem[106572] = 16'b0000000000000000;
	sram_mem[106573] = 16'b0000000000000000;
	sram_mem[106574] = 16'b0000000000000000;
	sram_mem[106575] = 16'b0000000000000000;
	sram_mem[106576] = 16'b0000000000000000;
	sram_mem[106577] = 16'b0000000000000000;
	sram_mem[106578] = 16'b0000000000000000;
	sram_mem[106579] = 16'b0000000000000000;
	sram_mem[106580] = 16'b0000000000000000;
	sram_mem[106581] = 16'b0000000000000000;
	sram_mem[106582] = 16'b0000000000000000;
	sram_mem[106583] = 16'b0000000000000000;
	sram_mem[106584] = 16'b0000000000000000;
	sram_mem[106585] = 16'b0000000000000000;
	sram_mem[106586] = 16'b0000000000000000;
	sram_mem[106587] = 16'b0000000000000000;
	sram_mem[106588] = 16'b0000000000000000;
	sram_mem[106589] = 16'b0000000000000000;
	sram_mem[106590] = 16'b0000000000000000;
	sram_mem[106591] = 16'b0000000000000000;
	sram_mem[106592] = 16'b0000000000000000;
	sram_mem[106593] = 16'b0000000000000000;
	sram_mem[106594] = 16'b0000000000000000;
	sram_mem[106595] = 16'b0000000000000000;
	sram_mem[106596] = 16'b0000000000000000;
	sram_mem[106597] = 16'b0000000000000000;
	sram_mem[106598] = 16'b0000000000000000;
	sram_mem[106599] = 16'b0000000000000000;
	sram_mem[106600] = 16'b0000000000000000;
	sram_mem[106601] = 16'b0000000000000000;
	sram_mem[106602] = 16'b0000000000000000;
	sram_mem[106603] = 16'b0000000000000000;
	sram_mem[106604] = 16'b0000000000000000;
	sram_mem[106605] = 16'b0000000000000000;
	sram_mem[106606] = 16'b0000000000000000;
	sram_mem[106607] = 16'b0000000000000000;
	sram_mem[106608] = 16'b0000000000000000;
	sram_mem[106609] = 16'b0000000000000000;
	sram_mem[106610] = 16'b0000000000000000;
	sram_mem[106611] = 16'b0000000000000000;
	sram_mem[106612] = 16'b0000000000000000;
	sram_mem[106613] = 16'b0000000000000000;
	sram_mem[106614] = 16'b0000000000000000;
	sram_mem[106615] = 16'b0000000000000000;
	sram_mem[106616] = 16'b0000000000000000;
	sram_mem[106617] = 16'b0000000000000000;
	sram_mem[106618] = 16'b0000000000000000;
	sram_mem[106619] = 16'b0000000000000000;
	sram_mem[106620] = 16'b0000000000000000;
	sram_mem[106621] = 16'b0000000000000000;
	sram_mem[106622] = 16'b0000000000000000;
	sram_mem[106623] = 16'b0000000000000000;
	sram_mem[106624] = 16'b0000000000000000;
	sram_mem[106625] = 16'b0000000000000000;
	sram_mem[106626] = 16'b0000000000000000;
	sram_mem[106627] = 16'b0000000000000000;
	sram_mem[106628] = 16'b0000000000000000;
	sram_mem[106629] = 16'b0000000000000000;
	sram_mem[106630] = 16'b0000000000000000;
	sram_mem[106631] = 16'b0000000000000000;
	sram_mem[106632] = 16'b0000000000000000;
	sram_mem[106633] = 16'b0000000000000000;
	sram_mem[106634] = 16'b0000000000000000;
	sram_mem[106635] = 16'b0000000000000000;
	sram_mem[106636] = 16'b0000000000000000;
	sram_mem[106637] = 16'b0000000000000000;
	sram_mem[106638] = 16'b0000000000000000;
	sram_mem[106639] = 16'b0000000000000000;
	sram_mem[106640] = 16'b0000000000000000;
	sram_mem[106641] = 16'b0000000000000000;
	sram_mem[106642] = 16'b0000000000000000;
	sram_mem[106643] = 16'b0000000000000000;
	sram_mem[106644] = 16'b0000000000000000;
	sram_mem[106645] = 16'b0000000000000000;
	sram_mem[106646] = 16'b0000000000000000;
	sram_mem[106647] = 16'b0000000000000000;
	sram_mem[106648] = 16'b0000000000000000;
	sram_mem[106649] = 16'b0000000000000000;
	sram_mem[106650] = 16'b0000000000000000;
	sram_mem[106651] = 16'b0000000000000000;
	sram_mem[106652] = 16'b0000000000000000;
	sram_mem[106653] = 16'b0000000000000000;
	sram_mem[106654] = 16'b0000000000000000;
	sram_mem[106655] = 16'b0000000000000000;
	sram_mem[106656] = 16'b0000000000000000;
	sram_mem[106657] = 16'b0000000000000000;
	sram_mem[106658] = 16'b0000000000000000;
	sram_mem[106659] = 16'b0000000000000000;
	sram_mem[106660] = 16'b0000000000000000;
	sram_mem[106661] = 16'b0000000000000000;
	sram_mem[106662] = 16'b0000000000000000;
	sram_mem[106663] = 16'b0000000000000000;
	sram_mem[106664] = 16'b0000000000000000;
	sram_mem[106665] = 16'b0000000000000000;
	sram_mem[106666] = 16'b0000000000000000;
	sram_mem[106667] = 16'b0000000000000000;
	sram_mem[106668] = 16'b0000000000000000;
	sram_mem[106669] = 16'b0000000000000000;
	sram_mem[106670] = 16'b0000000000000000;
	sram_mem[106671] = 16'b0000000000000000;
	sram_mem[106672] = 16'b0000000000000000;
	sram_mem[106673] = 16'b0000000000000000;
	sram_mem[106674] = 16'b0000000000000000;
	sram_mem[106675] = 16'b0000000000000000;
	sram_mem[106676] = 16'b0000000000000000;
	sram_mem[106677] = 16'b0000000000000000;
	sram_mem[106678] = 16'b0000000000000000;
	sram_mem[106679] = 16'b0000000000000000;
	sram_mem[106680] = 16'b0000000000000000;
	sram_mem[106681] = 16'b0000000000000000;
	sram_mem[106682] = 16'b0000000000000000;
	sram_mem[106683] = 16'b0000000000000000;
	sram_mem[106684] = 16'b0000000000000000;
	sram_mem[106685] = 16'b0000000000000000;
	sram_mem[106686] = 16'b0000000000000000;
	sram_mem[106687] = 16'b0000000000000000;
	sram_mem[106688] = 16'b0000000000000000;
	sram_mem[106689] = 16'b0000000000000000;
	sram_mem[106690] = 16'b0000000000000000;
	sram_mem[106691] = 16'b0000000000000000;
	sram_mem[106692] = 16'b0000000000000000;
	sram_mem[106693] = 16'b0000000000000000;
	sram_mem[106694] = 16'b0000000000000000;
	sram_mem[106695] = 16'b0000000000000000;
	sram_mem[106696] = 16'b0000000000000000;
	sram_mem[106697] = 16'b0000000000000000;
	sram_mem[106698] = 16'b0000000000000000;
	sram_mem[106699] = 16'b0000000000000000;
	sram_mem[106700] = 16'b0000000000000000;
	sram_mem[106701] = 16'b0000000000000000;
	sram_mem[106702] = 16'b0000000000000000;
	sram_mem[106703] = 16'b0000000000000000;
	sram_mem[106704] = 16'b0000000000000000;
	sram_mem[106705] = 16'b0000000000000000;
	sram_mem[106706] = 16'b0000000000000000;
	sram_mem[106707] = 16'b0000000000000000;
	sram_mem[106708] = 16'b0000000000000000;
	sram_mem[106709] = 16'b0000000000000000;
	sram_mem[106710] = 16'b0000000000000000;
	sram_mem[106711] = 16'b0000000000000000;
	sram_mem[106712] = 16'b0000000000000000;
	sram_mem[106713] = 16'b0000000000000000;
	sram_mem[106714] = 16'b0000000000000000;
	sram_mem[106715] = 16'b0000000000000000;
	sram_mem[106716] = 16'b0000000000000000;
	sram_mem[106717] = 16'b0000000000000000;
	sram_mem[106718] = 16'b0000000000000000;
	sram_mem[106719] = 16'b0000000000000000;
	sram_mem[106720] = 16'b0000000000000000;
	sram_mem[106721] = 16'b0000000000000000;
	sram_mem[106722] = 16'b0000000000000000;
	sram_mem[106723] = 16'b0000000000000000;
	sram_mem[106724] = 16'b0000000000000000;
	sram_mem[106725] = 16'b0000000000000000;
	sram_mem[106726] = 16'b0000000000000000;
	sram_mem[106727] = 16'b0000000000000000;
	sram_mem[106728] = 16'b0000000000000000;
	sram_mem[106729] = 16'b0000000000000000;
	sram_mem[106730] = 16'b0000000000000000;
	sram_mem[106731] = 16'b0000000000000000;
	sram_mem[106732] = 16'b0000000000000000;
	sram_mem[106733] = 16'b0000000000000000;
	sram_mem[106734] = 16'b0000000000000000;
	sram_mem[106735] = 16'b0000000000000000;
	sram_mem[106736] = 16'b0000000000000000;
	sram_mem[106737] = 16'b0000000000000000;
	sram_mem[106738] = 16'b0000000000000000;
	sram_mem[106739] = 16'b0000000000000000;
	sram_mem[106740] = 16'b0000000000000000;
	sram_mem[106741] = 16'b0000000000000000;
	sram_mem[106742] = 16'b0000000000000000;
	sram_mem[106743] = 16'b0000000000000000;
	sram_mem[106744] = 16'b0000000000000000;
	sram_mem[106745] = 16'b0000000000000000;
	sram_mem[106746] = 16'b0000000000000000;
	sram_mem[106747] = 16'b0000000000000000;
	sram_mem[106748] = 16'b0000000000000000;
	sram_mem[106749] = 16'b0000000000000000;
	sram_mem[106750] = 16'b0000000000000000;
	sram_mem[106751] = 16'b0000000000000000;
	sram_mem[106752] = 16'b0000000000000000;
	sram_mem[106753] = 16'b0000000000000000;
	sram_mem[106754] = 16'b0000000000000000;
	sram_mem[106755] = 16'b0000000000000000;
	sram_mem[106756] = 16'b0000000000000000;
	sram_mem[106757] = 16'b0000000000000000;
	sram_mem[106758] = 16'b0000000000000000;
	sram_mem[106759] = 16'b0000000000000000;
	sram_mem[106760] = 16'b0000000000000000;
	sram_mem[106761] = 16'b0000000000000000;
	sram_mem[106762] = 16'b0000000000000000;
	sram_mem[106763] = 16'b0000000000000000;
	sram_mem[106764] = 16'b0000000000000000;
	sram_mem[106765] = 16'b0000000000000000;
	sram_mem[106766] = 16'b0000000000000000;
	sram_mem[106767] = 16'b0000000000000000;
	sram_mem[106768] = 16'b0000000000000000;
	sram_mem[106769] = 16'b0000000000000000;
	sram_mem[106770] = 16'b0000000000000000;
	sram_mem[106771] = 16'b0000000000000000;
	sram_mem[106772] = 16'b0000000000000000;
	sram_mem[106773] = 16'b0000000000000000;
	sram_mem[106774] = 16'b0000000000000000;
	sram_mem[106775] = 16'b0000000000000000;
	sram_mem[106776] = 16'b0000000000000000;
	sram_mem[106777] = 16'b0000000000000000;
	sram_mem[106778] = 16'b0000000000000000;
	sram_mem[106779] = 16'b0000000000000000;
	sram_mem[106780] = 16'b0000000000000000;
	sram_mem[106781] = 16'b0000000000000000;
	sram_mem[106782] = 16'b0000000000000000;
	sram_mem[106783] = 16'b0000000000000000;
	sram_mem[106784] = 16'b0000000000000000;
	sram_mem[106785] = 16'b0000000000000000;
	sram_mem[106786] = 16'b0000000000000000;
	sram_mem[106787] = 16'b0000000000000000;
	sram_mem[106788] = 16'b0000000000000000;
	sram_mem[106789] = 16'b0000000000000000;
	sram_mem[106790] = 16'b0000000000000000;
	sram_mem[106791] = 16'b0000000000000000;
	sram_mem[106792] = 16'b0000000000000000;
	sram_mem[106793] = 16'b0000000000000000;
	sram_mem[106794] = 16'b0000000000000000;
	sram_mem[106795] = 16'b0000000000000000;
	sram_mem[106796] = 16'b0000000000000000;
	sram_mem[106797] = 16'b0000000000000000;
	sram_mem[106798] = 16'b0000000000000000;
	sram_mem[106799] = 16'b0000000000000000;
	sram_mem[106800] = 16'b0000000000000000;
	sram_mem[106801] = 16'b0000000000000000;
	sram_mem[106802] = 16'b0000000000000000;
	sram_mem[106803] = 16'b0000000000000000;
	sram_mem[106804] = 16'b0000000000000000;
	sram_mem[106805] = 16'b0000000000000000;
	sram_mem[106806] = 16'b0000000000000000;
	sram_mem[106807] = 16'b0000000000000000;
	sram_mem[106808] = 16'b0000000000000000;
	sram_mem[106809] = 16'b0000000000000000;
	sram_mem[106810] = 16'b0000000000000000;
	sram_mem[106811] = 16'b0000000000000000;
	sram_mem[106812] = 16'b0000000000000000;
	sram_mem[106813] = 16'b0000000000000000;
	sram_mem[106814] = 16'b0000000000000000;
	sram_mem[106815] = 16'b0000000000000000;
	sram_mem[106816] = 16'b0000000000000000;
	sram_mem[106817] = 16'b0000000000000000;
	sram_mem[106818] = 16'b0000000000000000;
	sram_mem[106819] = 16'b0000000000000000;
	sram_mem[106820] = 16'b0000000000000000;
	sram_mem[106821] = 16'b0000000000000000;
	sram_mem[106822] = 16'b0000000000000000;
	sram_mem[106823] = 16'b0000000000000000;
	sram_mem[106824] = 16'b0000000000000000;
	sram_mem[106825] = 16'b0000000000000000;
	sram_mem[106826] = 16'b0000000000000000;
	sram_mem[106827] = 16'b0000000000000000;
	sram_mem[106828] = 16'b0000000000000000;
	sram_mem[106829] = 16'b0000000000000000;
	sram_mem[106830] = 16'b0000000000000000;
	sram_mem[106831] = 16'b0000000000000000;
	sram_mem[106832] = 16'b0000000000000000;
	sram_mem[106833] = 16'b0000000000000000;
	sram_mem[106834] = 16'b0000000000000000;
	sram_mem[106835] = 16'b0000000000000000;
	sram_mem[106836] = 16'b0000000000000000;
	sram_mem[106837] = 16'b0000000000000000;
	sram_mem[106838] = 16'b0000000000000000;
	sram_mem[106839] = 16'b0000000000000000;
	sram_mem[106840] = 16'b0000000000000000;
	sram_mem[106841] = 16'b0000000000000000;
	sram_mem[106842] = 16'b0000000000000000;
	sram_mem[106843] = 16'b0000000000000000;
	sram_mem[106844] = 16'b0000000000000000;
	sram_mem[106845] = 16'b0000000000000000;
	sram_mem[106846] = 16'b0000000000000000;
	sram_mem[106847] = 16'b0000000000000000;
	sram_mem[106848] = 16'b0000000000000000;
	sram_mem[106849] = 16'b0000000000000000;
	sram_mem[106850] = 16'b0000000000000000;
	sram_mem[106851] = 16'b0000000000000000;
	sram_mem[106852] = 16'b0000000000000000;
	sram_mem[106853] = 16'b0000000000000000;
	sram_mem[106854] = 16'b0000000000000000;
	sram_mem[106855] = 16'b0000000000000000;
	sram_mem[106856] = 16'b0000000000000000;
	sram_mem[106857] = 16'b0000000000000000;
	sram_mem[106858] = 16'b0000000000000000;
	sram_mem[106859] = 16'b0000000000000000;
	sram_mem[106860] = 16'b0000000000000000;
	sram_mem[106861] = 16'b0000000000000000;
	sram_mem[106862] = 16'b0000000000000000;
	sram_mem[106863] = 16'b0000000000000000;
	sram_mem[106864] = 16'b0000000000000000;
	sram_mem[106865] = 16'b0000000000000000;
	sram_mem[106866] = 16'b0000000000000000;
	sram_mem[106867] = 16'b0000000000000000;
	sram_mem[106868] = 16'b0000000000000000;
	sram_mem[106869] = 16'b0000000000000000;
	sram_mem[106870] = 16'b0000000000000000;
	sram_mem[106871] = 16'b0000000000000000;
	sram_mem[106872] = 16'b0000000000000000;
	sram_mem[106873] = 16'b0000000000000000;
	sram_mem[106874] = 16'b0000000000000000;
	sram_mem[106875] = 16'b0000000000000000;
	sram_mem[106876] = 16'b0000000000000000;
	sram_mem[106877] = 16'b0000000000000000;
	sram_mem[106878] = 16'b0000000000000000;
	sram_mem[106879] = 16'b0000000000000000;
	sram_mem[106880] = 16'b0000000000000000;
	sram_mem[106881] = 16'b0000000000000000;
	sram_mem[106882] = 16'b0000000000000000;
	sram_mem[106883] = 16'b0000000000000000;
	sram_mem[106884] = 16'b0000000000000000;
	sram_mem[106885] = 16'b0000000000000000;
	sram_mem[106886] = 16'b0000000000000000;
	sram_mem[106887] = 16'b0000000000000000;
	sram_mem[106888] = 16'b0000000000000000;
	sram_mem[106889] = 16'b0000000000000000;
	sram_mem[106890] = 16'b0000000000000000;
	sram_mem[106891] = 16'b0000000000000000;
	sram_mem[106892] = 16'b0000000000000000;
	sram_mem[106893] = 16'b0000000000000000;
	sram_mem[106894] = 16'b0000000000000000;
	sram_mem[106895] = 16'b0000000000000000;
	sram_mem[106896] = 16'b0000000000000000;
	sram_mem[106897] = 16'b0000000000000000;
	sram_mem[106898] = 16'b0000000000000000;
	sram_mem[106899] = 16'b0000000000000000;
	sram_mem[106900] = 16'b0000000000000000;
	sram_mem[106901] = 16'b0000000000000000;
	sram_mem[106902] = 16'b0000000000000000;
	sram_mem[106903] = 16'b0000000000000000;
	sram_mem[106904] = 16'b0000000000000000;
	sram_mem[106905] = 16'b0000000000000000;
	sram_mem[106906] = 16'b0000000000000000;
	sram_mem[106907] = 16'b0000000000000000;
	sram_mem[106908] = 16'b0000000000000000;
	sram_mem[106909] = 16'b0000000000000000;
	sram_mem[106910] = 16'b0000000000000000;
	sram_mem[106911] = 16'b0000000000000000;
	sram_mem[106912] = 16'b0000000000000000;
	sram_mem[106913] = 16'b0000000000000000;
	sram_mem[106914] = 16'b0000000000000000;
	sram_mem[106915] = 16'b0000000000000000;
	sram_mem[106916] = 16'b0000000000000000;
	sram_mem[106917] = 16'b0000000000000000;
	sram_mem[106918] = 16'b0000000000000000;
	sram_mem[106919] = 16'b0000000000000000;
	sram_mem[106920] = 16'b0000000000000000;
	sram_mem[106921] = 16'b0000000000000000;
	sram_mem[106922] = 16'b0000000000000000;
	sram_mem[106923] = 16'b0000000000000000;
	sram_mem[106924] = 16'b0000000000000000;
	sram_mem[106925] = 16'b0000000000000000;
	sram_mem[106926] = 16'b0000000000000000;
	sram_mem[106927] = 16'b0000000000000000;
	sram_mem[106928] = 16'b0000000000000000;
	sram_mem[106929] = 16'b0000000000000000;
	sram_mem[106930] = 16'b0000000000000000;
	sram_mem[106931] = 16'b0000000000000000;
	sram_mem[106932] = 16'b0000000000000000;
	sram_mem[106933] = 16'b0000000000000000;
	sram_mem[106934] = 16'b0000000000000000;
	sram_mem[106935] = 16'b0000000000000000;
	sram_mem[106936] = 16'b0000000000000000;
	sram_mem[106937] = 16'b0000000000000000;
	sram_mem[106938] = 16'b0000000000000000;
	sram_mem[106939] = 16'b0000000000000000;
	sram_mem[106940] = 16'b0000000000000000;
	sram_mem[106941] = 16'b0000000000000000;
	sram_mem[106942] = 16'b0000000000000000;
	sram_mem[106943] = 16'b0000000000000000;
	sram_mem[106944] = 16'b0000000000000000;
	sram_mem[106945] = 16'b0000000000000000;
	sram_mem[106946] = 16'b0000000000000000;
	sram_mem[106947] = 16'b0000000000000000;
	sram_mem[106948] = 16'b0000000000000000;
	sram_mem[106949] = 16'b0000000000000000;
	sram_mem[106950] = 16'b0000000000000000;
	sram_mem[106951] = 16'b0000000000000000;
	sram_mem[106952] = 16'b0000000000000000;
	sram_mem[106953] = 16'b0000000000000000;
	sram_mem[106954] = 16'b0000000000000000;
	sram_mem[106955] = 16'b0000000000000000;
	sram_mem[106956] = 16'b0000000000000000;
	sram_mem[106957] = 16'b0000000000000000;
	sram_mem[106958] = 16'b0000000000000000;
	sram_mem[106959] = 16'b0000000000000000;
	sram_mem[106960] = 16'b0000000000000000;
	sram_mem[106961] = 16'b0000000000000000;
	sram_mem[106962] = 16'b0000000000000000;
	sram_mem[106963] = 16'b0000000000000000;
	sram_mem[106964] = 16'b0000000000000000;
	sram_mem[106965] = 16'b0000000000000000;
	sram_mem[106966] = 16'b0000000000000000;
	sram_mem[106967] = 16'b0000000000000000;
	sram_mem[106968] = 16'b0000000000000000;
	sram_mem[106969] = 16'b0000000000000000;
	sram_mem[106970] = 16'b0000000000000000;
	sram_mem[106971] = 16'b0000000000000000;
	sram_mem[106972] = 16'b0000000000000000;
	sram_mem[106973] = 16'b0000000000000000;
	sram_mem[106974] = 16'b0000000000000000;
	sram_mem[106975] = 16'b0000000000000000;
	sram_mem[106976] = 16'b0000000000000000;
	sram_mem[106977] = 16'b0000000000000000;
	sram_mem[106978] = 16'b0000000000000000;
	sram_mem[106979] = 16'b0000000000000000;
	sram_mem[106980] = 16'b0000000000000000;
	sram_mem[106981] = 16'b0000000000000000;
	sram_mem[106982] = 16'b0000000000000000;
	sram_mem[106983] = 16'b0000000000000000;
	sram_mem[106984] = 16'b0000000000000000;
	sram_mem[106985] = 16'b0000000000000000;
	sram_mem[106986] = 16'b0000000000000000;
	sram_mem[106987] = 16'b0000000000000000;
	sram_mem[106988] = 16'b0000000000000000;
	sram_mem[106989] = 16'b0000000000000000;
	sram_mem[106990] = 16'b0000000000000000;
	sram_mem[106991] = 16'b0000000000000000;
	sram_mem[106992] = 16'b0000000000000000;
	sram_mem[106993] = 16'b0000000000000000;
	sram_mem[106994] = 16'b0000000000000000;
	sram_mem[106995] = 16'b0000000000000000;
	sram_mem[106996] = 16'b0000000000000000;
	sram_mem[106997] = 16'b0000000000000000;
	sram_mem[106998] = 16'b0000000000000000;
	sram_mem[106999] = 16'b0000000000000000;
	sram_mem[107000] = 16'b0000000000000000;
	sram_mem[107001] = 16'b0000000000000000;
	sram_mem[107002] = 16'b0000000000000000;
	sram_mem[107003] = 16'b0000000000000000;
	sram_mem[107004] = 16'b0000000000000000;
	sram_mem[107005] = 16'b0000000000000000;
	sram_mem[107006] = 16'b0000000000000000;
	sram_mem[107007] = 16'b0000000000000000;
	sram_mem[107008] = 16'b0000000000000000;
	sram_mem[107009] = 16'b0000000000000000;
	sram_mem[107010] = 16'b0000000000000000;
	sram_mem[107011] = 16'b0000000000000000;
	sram_mem[107012] = 16'b0000000000000000;
	sram_mem[107013] = 16'b0000000000000000;
	sram_mem[107014] = 16'b0000000000000000;
	sram_mem[107015] = 16'b0000000000000000;
	sram_mem[107016] = 16'b0000000000000000;
	sram_mem[107017] = 16'b0000000000000000;
	sram_mem[107018] = 16'b0000000000000000;
	sram_mem[107019] = 16'b0000000000000000;
	sram_mem[107020] = 16'b0000000000000000;
	sram_mem[107021] = 16'b0000000000000000;
	sram_mem[107022] = 16'b0000000000000000;
	sram_mem[107023] = 16'b0000000000000000;
	sram_mem[107024] = 16'b0000000000000000;
	sram_mem[107025] = 16'b0000000000000000;
	sram_mem[107026] = 16'b0000000000000000;
	sram_mem[107027] = 16'b0000000000000000;
	sram_mem[107028] = 16'b0000000000000000;
	sram_mem[107029] = 16'b0000000000000000;
	sram_mem[107030] = 16'b0000000000000000;
	sram_mem[107031] = 16'b0000000000000000;
	sram_mem[107032] = 16'b0000000000000000;
	sram_mem[107033] = 16'b0000000000000000;
	sram_mem[107034] = 16'b0000000000000000;
	sram_mem[107035] = 16'b0000000000000000;
	sram_mem[107036] = 16'b0000000000000000;
	sram_mem[107037] = 16'b0000000000000000;
	sram_mem[107038] = 16'b0000000000000000;
	sram_mem[107039] = 16'b0000000000000000;
	sram_mem[107040] = 16'b0000000000000000;
	sram_mem[107041] = 16'b0000000000000000;
	sram_mem[107042] = 16'b0000000000000000;
	sram_mem[107043] = 16'b0000000000000000;
	sram_mem[107044] = 16'b0000000000000000;
	sram_mem[107045] = 16'b0000000000000000;
	sram_mem[107046] = 16'b0000000000000000;
	sram_mem[107047] = 16'b0000000000000000;
	sram_mem[107048] = 16'b0000000000000000;
	sram_mem[107049] = 16'b0000000000000000;
	sram_mem[107050] = 16'b0000000000000000;
	sram_mem[107051] = 16'b0000000000000000;
	sram_mem[107052] = 16'b0000000000000000;
	sram_mem[107053] = 16'b0000000000000000;
	sram_mem[107054] = 16'b0000000000000000;
	sram_mem[107055] = 16'b0000000000000000;
	sram_mem[107056] = 16'b0000000000000000;
	sram_mem[107057] = 16'b0000000000000000;
	sram_mem[107058] = 16'b0000000000000000;
	sram_mem[107059] = 16'b0000000000000000;
	sram_mem[107060] = 16'b0000000000000000;
	sram_mem[107061] = 16'b0000000000000000;
	sram_mem[107062] = 16'b0000000000000000;
	sram_mem[107063] = 16'b0000000000000000;
	sram_mem[107064] = 16'b0000000000000000;
	sram_mem[107065] = 16'b0000000000000000;
	sram_mem[107066] = 16'b0000000000000000;
	sram_mem[107067] = 16'b0000000000000000;
	sram_mem[107068] = 16'b0000000000000000;
	sram_mem[107069] = 16'b0000000000000000;
	sram_mem[107070] = 16'b0000000000000000;
	sram_mem[107071] = 16'b0000000000000000;
	sram_mem[107072] = 16'b0000000000000000;
	sram_mem[107073] = 16'b0000000000000000;
	sram_mem[107074] = 16'b0000000000000000;
	sram_mem[107075] = 16'b0000000000000000;
	sram_mem[107076] = 16'b0000000000000000;
	sram_mem[107077] = 16'b0000000000000000;
	sram_mem[107078] = 16'b0000000000000000;
	sram_mem[107079] = 16'b0000000000000000;
	sram_mem[107080] = 16'b0000000000000000;
	sram_mem[107081] = 16'b0000000000000000;
	sram_mem[107082] = 16'b0000000000000000;
	sram_mem[107083] = 16'b0000000000000000;
	sram_mem[107084] = 16'b0000000000000000;
	sram_mem[107085] = 16'b0000000000000000;
	sram_mem[107086] = 16'b0000000000000000;
	sram_mem[107087] = 16'b0000000000000000;
	sram_mem[107088] = 16'b0000000000000000;
	sram_mem[107089] = 16'b0000000000000000;
	sram_mem[107090] = 16'b0000000000000000;
	sram_mem[107091] = 16'b0000000000000000;
	sram_mem[107092] = 16'b0000000000000000;
	sram_mem[107093] = 16'b0000000000000000;
	sram_mem[107094] = 16'b0000000000000000;
	sram_mem[107095] = 16'b0000000000000000;
	sram_mem[107096] = 16'b0000000000000000;
	sram_mem[107097] = 16'b0000000000000000;
	sram_mem[107098] = 16'b0000000000000000;
	sram_mem[107099] = 16'b0000000000000000;
	sram_mem[107100] = 16'b0000000000000000;
	sram_mem[107101] = 16'b0000000000000000;
	sram_mem[107102] = 16'b0000000000000000;
	sram_mem[107103] = 16'b0000000000000000;
	sram_mem[107104] = 16'b0000000000000000;
	sram_mem[107105] = 16'b0000000000000000;
	sram_mem[107106] = 16'b0000000000000000;
	sram_mem[107107] = 16'b0000000000000000;
	sram_mem[107108] = 16'b0000000000000000;
	sram_mem[107109] = 16'b0000000000000000;
	sram_mem[107110] = 16'b0000000000000000;
	sram_mem[107111] = 16'b0000000000000000;
	sram_mem[107112] = 16'b0000000000000000;
	sram_mem[107113] = 16'b0000000000000000;
	sram_mem[107114] = 16'b0000000000000000;
	sram_mem[107115] = 16'b0000000000000000;
	sram_mem[107116] = 16'b0000000000000000;
	sram_mem[107117] = 16'b0000000000000000;
	sram_mem[107118] = 16'b0000000000000000;
	sram_mem[107119] = 16'b0000000000000000;
	sram_mem[107120] = 16'b0000000000000000;
	sram_mem[107121] = 16'b0000000000000000;
	sram_mem[107122] = 16'b0000000000000000;
	sram_mem[107123] = 16'b0000000000000000;
	sram_mem[107124] = 16'b0000000000000000;
	sram_mem[107125] = 16'b0000000000000000;
	sram_mem[107126] = 16'b0000000000000000;
	sram_mem[107127] = 16'b0000000000000000;
	sram_mem[107128] = 16'b0000000000000000;
	sram_mem[107129] = 16'b0000000000000000;
	sram_mem[107130] = 16'b0000000000000000;
	sram_mem[107131] = 16'b0000000000000000;
	sram_mem[107132] = 16'b0000000000000000;
	sram_mem[107133] = 16'b0000000000000000;
	sram_mem[107134] = 16'b0000000000000000;
	sram_mem[107135] = 16'b0000000000000000;
	sram_mem[107136] = 16'b0000000000000000;
	sram_mem[107137] = 16'b0000000000000000;
	sram_mem[107138] = 16'b0000000000000000;
	sram_mem[107139] = 16'b0000000000000000;
	sram_mem[107140] = 16'b0000000000000000;
	sram_mem[107141] = 16'b0000000000000000;
	sram_mem[107142] = 16'b0000000000000000;
	sram_mem[107143] = 16'b0000000000000000;
	sram_mem[107144] = 16'b0000000000000000;
	sram_mem[107145] = 16'b0000000000000000;
	sram_mem[107146] = 16'b0000000000000000;
	sram_mem[107147] = 16'b0000000000000000;
	sram_mem[107148] = 16'b0000000000000000;
	sram_mem[107149] = 16'b0000000000000000;
	sram_mem[107150] = 16'b0000000000000000;
	sram_mem[107151] = 16'b0000000000000000;
	sram_mem[107152] = 16'b0000000000000000;
	sram_mem[107153] = 16'b0000000000000000;
	sram_mem[107154] = 16'b0000000000000000;
	sram_mem[107155] = 16'b0000000000000000;
	sram_mem[107156] = 16'b0000000000000000;
	sram_mem[107157] = 16'b0000000000000000;
	sram_mem[107158] = 16'b0000000000000000;
	sram_mem[107159] = 16'b0000000000000000;
	sram_mem[107160] = 16'b0000000000000000;
	sram_mem[107161] = 16'b0000000000000000;
	sram_mem[107162] = 16'b0000000000000000;
	sram_mem[107163] = 16'b0000000000000000;
	sram_mem[107164] = 16'b0000000000000000;
	sram_mem[107165] = 16'b0000000000000000;
	sram_mem[107166] = 16'b0000000000000000;
	sram_mem[107167] = 16'b0000000000000000;
	sram_mem[107168] = 16'b0000000000000000;
	sram_mem[107169] = 16'b0000000000000000;
	sram_mem[107170] = 16'b0000000000000000;
	sram_mem[107171] = 16'b0000000000000000;
	sram_mem[107172] = 16'b0000000000000000;
	sram_mem[107173] = 16'b0000000000000000;
	sram_mem[107174] = 16'b0000000000000000;
	sram_mem[107175] = 16'b0000000000000000;
	sram_mem[107176] = 16'b0000000000000000;
	sram_mem[107177] = 16'b0000000000000000;
	sram_mem[107178] = 16'b0000000000000000;
	sram_mem[107179] = 16'b0000000000000000;
	sram_mem[107180] = 16'b0000000000000000;
	sram_mem[107181] = 16'b0000000000000000;
	sram_mem[107182] = 16'b0000000000000000;
	sram_mem[107183] = 16'b0000000000000000;
	sram_mem[107184] = 16'b0000000000000000;
	sram_mem[107185] = 16'b0000000000000000;
	sram_mem[107186] = 16'b0000000000000000;
	sram_mem[107187] = 16'b0000000000000000;
	sram_mem[107188] = 16'b0000000000000000;
	sram_mem[107189] = 16'b0000000000000000;
	sram_mem[107190] = 16'b0000000000000000;
	sram_mem[107191] = 16'b0000000000000000;
	sram_mem[107192] = 16'b0000000000000000;
	sram_mem[107193] = 16'b0000000000000000;
	sram_mem[107194] = 16'b0000000000000000;
	sram_mem[107195] = 16'b0000000000000000;
	sram_mem[107196] = 16'b0000000000000000;
	sram_mem[107197] = 16'b0000000000000000;
	sram_mem[107198] = 16'b0000000000000000;
	sram_mem[107199] = 16'b0000000000000000;
	sram_mem[107200] = 16'b0000000000000000;
	sram_mem[107201] = 16'b0000000000000000;
	sram_mem[107202] = 16'b0000000000000000;
	sram_mem[107203] = 16'b0000000000000000;
	sram_mem[107204] = 16'b0000000000000000;
	sram_mem[107205] = 16'b0000000000000000;
	sram_mem[107206] = 16'b0000000000000000;
	sram_mem[107207] = 16'b0000000000000000;
	sram_mem[107208] = 16'b0000000000000000;
	sram_mem[107209] = 16'b0000000000000000;
	sram_mem[107210] = 16'b0000000000000000;
	sram_mem[107211] = 16'b0000000000000000;
	sram_mem[107212] = 16'b0000000000000000;
	sram_mem[107213] = 16'b0000000000000000;
	sram_mem[107214] = 16'b0000000000000000;
	sram_mem[107215] = 16'b0000000000000000;
	sram_mem[107216] = 16'b0000000000000000;
	sram_mem[107217] = 16'b0000000000000000;
	sram_mem[107218] = 16'b0000000000000000;
	sram_mem[107219] = 16'b0000000000000000;
	sram_mem[107220] = 16'b0000000000000000;
	sram_mem[107221] = 16'b0000000000000000;
	sram_mem[107222] = 16'b0000000000000000;
	sram_mem[107223] = 16'b0000000000000000;
	sram_mem[107224] = 16'b0000000000000000;
	sram_mem[107225] = 16'b0000000000000000;
	sram_mem[107226] = 16'b0000000000000000;
	sram_mem[107227] = 16'b0000000000000000;
	sram_mem[107228] = 16'b0000000000000000;
	sram_mem[107229] = 16'b0000000000000000;
	sram_mem[107230] = 16'b0000000000000000;
	sram_mem[107231] = 16'b0000000000000000;
	sram_mem[107232] = 16'b0000000000000000;
	sram_mem[107233] = 16'b0000000000000000;
	sram_mem[107234] = 16'b0000000000000000;
	sram_mem[107235] = 16'b0000000000000000;
	sram_mem[107236] = 16'b0000000000000000;
	sram_mem[107237] = 16'b0000000000000000;
	sram_mem[107238] = 16'b0000000000000000;
	sram_mem[107239] = 16'b0000000000000000;
	sram_mem[107240] = 16'b0000000000000000;
	sram_mem[107241] = 16'b0000000000000000;
	sram_mem[107242] = 16'b0000000000000000;
	sram_mem[107243] = 16'b0000000000000000;
	sram_mem[107244] = 16'b0000000000000000;
	sram_mem[107245] = 16'b0000000000000000;
	sram_mem[107246] = 16'b0000000000000000;
	sram_mem[107247] = 16'b0000000000000000;
	sram_mem[107248] = 16'b0000000000000000;
	sram_mem[107249] = 16'b0000000000000000;
	sram_mem[107250] = 16'b0000000000000000;
	sram_mem[107251] = 16'b0000000000000000;
	sram_mem[107252] = 16'b0000000000000000;
	sram_mem[107253] = 16'b0000000000000000;
	sram_mem[107254] = 16'b0000000000000000;
	sram_mem[107255] = 16'b0000000000000000;
	sram_mem[107256] = 16'b0000000000000000;
	sram_mem[107257] = 16'b0000000000000000;
	sram_mem[107258] = 16'b0000000000000000;
	sram_mem[107259] = 16'b0000000000000000;
	sram_mem[107260] = 16'b0000000000000000;
	sram_mem[107261] = 16'b0000000000000000;
	sram_mem[107262] = 16'b0000000000000000;
	sram_mem[107263] = 16'b0000000000000000;
	sram_mem[107264] = 16'b0000000000000000;
	sram_mem[107265] = 16'b0000000000000000;
	sram_mem[107266] = 16'b0000000000000000;
	sram_mem[107267] = 16'b0000000000000000;
	sram_mem[107268] = 16'b0000000000000000;
	sram_mem[107269] = 16'b0000000000000000;
	sram_mem[107270] = 16'b0000000000000000;
	sram_mem[107271] = 16'b0000000000000000;
	sram_mem[107272] = 16'b0000000000000000;
	sram_mem[107273] = 16'b0000000000000000;
	sram_mem[107274] = 16'b0000000000000000;
	sram_mem[107275] = 16'b0000000000000000;
	sram_mem[107276] = 16'b0000000000000000;
	sram_mem[107277] = 16'b0000000000000000;
	sram_mem[107278] = 16'b0000000000000000;
	sram_mem[107279] = 16'b0000000000000000;
	sram_mem[107280] = 16'b0000000000000000;
	sram_mem[107281] = 16'b0000000000000000;
	sram_mem[107282] = 16'b0000000000000000;
	sram_mem[107283] = 16'b0000000000000000;
	sram_mem[107284] = 16'b0000000000000000;
	sram_mem[107285] = 16'b0000000000000000;
	sram_mem[107286] = 16'b0000000000000000;
	sram_mem[107287] = 16'b0000000000000000;
	sram_mem[107288] = 16'b0000000000000000;
	sram_mem[107289] = 16'b0000000000000000;
	sram_mem[107290] = 16'b0000000000000000;
	sram_mem[107291] = 16'b0000000000000000;
	sram_mem[107292] = 16'b0000000000000000;
	sram_mem[107293] = 16'b0000000000000000;
	sram_mem[107294] = 16'b0000000000000000;
	sram_mem[107295] = 16'b0000000000000000;
	sram_mem[107296] = 16'b0000000000000000;
	sram_mem[107297] = 16'b0000000000000000;
	sram_mem[107298] = 16'b0000000000000000;
	sram_mem[107299] = 16'b0000000000000000;
	sram_mem[107300] = 16'b0000000000000000;
	sram_mem[107301] = 16'b0000000000000000;
	sram_mem[107302] = 16'b0000000000000000;
	sram_mem[107303] = 16'b0000000000000000;
	sram_mem[107304] = 16'b0000000000000000;
	sram_mem[107305] = 16'b0000000000000000;
	sram_mem[107306] = 16'b0000000000000000;
	sram_mem[107307] = 16'b0000000000000000;
	sram_mem[107308] = 16'b0000000000000000;
	sram_mem[107309] = 16'b0000000000000000;
	sram_mem[107310] = 16'b0000000000000000;
	sram_mem[107311] = 16'b0000000000000000;
	sram_mem[107312] = 16'b0000000000000000;
	sram_mem[107313] = 16'b0000000000000000;
	sram_mem[107314] = 16'b0000000000000000;
	sram_mem[107315] = 16'b0000000000000000;
	sram_mem[107316] = 16'b0000000000000000;
	sram_mem[107317] = 16'b0000000000000000;
	sram_mem[107318] = 16'b0000000000000000;
	sram_mem[107319] = 16'b0000000000000000;
	sram_mem[107320] = 16'b0000000000000000;
	sram_mem[107321] = 16'b0000000000000000;
	sram_mem[107322] = 16'b0000000000000000;
	sram_mem[107323] = 16'b0000000000000000;
	sram_mem[107324] = 16'b0000000000000000;
	sram_mem[107325] = 16'b0000000000000000;
	sram_mem[107326] = 16'b0000000000000000;
	sram_mem[107327] = 16'b0000000000000000;
	sram_mem[107328] = 16'b0000000000000000;
	sram_mem[107329] = 16'b0000000000000000;
	sram_mem[107330] = 16'b0000000000000000;
	sram_mem[107331] = 16'b0000000000000000;
	sram_mem[107332] = 16'b0000000000000000;
	sram_mem[107333] = 16'b0000000000000000;
	sram_mem[107334] = 16'b0000000000000000;
	sram_mem[107335] = 16'b0000000000000000;
	sram_mem[107336] = 16'b0000000000000000;
	sram_mem[107337] = 16'b0000000000000000;
	sram_mem[107338] = 16'b0000000000000000;
	sram_mem[107339] = 16'b0000000000000000;
	sram_mem[107340] = 16'b0000000000000000;
	sram_mem[107341] = 16'b0000000000000000;
	sram_mem[107342] = 16'b0000000000000000;
	sram_mem[107343] = 16'b0000000000000000;
	sram_mem[107344] = 16'b0000000000000000;
	sram_mem[107345] = 16'b0000000000000000;
	sram_mem[107346] = 16'b0000000000000000;
	sram_mem[107347] = 16'b0000000000000000;
	sram_mem[107348] = 16'b0000000000000000;
	sram_mem[107349] = 16'b0000000000000000;
	sram_mem[107350] = 16'b0000000000000000;
	sram_mem[107351] = 16'b0000000000000000;
	sram_mem[107352] = 16'b0000000000000000;
	sram_mem[107353] = 16'b0000000000000000;
	sram_mem[107354] = 16'b0000000000000000;
	sram_mem[107355] = 16'b0000000000000000;
	sram_mem[107356] = 16'b0000000000000000;
	sram_mem[107357] = 16'b0000000000000000;
	sram_mem[107358] = 16'b0000000000000000;
	sram_mem[107359] = 16'b0000000000000000;
	sram_mem[107360] = 16'b0000000000000000;
	sram_mem[107361] = 16'b0000000000000000;
	sram_mem[107362] = 16'b0000000000000000;
	sram_mem[107363] = 16'b0000000000000000;
	sram_mem[107364] = 16'b0000000000000000;
	sram_mem[107365] = 16'b0000000000000000;
	sram_mem[107366] = 16'b0000000000000000;
	sram_mem[107367] = 16'b0000000000000000;
	sram_mem[107368] = 16'b0000000000000000;
	sram_mem[107369] = 16'b0000000000000000;
	sram_mem[107370] = 16'b0000000000000000;
	sram_mem[107371] = 16'b0000000000000000;
	sram_mem[107372] = 16'b0000000000000000;
	sram_mem[107373] = 16'b0000000000000000;
	sram_mem[107374] = 16'b0000000000000000;
	sram_mem[107375] = 16'b0000000000000000;
	sram_mem[107376] = 16'b0000000000000000;
	sram_mem[107377] = 16'b0000000000000000;
	sram_mem[107378] = 16'b0000000000000000;
	sram_mem[107379] = 16'b0000000000000000;
	sram_mem[107380] = 16'b0000000000000000;
	sram_mem[107381] = 16'b0000000000000000;
	sram_mem[107382] = 16'b0000000000000000;
	sram_mem[107383] = 16'b0000000000000000;
	sram_mem[107384] = 16'b0000000000000000;
	sram_mem[107385] = 16'b0000000000000000;
	sram_mem[107386] = 16'b0000000000000000;
	sram_mem[107387] = 16'b0000000000000000;
	sram_mem[107388] = 16'b0000000000000000;
	sram_mem[107389] = 16'b0000000000000000;
	sram_mem[107390] = 16'b0000000000000000;
	sram_mem[107391] = 16'b0000000000000000;
	sram_mem[107392] = 16'b0000000000000000;
	sram_mem[107393] = 16'b0000000000000000;
	sram_mem[107394] = 16'b0000000000000000;
	sram_mem[107395] = 16'b0000000000000000;
	sram_mem[107396] = 16'b0000000000000000;
	sram_mem[107397] = 16'b0000000000000000;
	sram_mem[107398] = 16'b0000000000000000;
	sram_mem[107399] = 16'b0000000000000000;
	sram_mem[107400] = 16'b0000000000000000;
	sram_mem[107401] = 16'b0000000000000000;
	sram_mem[107402] = 16'b0000000000000000;
	sram_mem[107403] = 16'b0000000000000000;
	sram_mem[107404] = 16'b0000000000000000;
	sram_mem[107405] = 16'b0000000000000000;
	sram_mem[107406] = 16'b0000000000000000;
	sram_mem[107407] = 16'b0000000000000000;
	sram_mem[107408] = 16'b0000000000000000;
	sram_mem[107409] = 16'b0000000000000000;
	sram_mem[107410] = 16'b0000000000000000;
	sram_mem[107411] = 16'b0000000000000000;
	sram_mem[107412] = 16'b0000000000000000;
	sram_mem[107413] = 16'b0000000000000000;
	sram_mem[107414] = 16'b0000000000000000;
	sram_mem[107415] = 16'b0000000000000000;
	sram_mem[107416] = 16'b0000000000000000;
	sram_mem[107417] = 16'b0000000000000000;
	sram_mem[107418] = 16'b0000000000000000;
	sram_mem[107419] = 16'b0000000000000000;
	sram_mem[107420] = 16'b0000000000000000;
	sram_mem[107421] = 16'b0000000000000000;
	sram_mem[107422] = 16'b0000000000000000;
	sram_mem[107423] = 16'b0000000000000000;
	sram_mem[107424] = 16'b0000000000000000;
	sram_mem[107425] = 16'b0000000000000000;
	sram_mem[107426] = 16'b0000000000000000;
	sram_mem[107427] = 16'b0000000000000000;
	sram_mem[107428] = 16'b0000000000000000;
	sram_mem[107429] = 16'b0000000000000000;
	sram_mem[107430] = 16'b0000000000000000;
	sram_mem[107431] = 16'b0000000000000000;
	sram_mem[107432] = 16'b0000000000000000;
	sram_mem[107433] = 16'b0000000000000000;
	sram_mem[107434] = 16'b0000000000000000;
	sram_mem[107435] = 16'b0000000000000000;
	sram_mem[107436] = 16'b0000000000000000;
	sram_mem[107437] = 16'b0000000000000000;
	sram_mem[107438] = 16'b0000000000000000;
	sram_mem[107439] = 16'b0000000000000000;
	sram_mem[107440] = 16'b0000000000000000;
	sram_mem[107441] = 16'b0000000000000000;
	sram_mem[107442] = 16'b0000000000000000;
	sram_mem[107443] = 16'b0000000000000000;
	sram_mem[107444] = 16'b0000000000000000;
	sram_mem[107445] = 16'b0000000000000000;
	sram_mem[107446] = 16'b0000000000000000;
	sram_mem[107447] = 16'b0000000000000000;
	sram_mem[107448] = 16'b0000000000000000;
	sram_mem[107449] = 16'b0000000000000000;
	sram_mem[107450] = 16'b0000000000000000;
	sram_mem[107451] = 16'b0000000000000000;
	sram_mem[107452] = 16'b0000000000000000;
	sram_mem[107453] = 16'b0000000000000000;
	sram_mem[107454] = 16'b0000000000000000;
	sram_mem[107455] = 16'b0000000000000000;
	sram_mem[107456] = 16'b0000000000000000;
	sram_mem[107457] = 16'b0000000000000000;
	sram_mem[107458] = 16'b0000000000000000;
	sram_mem[107459] = 16'b0000000000000000;
	sram_mem[107460] = 16'b0000000000000000;
	sram_mem[107461] = 16'b0000000000000000;
	sram_mem[107462] = 16'b0000000000000000;
	sram_mem[107463] = 16'b0000000000000000;
	sram_mem[107464] = 16'b0000000000000000;
	sram_mem[107465] = 16'b0000000000000000;
	sram_mem[107466] = 16'b0000000000000000;
	sram_mem[107467] = 16'b0000000000000000;
	sram_mem[107468] = 16'b0000000000000000;
	sram_mem[107469] = 16'b0000000000000000;
	sram_mem[107470] = 16'b0000000000000000;
	sram_mem[107471] = 16'b0000000000000000;
	sram_mem[107472] = 16'b0000000000000000;
	sram_mem[107473] = 16'b0000000000000000;
	sram_mem[107474] = 16'b0000000000000000;
	sram_mem[107475] = 16'b0000000000000000;
	sram_mem[107476] = 16'b0000000000000000;
	sram_mem[107477] = 16'b0000000000000000;
	sram_mem[107478] = 16'b0000000000000000;
	sram_mem[107479] = 16'b0000000000000000;
	sram_mem[107480] = 16'b0000000000000000;
	sram_mem[107481] = 16'b0000000000000000;
	sram_mem[107482] = 16'b0000000000000000;
	sram_mem[107483] = 16'b0000000000000000;
	sram_mem[107484] = 16'b0000000000000000;
	sram_mem[107485] = 16'b0000000000000000;
	sram_mem[107486] = 16'b0000000000000000;
	sram_mem[107487] = 16'b0000000000000000;
	sram_mem[107488] = 16'b0000000000000000;
	sram_mem[107489] = 16'b0000000000000000;
	sram_mem[107490] = 16'b0000000000000000;
	sram_mem[107491] = 16'b0000000000000000;
	sram_mem[107492] = 16'b0000000000000000;
	sram_mem[107493] = 16'b0000000000000000;
	sram_mem[107494] = 16'b0000000000000000;
	sram_mem[107495] = 16'b0000000000000000;
	sram_mem[107496] = 16'b0000000000000000;
	sram_mem[107497] = 16'b0000000000000000;
	sram_mem[107498] = 16'b0000000000000000;
	sram_mem[107499] = 16'b0000000000000000;
	sram_mem[107500] = 16'b0000000000000000;
	sram_mem[107501] = 16'b0000000000000000;
	sram_mem[107502] = 16'b0000000000000000;
	sram_mem[107503] = 16'b0000000000000000;
	sram_mem[107504] = 16'b0000000000000000;
	sram_mem[107505] = 16'b0000000000000000;
	sram_mem[107506] = 16'b0000000000000000;
	sram_mem[107507] = 16'b0000000000000000;
	sram_mem[107508] = 16'b0000000000000000;
	sram_mem[107509] = 16'b0000000000000000;
	sram_mem[107510] = 16'b0000000000000000;
	sram_mem[107511] = 16'b0000000000000000;
	sram_mem[107512] = 16'b0000000000000000;
	sram_mem[107513] = 16'b0000000000000000;
	sram_mem[107514] = 16'b0000000000000000;
	sram_mem[107515] = 16'b0000000000000000;
	sram_mem[107516] = 16'b0000000000000000;
	sram_mem[107517] = 16'b0000000000000000;
	sram_mem[107518] = 16'b0000000000000000;
	sram_mem[107519] = 16'b0000000000000000;
	sram_mem[107520] = 16'b0000000000000000;
	sram_mem[107521] = 16'b0000000000000000;
	sram_mem[107522] = 16'b0000000000000000;
	sram_mem[107523] = 16'b0000000000000000;
	sram_mem[107524] = 16'b0000000000000000;
	sram_mem[107525] = 16'b0000000000000000;
	sram_mem[107526] = 16'b0000000000000000;
	sram_mem[107527] = 16'b0000000000000000;
	sram_mem[107528] = 16'b0000000000000000;
	sram_mem[107529] = 16'b0000000000000000;
	sram_mem[107530] = 16'b0000000000000000;
	sram_mem[107531] = 16'b0000000000000000;
	sram_mem[107532] = 16'b0000000000000000;
	sram_mem[107533] = 16'b0000000000000000;
	sram_mem[107534] = 16'b0000000000000000;
	sram_mem[107535] = 16'b0000000000000000;
	sram_mem[107536] = 16'b0000000000000000;
	sram_mem[107537] = 16'b0000000000000000;
	sram_mem[107538] = 16'b0000000000000000;
	sram_mem[107539] = 16'b0000000000000000;
	sram_mem[107540] = 16'b0000000000000000;
	sram_mem[107541] = 16'b0000000000000000;
	sram_mem[107542] = 16'b0000000000000000;
	sram_mem[107543] = 16'b0000000000000000;
	sram_mem[107544] = 16'b0000000000000000;
	sram_mem[107545] = 16'b0000000000000000;
	sram_mem[107546] = 16'b0000000000000000;
	sram_mem[107547] = 16'b0000000000000000;
	sram_mem[107548] = 16'b0000000000000000;
	sram_mem[107549] = 16'b0000000000000000;
	sram_mem[107550] = 16'b0000000000000000;
	sram_mem[107551] = 16'b0000000000000000;
	sram_mem[107552] = 16'b0000000000000000;
	sram_mem[107553] = 16'b0000000000000000;
	sram_mem[107554] = 16'b0000000000000000;
	sram_mem[107555] = 16'b0000000000000000;
	sram_mem[107556] = 16'b0000000000000000;
	sram_mem[107557] = 16'b0000000000000000;
	sram_mem[107558] = 16'b0000000000000000;
	sram_mem[107559] = 16'b0000000000000000;
	sram_mem[107560] = 16'b0000000000000000;
	sram_mem[107561] = 16'b0000000000000000;
	sram_mem[107562] = 16'b0000000000000000;
	sram_mem[107563] = 16'b0000000000000000;
	sram_mem[107564] = 16'b0000000000000000;
	sram_mem[107565] = 16'b0000000000000000;
	sram_mem[107566] = 16'b0000000000000000;
	sram_mem[107567] = 16'b0000000000000000;
	sram_mem[107568] = 16'b0000000000000000;
	sram_mem[107569] = 16'b0000000000000000;
	sram_mem[107570] = 16'b0000000000000000;
	sram_mem[107571] = 16'b0000000000000000;
	sram_mem[107572] = 16'b0000000000000000;
	sram_mem[107573] = 16'b0000000000000000;
	sram_mem[107574] = 16'b0000000000000000;
	sram_mem[107575] = 16'b0000000000000000;
	sram_mem[107576] = 16'b0000000000000000;
	sram_mem[107577] = 16'b0000000000000000;
	sram_mem[107578] = 16'b0000000000000000;
	sram_mem[107579] = 16'b0000000000000000;
	sram_mem[107580] = 16'b0000000000000000;
	sram_mem[107581] = 16'b0000000000000000;
	sram_mem[107582] = 16'b0000000000000000;
	sram_mem[107583] = 16'b0000000000000000;
	sram_mem[107584] = 16'b0000000000000000;
	sram_mem[107585] = 16'b0000000000000000;
	sram_mem[107586] = 16'b0000000000000000;
	sram_mem[107587] = 16'b0000000000000000;
	sram_mem[107588] = 16'b0000000000000000;
	sram_mem[107589] = 16'b0000000000000000;
	sram_mem[107590] = 16'b0000000000000000;
	sram_mem[107591] = 16'b0000000000000000;
	sram_mem[107592] = 16'b0000000000000000;
	sram_mem[107593] = 16'b0000000000000000;
	sram_mem[107594] = 16'b0000000000000000;
	sram_mem[107595] = 16'b0000000000000000;
	sram_mem[107596] = 16'b0000000000000000;
	sram_mem[107597] = 16'b0000000000000000;
	sram_mem[107598] = 16'b0000000000000000;
	sram_mem[107599] = 16'b0000000000000000;
	sram_mem[107600] = 16'b0000000000000000;
	sram_mem[107601] = 16'b0000000000000000;
	sram_mem[107602] = 16'b0000000000000000;
	sram_mem[107603] = 16'b0000000000000000;
	sram_mem[107604] = 16'b0000000000000000;
	sram_mem[107605] = 16'b0000000000000000;
	sram_mem[107606] = 16'b0000000000000000;
	sram_mem[107607] = 16'b0000000000000000;
	sram_mem[107608] = 16'b0000000000000000;
	sram_mem[107609] = 16'b0000000000000000;
	sram_mem[107610] = 16'b0000000000000000;
	sram_mem[107611] = 16'b0000000000000000;
	sram_mem[107612] = 16'b0000000000000000;
	sram_mem[107613] = 16'b0000000000000000;
	sram_mem[107614] = 16'b0000000000000000;
	sram_mem[107615] = 16'b0000000000000000;
	sram_mem[107616] = 16'b0000000000000000;
	sram_mem[107617] = 16'b0000000000000000;
	sram_mem[107618] = 16'b0000000000000000;
	sram_mem[107619] = 16'b0000000000000000;
	sram_mem[107620] = 16'b0000000000000000;
	sram_mem[107621] = 16'b0000000000000000;
	sram_mem[107622] = 16'b0000000000000000;
	sram_mem[107623] = 16'b0000000000000000;
	sram_mem[107624] = 16'b0000000000000000;
	sram_mem[107625] = 16'b0000000000000000;
	sram_mem[107626] = 16'b0000000000000000;
	sram_mem[107627] = 16'b0000000000000000;
	sram_mem[107628] = 16'b0000000000000000;
	sram_mem[107629] = 16'b0000000000000000;
	sram_mem[107630] = 16'b0000000000000000;
	sram_mem[107631] = 16'b0000000000000000;
	sram_mem[107632] = 16'b0000000000000000;
	sram_mem[107633] = 16'b0000000000000000;
	sram_mem[107634] = 16'b0000000000000000;
	sram_mem[107635] = 16'b0000000000000000;
	sram_mem[107636] = 16'b0000000000000000;
	sram_mem[107637] = 16'b0000000000000000;
	sram_mem[107638] = 16'b0000000000000000;
	sram_mem[107639] = 16'b0000000000000000;
	sram_mem[107640] = 16'b0000000000000000;
	sram_mem[107641] = 16'b0000000000000000;
	sram_mem[107642] = 16'b0000000000000000;
	sram_mem[107643] = 16'b0000000000000000;
	sram_mem[107644] = 16'b0000000000000000;
	sram_mem[107645] = 16'b0000000000000000;
	sram_mem[107646] = 16'b0000000000000000;
	sram_mem[107647] = 16'b0000000000000000;
	sram_mem[107648] = 16'b0000000000000000;
	sram_mem[107649] = 16'b0000000000000000;
	sram_mem[107650] = 16'b0000000000000000;
	sram_mem[107651] = 16'b0000000000000000;
	sram_mem[107652] = 16'b0000000000000000;
	sram_mem[107653] = 16'b0000000000000000;
	sram_mem[107654] = 16'b0000000000000000;
	sram_mem[107655] = 16'b0000000000000000;
	sram_mem[107656] = 16'b0000000000000000;
	sram_mem[107657] = 16'b0000000000000000;
	sram_mem[107658] = 16'b0000000000000000;
	sram_mem[107659] = 16'b0000000000000000;
	sram_mem[107660] = 16'b0000000000000000;
	sram_mem[107661] = 16'b0000000000000000;
	sram_mem[107662] = 16'b0000000000000000;
	sram_mem[107663] = 16'b0000000000000000;
	sram_mem[107664] = 16'b0000000000000000;
	sram_mem[107665] = 16'b0000000000000000;
	sram_mem[107666] = 16'b0000000000000000;
	sram_mem[107667] = 16'b0000000000000000;
	sram_mem[107668] = 16'b0000000000000000;
	sram_mem[107669] = 16'b0000000000000000;
	sram_mem[107670] = 16'b0000000000000000;
	sram_mem[107671] = 16'b0000000000000000;
	sram_mem[107672] = 16'b0000000000000000;
	sram_mem[107673] = 16'b0000000000000000;
	sram_mem[107674] = 16'b0000000000000000;
	sram_mem[107675] = 16'b0000000000000000;
	sram_mem[107676] = 16'b0000000000000000;
	sram_mem[107677] = 16'b0000000000000000;
	sram_mem[107678] = 16'b0000000000000000;
	sram_mem[107679] = 16'b0000000000000000;
	sram_mem[107680] = 16'b0000000000000000;
	sram_mem[107681] = 16'b0000000000000000;
	sram_mem[107682] = 16'b0000000000000000;
	sram_mem[107683] = 16'b0000000000000000;
	sram_mem[107684] = 16'b0000000000000000;
	sram_mem[107685] = 16'b0000000000000000;
	sram_mem[107686] = 16'b0000000000000000;
	sram_mem[107687] = 16'b0000000000000000;
	sram_mem[107688] = 16'b0000000000000000;
	sram_mem[107689] = 16'b0000000000000000;
	sram_mem[107690] = 16'b0000000000000000;
	sram_mem[107691] = 16'b0000000000000000;
	sram_mem[107692] = 16'b0000000000000000;
	sram_mem[107693] = 16'b0000000000000000;
	sram_mem[107694] = 16'b0000000000000000;
	sram_mem[107695] = 16'b0000000000000000;
	sram_mem[107696] = 16'b0000000000000000;
	sram_mem[107697] = 16'b0000000000000000;
	sram_mem[107698] = 16'b0000000000000000;
	sram_mem[107699] = 16'b0000000000000000;
	sram_mem[107700] = 16'b0000000000000000;
	sram_mem[107701] = 16'b0000000000000000;
	sram_mem[107702] = 16'b0000000000000000;
	sram_mem[107703] = 16'b0000000000000000;
	sram_mem[107704] = 16'b0000000000000000;
	sram_mem[107705] = 16'b0000000000000000;
	sram_mem[107706] = 16'b0000000000000000;
	sram_mem[107707] = 16'b0000000000000000;
	sram_mem[107708] = 16'b0000000000000000;
	sram_mem[107709] = 16'b0000000000000000;
	sram_mem[107710] = 16'b0000000000000000;
	sram_mem[107711] = 16'b0000000000000000;
	sram_mem[107712] = 16'b0000000000000000;
	sram_mem[107713] = 16'b0000000000000000;
	sram_mem[107714] = 16'b0000000000000000;
	sram_mem[107715] = 16'b0000000000000000;
	sram_mem[107716] = 16'b0000000000000000;
	sram_mem[107717] = 16'b0000000000000000;
	sram_mem[107718] = 16'b0000000000000000;
	sram_mem[107719] = 16'b0000000000000000;
	sram_mem[107720] = 16'b0000000000000000;
	sram_mem[107721] = 16'b0000000000000000;
	sram_mem[107722] = 16'b0000000000000000;
	sram_mem[107723] = 16'b0000000000000000;
	sram_mem[107724] = 16'b0000000000000000;
	sram_mem[107725] = 16'b0000000000000000;
	sram_mem[107726] = 16'b0000000000000000;
	sram_mem[107727] = 16'b0000000000000000;
	sram_mem[107728] = 16'b0000000000000000;
	sram_mem[107729] = 16'b0000000000000000;
	sram_mem[107730] = 16'b0000000000000000;
	sram_mem[107731] = 16'b0000000000000000;
	sram_mem[107732] = 16'b0000000000000000;
	sram_mem[107733] = 16'b0000000000000000;
	sram_mem[107734] = 16'b0000000000000000;
	sram_mem[107735] = 16'b0000000000000000;
	sram_mem[107736] = 16'b0000000000000000;
	sram_mem[107737] = 16'b0000000000000000;
	sram_mem[107738] = 16'b0000000000000000;
	sram_mem[107739] = 16'b0000000000000000;
	sram_mem[107740] = 16'b0000000000000000;
	sram_mem[107741] = 16'b0000000000000000;
	sram_mem[107742] = 16'b0000000000000000;
	sram_mem[107743] = 16'b0000000000000000;
	sram_mem[107744] = 16'b0000000000000000;
	sram_mem[107745] = 16'b0000000000000000;
	sram_mem[107746] = 16'b0000000000000000;
	sram_mem[107747] = 16'b0000000000000000;
	sram_mem[107748] = 16'b0000000000000000;
	sram_mem[107749] = 16'b0000000000000000;
	sram_mem[107750] = 16'b0000000000000000;
	sram_mem[107751] = 16'b0000000000000000;
	sram_mem[107752] = 16'b0000000000000000;
	sram_mem[107753] = 16'b0000000000000000;
	sram_mem[107754] = 16'b0000000000000000;
	sram_mem[107755] = 16'b0000000000000000;
	sram_mem[107756] = 16'b0000000000000000;
	sram_mem[107757] = 16'b0000000000000000;
	sram_mem[107758] = 16'b0000000000000000;
	sram_mem[107759] = 16'b0000000000000000;
	sram_mem[107760] = 16'b0000000000000000;
	sram_mem[107761] = 16'b0000000000000000;
	sram_mem[107762] = 16'b0000000000000000;
	sram_mem[107763] = 16'b0000000000000000;
	sram_mem[107764] = 16'b0000000000000000;
	sram_mem[107765] = 16'b0000000000000000;
	sram_mem[107766] = 16'b0000000000000000;
	sram_mem[107767] = 16'b0000000000000000;
	sram_mem[107768] = 16'b0000000000000000;
	sram_mem[107769] = 16'b0000000000000000;
	sram_mem[107770] = 16'b0000000000000000;
	sram_mem[107771] = 16'b0000000000000000;
	sram_mem[107772] = 16'b0000000000000000;
	sram_mem[107773] = 16'b0000000000000000;
	sram_mem[107774] = 16'b0000000000000000;
	sram_mem[107775] = 16'b0000000000000000;
	sram_mem[107776] = 16'b0000000000000000;
	sram_mem[107777] = 16'b0000000000000000;
	sram_mem[107778] = 16'b0000000000000000;
	sram_mem[107779] = 16'b0000000000000000;
	sram_mem[107780] = 16'b0000000000000000;
	sram_mem[107781] = 16'b0000000000000000;
	sram_mem[107782] = 16'b0000000000000000;
	sram_mem[107783] = 16'b0000000000000000;
	sram_mem[107784] = 16'b0000000000000000;
	sram_mem[107785] = 16'b0000000000000000;
	sram_mem[107786] = 16'b0000000000000000;
	sram_mem[107787] = 16'b0000000000000000;
	sram_mem[107788] = 16'b0000000000000000;
	sram_mem[107789] = 16'b0000000000000000;
	sram_mem[107790] = 16'b0000000000000000;
	sram_mem[107791] = 16'b0000000000000000;
	sram_mem[107792] = 16'b0000000000000000;
	sram_mem[107793] = 16'b0000000000000000;
	sram_mem[107794] = 16'b0000000000000000;
	sram_mem[107795] = 16'b0000000000000000;
	sram_mem[107796] = 16'b0000000000000000;
	sram_mem[107797] = 16'b0000000000000000;
	sram_mem[107798] = 16'b0000000000000000;
	sram_mem[107799] = 16'b0000000000000000;
	sram_mem[107800] = 16'b0000000000000000;
	sram_mem[107801] = 16'b0000000000000000;
	sram_mem[107802] = 16'b0000000000000000;
	sram_mem[107803] = 16'b0000000000000000;
	sram_mem[107804] = 16'b0000000000000000;
	sram_mem[107805] = 16'b0000000000000000;
	sram_mem[107806] = 16'b0000000000000000;
	sram_mem[107807] = 16'b0000000000000000;
	sram_mem[107808] = 16'b0000000000000000;
	sram_mem[107809] = 16'b0000000000000000;
	sram_mem[107810] = 16'b0000000000000000;
	sram_mem[107811] = 16'b0000000000000000;
	sram_mem[107812] = 16'b0000000000000000;
	sram_mem[107813] = 16'b0000000000000000;
	sram_mem[107814] = 16'b0000000000000000;
	sram_mem[107815] = 16'b0000000000000000;
	sram_mem[107816] = 16'b0000000000000000;
	sram_mem[107817] = 16'b0000000000000000;
	sram_mem[107818] = 16'b0000000000000000;
	sram_mem[107819] = 16'b0000000000000000;
	sram_mem[107820] = 16'b0000000000000000;
	sram_mem[107821] = 16'b0000000000000000;
	sram_mem[107822] = 16'b0000000000000000;
	sram_mem[107823] = 16'b0000000000000000;
	sram_mem[107824] = 16'b0000000000000000;
	sram_mem[107825] = 16'b0000000000000000;
	sram_mem[107826] = 16'b0000000000000000;
	sram_mem[107827] = 16'b0000000000000000;
	sram_mem[107828] = 16'b0000000000000000;
	sram_mem[107829] = 16'b0000000000000000;
	sram_mem[107830] = 16'b0000000000000000;
	sram_mem[107831] = 16'b0000000000000000;
	sram_mem[107832] = 16'b0000000000000000;
	sram_mem[107833] = 16'b0000000000000000;
	sram_mem[107834] = 16'b0000000000000000;
	sram_mem[107835] = 16'b0000000000000000;
	sram_mem[107836] = 16'b0000000000000000;
	sram_mem[107837] = 16'b0000000000000000;
	sram_mem[107838] = 16'b0000000000000000;
	sram_mem[107839] = 16'b0000000000000000;
	sram_mem[107840] = 16'b0000000000000000;
	sram_mem[107841] = 16'b0000000000000000;
	sram_mem[107842] = 16'b0000000000000000;
	sram_mem[107843] = 16'b0000000000000000;
	sram_mem[107844] = 16'b0000000000000000;
	sram_mem[107845] = 16'b0000000000000000;
	sram_mem[107846] = 16'b0000000000000000;
	sram_mem[107847] = 16'b0000000000000000;
	sram_mem[107848] = 16'b0000000000000000;
	sram_mem[107849] = 16'b0000000000000000;
	sram_mem[107850] = 16'b0000000000000000;
	sram_mem[107851] = 16'b0000000000000000;
	sram_mem[107852] = 16'b0000000000000000;
	sram_mem[107853] = 16'b0000000000000000;
	sram_mem[107854] = 16'b0000000000000000;
	sram_mem[107855] = 16'b0000000000000000;
	sram_mem[107856] = 16'b0000000000000000;
	sram_mem[107857] = 16'b0000000000000000;
	sram_mem[107858] = 16'b0000000000000000;
	sram_mem[107859] = 16'b0000000000000000;
	sram_mem[107860] = 16'b0000000000000000;
	sram_mem[107861] = 16'b0000000000000000;
	sram_mem[107862] = 16'b0000000000000000;
	sram_mem[107863] = 16'b0000000000000000;
	sram_mem[107864] = 16'b0000000000000000;
	sram_mem[107865] = 16'b0000000000000000;
	sram_mem[107866] = 16'b0000000000000000;
	sram_mem[107867] = 16'b0000000000000000;
	sram_mem[107868] = 16'b0000000000000000;
	sram_mem[107869] = 16'b0000000000000000;
	sram_mem[107870] = 16'b0000000000000000;
	sram_mem[107871] = 16'b0000000000000000;
	sram_mem[107872] = 16'b0000000000000000;
	sram_mem[107873] = 16'b0000000000000000;
	sram_mem[107874] = 16'b0000000000000000;
	sram_mem[107875] = 16'b0000000000000000;
	sram_mem[107876] = 16'b0000000000000000;
	sram_mem[107877] = 16'b0000000000000000;
	sram_mem[107878] = 16'b0000000000000000;
	sram_mem[107879] = 16'b0000000000000000;
	sram_mem[107880] = 16'b0000000000000000;
	sram_mem[107881] = 16'b0000000000000000;
	sram_mem[107882] = 16'b0000000000000000;
	sram_mem[107883] = 16'b0000000000000000;
	sram_mem[107884] = 16'b0000000000000000;
	sram_mem[107885] = 16'b0000000000000000;
	sram_mem[107886] = 16'b0000000000000000;
	sram_mem[107887] = 16'b0000000000000000;
	sram_mem[107888] = 16'b0000000000000000;
	sram_mem[107889] = 16'b0000000000000000;
	sram_mem[107890] = 16'b0000000000000000;
	sram_mem[107891] = 16'b0000000000000000;
	sram_mem[107892] = 16'b0000000000000000;
	sram_mem[107893] = 16'b0000000000000000;
	sram_mem[107894] = 16'b0000000000000000;
	sram_mem[107895] = 16'b0000000000000000;
	sram_mem[107896] = 16'b0000000000000000;
	sram_mem[107897] = 16'b0000000000000000;
	sram_mem[107898] = 16'b0000000000000000;
	sram_mem[107899] = 16'b0000000000000000;
	sram_mem[107900] = 16'b0000000000000000;
	sram_mem[107901] = 16'b0000000000000000;
	sram_mem[107902] = 16'b0000000000000000;
	sram_mem[107903] = 16'b0000000000000000;
	sram_mem[107904] = 16'b0000000000000000;
	sram_mem[107905] = 16'b0000000000000000;
	sram_mem[107906] = 16'b0000000000000000;
	sram_mem[107907] = 16'b0000000000000000;
	sram_mem[107908] = 16'b0000000000000000;
	sram_mem[107909] = 16'b0000000000000000;
	sram_mem[107910] = 16'b0000000000000000;
	sram_mem[107911] = 16'b0000000000000000;
	sram_mem[107912] = 16'b0000000000000000;
	sram_mem[107913] = 16'b0000000000000000;
	sram_mem[107914] = 16'b0000000000000000;
	sram_mem[107915] = 16'b0000000000000000;
	sram_mem[107916] = 16'b0000000000000000;
	sram_mem[107917] = 16'b0000000000000000;
	sram_mem[107918] = 16'b0000000000000000;
	sram_mem[107919] = 16'b0000000000000000;
	sram_mem[107920] = 16'b0000000000000000;
	sram_mem[107921] = 16'b0000000000000000;
	sram_mem[107922] = 16'b0000000000000000;
	sram_mem[107923] = 16'b0000000000000000;
	sram_mem[107924] = 16'b0000000000000000;
	sram_mem[107925] = 16'b0000000000000000;
	sram_mem[107926] = 16'b0000000000000000;
	sram_mem[107927] = 16'b0000000000000000;
	sram_mem[107928] = 16'b0000000000000000;
	sram_mem[107929] = 16'b0000000000000000;
	sram_mem[107930] = 16'b0000000000000000;
	sram_mem[107931] = 16'b0000000000000000;
	sram_mem[107932] = 16'b0000000000000000;
	sram_mem[107933] = 16'b0000000000000000;
	sram_mem[107934] = 16'b0000000000000000;
	sram_mem[107935] = 16'b0000000000000000;
	sram_mem[107936] = 16'b0000000000000000;
	sram_mem[107937] = 16'b0000000000000000;
	sram_mem[107938] = 16'b0000000000000000;
	sram_mem[107939] = 16'b0000000000000000;
	sram_mem[107940] = 16'b0000000000000000;
	sram_mem[107941] = 16'b0000000000000000;
	sram_mem[107942] = 16'b0000000000000000;
	sram_mem[107943] = 16'b0000000000000000;
	sram_mem[107944] = 16'b0000000000000000;
	sram_mem[107945] = 16'b0000000000000000;
	sram_mem[107946] = 16'b0000000000000000;
	sram_mem[107947] = 16'b0000000000000000;
	sram_mem[107948] = 16'b0000000000000000;
	sram_mem[107949] = 16'b0000000000000000;
	sram_mem[107950] = 16'b0000000000000000;
	sram_mem[107951] = 16'b0000000000000000;
	sram_mem[107952] = 16'b0000000000000000;
	sram_mem[107953] = 16'b0000000000000000;
	sram_mem[107954] = 16'b0000000000000000;
	sram_mem[107955] = 16'b0000000000000000;
	sram_mem[107956] = 16'b0000000000000000;
	sram_mem[107957] = 16'b0000000000000000;
	sram_mem[107958] = 16'b0000000000000000;
	sram_mem[107959] = 16'b0000000000000000;
	sram_mem[107960] = 16'b0000000000000000;
	sram_mem[107961] = 16'b0000000000000000;
	sram_mem[107962] = 16'b0000000000000000;
	sram_mem[107963] = 16'b0000000000000000;
	sram_mem[107964] = 16'b0000000000000000;
	sram_mem[107965] = 16'b0000000000000000;
	sram_mem[107966] = 16'b0000000000000000;
	sram_mem[107967] = 16'b0000000000000000;
	sram_mem[107968] = 16'b0000000000000000;
	sram_mem[107969] = 16'b0000000000000000;
	sram_mem[107970] = 16'b0000000000000000;
	sram_mem[107971] = 16'b0000000000000000;
	sram_mem[107972] = 16'b0000000000000000;
	sram_mem[107973] = 16'b0000000000000000;
	sram_mem[107974] = 16'b0000000000000000;
	sram_mem[107975] = 16'b0000000000000000;
	sram_mem[107976] = 16'b0000000000000000;
	sram_mem[107977] = 16'b0000000000000000;
	sram_mem[107978] = 16'b0000000000000000;
	sram_mem[107979] = 16'b0000000000000000;
	sram_mem[107980] = 16'b0000000000000000;
	sram_mem[107981] = 16'b0000000000000000;
	sram_mem[107982] = 16'b0000000000000000;
	sram_mem[107983] = 16'b0000000000000000;
	sram_mem[107984] = 16'b0000000000000000;
	sram_mem[107985] = 16'b0000000000000000;
	sram_mem[107986] = 16'b0000000000000000;
	sram_mem[107987] = 16'b0000000000000000;
	sram_mem[107988] = 16'b0000000000000000;
	sram_mem[107989] = 16'b0000000000000000;
	sram_mem[107990] = 16'b0000000000000000;
	sram_mem[107991] = 16'b0000000000000000;
	sram_mem[107992] = 16'b0000000000000000;
	sram_mem[107993] = 16'b0000000000000000;
	sram_mem[107994] = 16'b0000000000000000;
	sram_mem[107995] = 16'b0000000000000000;
	sram_mem[107996] = 16'b0000000000000000;
	sram_mem[107997] = 16'b0000000000000000;
	sram_mem[107998] = 16'b0000000000000000;
	sram_mem[107999] = 16'b0000000000000000;
	sram_mem[108000] = 16'b0000000000000000;
	sram_mem[108001] = 16'b0000000000000000;
	sram_mem[108002] = 16'b0000000000000000;
	sram_mem[108003] = 16'b0000000000000000;
	sram_mem[108004] = 16'b0000000000000000;
	sram_mem[108005] = 16'b0000000000000000;
	sram_mem[108006] = 16'b0000000000000000;
	sram_mem[108007] = 16'b0000000000000000;
	sram_mem[108008] = 16'b0000000000000000;
	sram_mem[108009] = 16'b0000000000000000;
	sram_mem[108010] = 16'b0000000000000000;
	sram_mem[108011] = 16'b0000000000000000;
	sram_mem[108012] = 16'b0000000000000000;
	sram_mem[108013] = 16'b0000000000000000;
	sram_mem[108014] = 16'b0000000000000000;
	sram_mem[108015] = 16'b0000000000000000;
	sram_mem[108016] = 16'b0000000000000000;
	sram_mem[108017] = 16'b0000000000000000;
	sram_mem[108018] = 16'b0000000000000000;
	sram_mem[108019] = 16'b0000000000000000;
	sram_mem[108020] = 16'b0000000000000000;
	sram_mem[108021] = 16'b0000000000000000;
	sram_mem[108022] = 16'b0000000000000000;
	sram_mem[108023] = 16'b0000000000000000;
	sram_mem[108024] = 16'b0000000000000000;
	sram_mem[108025] = 16'b0000000000000000;
	sram_mem[108026] = 16'b0000000000000000;
	sram_mem[108027] = 16'b0000000000000000;
	sram_mem[108028] = 16'b0000000000000000;
	sram_mem[108029] = 16'b0000000000000000;
	sram_mem[108030] = 16'b0000000000000000;
	sram_mem[108031] = 16'b0000000000000000;
	sram_mem[108032] = 16'b0000000000000000;
	sram_mem[108033] = 16'b0000000000000000;
	sram_mem[108034] = 16'b0000000000000000;
	sram_mem[108035] = 16'b0000000000000000;
	sram_mem[108036] = 16'b0000000000000000;
	sram_mem[108037] = 16'b0000000000000000;
	sram_mem[108038] = 16'b0000000000000000;
	sram_mem[108039] = 16'b0000000000000000;
	sram_mem[108040] = 16'b0000000000000000;
	sram_mem[108041] = 16'b0000000000000000;
	sram_mem[108042] = 16'b0000000000000000;
	sram_mem[108043] = 16'b0000000000000000;
	sram_mem[108044] = 16'b0000000000000000;
	sram_mem[108045] = 16'b0000000000000000;
	sram_mem[108046] = 16'b0000000000000000;
	sram_mem[108047] = 16'b0000000000000000;
	sram_mem[108048] = 16'b0000000000000000;
	sram_mem[108049] = 16'b0000000000000000;
	sram_mem[108050] = 16'b0000000000000000;
	sram_mem[108051] = 16'b0000000000000000;
	sram_mem[108052] = 16'b0000000000000000;
	sram_mem[108053] = 16'b0000000000000000;
	sram_mem[108054] = 16'b0000000000000000;
	sram_mem[108055] = 16'b0000000000000000;
	sram_mem[108056] = 16'b0000000000000000;
	sram_mem[108057] = 16'b0000000000000000;
	sram_mem[108058] = 16'b0000000000000000;
	sram_mem[108059] = 16'b0000000000000000;
	sram_mem[108060] = 16'b0000000000000000;
	sram_mem[108061] = 16'b0000000000000000;
	sram_mem[108062] = 16'b0000000000000000;
	sram_mem[108063] = 16'b0000000000000000;
	sram_mem[108064] = 16'b0000000000000000;
	sram_mem[108065] = 16'b0000000000000000;
	sram_mem[108066] = 16'b0000000000000000;
	sram_mem[108067] = 16'b0000000000000000;
	sram_mem[108068] = 16'b0000000000000000;
	sram_mem[108069] = 16'b0000000000000000;
	sram_mem[108070] = 16'b0000000000000000;
	sram_mem[108071] = 16'b0000000000000000;
	sram_mem[108072] = 16'b0000000000000000;
	sram_mem[108073] = 16'b0000000000000000;
	sram_mem[108074] = 16'b0000000000000000;
	sram_mem[108075] = 16'b0000000000000000;
	sram_mem[108076] = 16'b0000000000000000;
	sram_mem[108077] = 16'b0000000000000000;
	sram_mem[108078] = 16'b0000000000000000;
	sram_mem[108079] = 16'b0000000000000000;
	sram_mem[108080] = 16'b0000000000000000;
	sram_mem[108081] = 16'b0000000000000000;
	sram_mem[108082] = 16'b0000000000000000;
	sram_mem[108083] = 16'b0000000000000000;
	sram_mem[108084] = 16'b0000000000000000;
	sram_mem[108085] = 16'b0000000000000000;
	sram_mem[108086] = 16'b0000000000000000;
	sram_mem[108087] = 16'b0000000000000000;
	sram_mem[108088] = 16'b0000000000000000;
	sram_mem[108089] = 16'b0000000000000000;
	sram_mem[108090] = 16'b0000000000000000;
	sram_mem[108091] = 16'b0000000000000000;
	sram_mem[108092] = 16'b0000000000000000;
	sram_mem[108093] = 16'b0000000000000000;
	sram_mem[108094] = 16'b0000000000000000;
	sram_mem[108095] = 16'b0000000000000000;
	sram_mem[108096] = 16'b0000000000000000;
	sram_mem[108097] = 16'b0000000000000000;
	sram_mem[108098] = 16'b0000000000000000;
	sram_mem[108099] = 16'b0000000000000000;
	sram_mem[108100] = 16'b0000000000000000;
	sram_mem[108101] = 16'b0000000000000000;
	sram_mem[108102] = 16'b0000000000000000;
	sram_mem[108103] = 16'b0000000000000000;
	sram_mem[108104] = 16'b0000000000000000;
	sram_mem[108105] = 16'b0000000000000000;
	sram_mem[108106] = 16'b0000000000000000;
	sram_mem[108107] = 16'b0000000000000000;
	sram_mem[108108] = 16'b0000000000000000;
	sram_mem[108109] = 16'b0000000000000000;
	sram_mem[108110] = 16'b0000000000000000;
	sram_mem[108111] = 16'b0000000000000000;
	sram_mem[108112] = 16'b0000000000000000;
	sram_mem[108113] = 16'b0000000000000000;
	sram_mem[108114] = 16'b0000000000000000;
	sram_mem[108115] = 16'b0000000000000000;
	sram_mem[108116] = 16'b0000000000000000;
	sram_mem[108117] = 16'b0000000000000000;
	sram_mem[108118] = 16'b0000000000000000;
	sram_mem[108119] = 16'b0000000000000000;
	sram_mem[108120] = 16'b0000000000000000;
	sram_mem[108121] = 16'b0000000000000000;
	sram_mem[108122] = 16'b0000000000000000;
	sram_mem[108123] = 16'b0000000000000000;
	sram_mem[108124] = 16'b0000000000000000;
	sram_mem[108125] = 16'b0000000000000000;
	sram_mem[108126] = 16'b0000000000000000;
	sram_mem[108127] = 16'b0000000000000000;
	sram_mem[108128] = 16'b0000000000000000;
	sram_mem[108129] = 16'b0000000000000000;
	sram_mem[108130] = 16'b0000000000000000;
	sram_mem[108131] = 16'b0000000000000000;
	sram_mem[108132] = 16'b0000000000000000;
	sram_mem[108133] = 16'b0000000000000000;
	sram_mem[108134] = 16'b0000000000000000;
	sram_mem[108135] = 16'b0000000000000000;
	sram_mem[108136] = 16'b0000000000000000;
	sram_mem[108137] = 16'b0000000000000000;
	sram_mem[108138] = 16'b0000000000000000;
	sram_mem[108139] = 16'b0000000000000000;
	sram_mem[108140] = 16'b0000000000000000;
	sram_mem[108141] = 16'b0000000000000000;
	sram_mem[108142] = 16'b0000000000000000;
	sram_mem[108143] = 16'b0000000000000000;
	sram_mem[108144] = 16'b0000000000000000;
	sram_mem[108145] = 16'b0000000000000000;
	sram_mem[108146] = 16'b0000000000000000;
	sram_mem[108147] = 16'b0000000000000000;
	sram_mem[108148] = 16'b0000000000000000;
	sram_mem[108149] = 16'b0000000000000000;
	sram_mem[108150] = 16'b0000000000000000;
	sram_mem[108151] = 16'b0000000000000000;
	sram_mem[108152] = 16'b0000000000000000;
	sram_mem[108153] = 16'b0000000000000000;
	sram_mem[108154] = 16'b0000000000000000;
	sram_mem[108155] = 16'b0000000000000000;
	sram_mem[108156] = 16'b0000000000000000;
	sram_mem[108157] = 16'b0000000000000000;
	sram_mem[108158] = 16'b0000000000000000;
	sram_mem[108159] = 16'b0000000000000000;
	sram_mem[108160] = 16'b0000000000000000;
	sram_mem[108161] = 16'b0000000000000000;
	sram_mem[108162] = 16'b0000000000000000;
	sram_mem[108163] = 16'b0000000000000000;
	sram_mem[108164] = 16'b0000000000000000;
	sram_mem[108165] = 16'b0000000000000000;
	sram_mem[108166] = 16'b0000000000000000;
	sram_mem[108167] = 16'b0000000000000000;
	sram_mem[108168] = 16'b0000000000000000;
	sram_mem[108169] = 16'b0000000000000000;
	sram_mem[108170] = 16'b0000000000000000;
	sram_mem[108171] = 16'b0000000000000000;
	sram_mem[108172] = 16'b0000000000000000;
	sram_mem[108173] = 16'b0000000000000000;
	sram_mem[108174] = 16'b0000000000000000;
	sram_mem[108175] = 16'b0000000000000000;
	sram_mem[108176] = 16'b0000000000000000;
	sram_mem[108177] = 16'b0000000000000000;
	sram_mem[108178] = 16'b0000000000000000;
	sram_mem[108179] = 16'b0000000000000000;
	sram_mem[108180] = 16'b0000000000000000;
	sram_mem[108181] = 16'b0000000000000000;
	sram_mem[108182] = 16'b0000000000000000;
	sram_mem[108183] = 16'b0000000000000000;
	sram_mem[108184] = 16'b0000000000000000;
	sram_mem[108185] = 16'b0000000000000000;
	sram_mem[108186] = 16'b0000000000000000;
	sram_mem[108187] = 16'b0000000000000000;
	sram_mem[108188] = 16'b0000000000000000;
	sram_mem[108189] = 16'b0000000000000000;
	sram_mem[108190] = 16'b0000000000000000;
	sram_mem[108191] = 16'b0000000000000000;
	sram_mem[108192] = 16'b0000000000000000;
	sram_mem[108193] = 16'b0000000000000000;
	sram_mem[108194] = 16'b0000000000000000;
	sram_mem[108195] = 16'b0000000000000000;
	sram_mem[108196] = 16'b0000000000000000;
	sram_mem[108197] = 16'b0000000000000000;
	sram_mem[108198] = 16'b0000000000000000;
	sram_mem[108199] = 16'b0000000000000000;
	sram_mem[108200] = 16'b0000000000000000;
	sram_mem[108201] = 16'b0000000000000000;
	sram_mem[108202] = 16'b0000000000000000;
	sram_mem[108203] = 16'b0000000000000000;
	sram_mem[108204] = 16'b0000000000000000;
	sram_mem[108205] = 16'b0000000000000000;
	sram_mem[108206] = 16'b0000000000000000;
	sram_mem[108207] = 16'b0000000000000000;
	sram_mem[108208] = 16'b0000000000000000;
	sram_mem[108209] = 16'b0000000000000000;
	sram_mem[108210] = 16'b0000000000000000;
	sram_mem[108211] = 16'b0000000000000000;
	sram_mem[108212] = 16'b0000000000000000;
	sram_mem[108213] = 16'b0000000000000000;
	sram_mem[108214] = 16'b0000000000000000;
	sram_mem[108215] = 16'b0000000000000000;
	sram_mem[108216] = 16'b0000000000000000;
	sram_mem[108217] = 16'b0000000000000000;
	sram_mem[108218] = 16'b0000000000000000;
	sram_mem[108219] = 16'b0000000000000000;
	sram_mem[108220] = 16'b0000000000000000;
	sram_mem[108221] = 16'b0000000000000000;
	sram_mem[108222] = 16'b0000000000000000;
	sram_mem[108223] = 16'b0000000000000000;
	sram_mem[108224] = 16'b0000000000000000;
	sram_mem[108225] = 16'b0000000000000000;
	sram_mem[108226] = 16'b0000000000000000;
	sram_mem[108227] = 16'b0000000000000000;
	sram_mem[108228] = 16'b0000000000000000;
	sram_mem[108229] = 16'b0000000000000000;
	sram_mem[108230] = 16'b0000000000000000;
	sram_mem[108231] = 16'b0000000000000000;
	sram_mem[108232] = 16'b0000000000000000;
	sram_mem[108233] = 16'b0000000000000000;
	sram_mem[108234] = 16'b0000000000000000;
	sram_mem[108235] = 16'b0000000000000000;
	sram_mem[108236] = 16'b0000000000000000;
	sram_mem[108237] = 16'b0000000000000000;
	sram_mem[108238] = 16'b0000000000000000;
	sram_mem[108239] = 16'b0000000000000000;
	sram_mem[108240] = 16'b0000000000000000;
	sram_mem[108241] = 16'b0000000000000000;
	sram_mem[108242] = 16'b0000000000000000;
	sram_mem[108243] = 16'b0000000000000000;
	sram_mem[108244] = 16'b0000000000000000;
	sram_mem[108245] = 16'b0000000000000000;
	sram_mem[108246] = 16'b0000000000000000;
	sram_mem[108247] = 16'b0000000000000000;
	sram_mem[108248] = 16'b0000000000000000;
	sram_mem[108249] = 16'b0000000000000000;
	sram_mem[108250] = 16'b0000000000000000;
	sram_mem[108251] = 16'b0000000000000000;
	sram_mem[108252] = 16'b0000000000000000;
	sram_mem[108253] = 16'b0000000000000000;
	sram_mem[108254] = 16'b0000000000000000;
	sram_mem[108255] = 16'b0000000000000000;
	sram_mem[108256] = 16'b0000000000000000;
	sram_mem[108257] = 16'b0000000000000000;
	sram_mem[108258] = 16'b0000000000000000;
	sram_mem[108259] = 16'b0000000000000000;
	sram_mem[108260] = 16'b0000000000000000;
	sram_mem[108261] = 16'b0000000000000000;
	sram_mem[108262] = 16'b0000000000000000;
	sram_mem[108263] = 16'b0000000000000000;
	sram_mem[108264] = 16'b0000000000000000;
	sram_mem[108265] = 16'b0000000000000000;
	sram_mem[108266] = 16'b0000000000000000;
	sram_mem[108267] = 16'b0000000000000000;
	sram_mem[108268] = 16'b0000000000000000;
	sram_mem[108269] = 16'b0000000000000000;
	sram_mem[108270] = 16'b0000000000000000;
	sram_mem[108271] = 16'b0000000000000000;
	sram_mem[108272] = 16'b0000000000000000;
	sram_mem[108273] = 16'b0000000000000000;
	sram_mem[108274] = 16'b0000000000000000;
	sram_mem[108275] = 16'b0000000000000000;
	sram_mem[108276] = 16'b0000000000000000;
	sram_mem[108277] = 16'b0000000000000000;
	sram_mem[108278] = 16'b0000000000000000;
	sram_mem[108279] = 16'b0000000000000000;
	sram_mem[108280] = 16'b0000000000000000;
	sram_mem[108281] = 16'b0000000000000000;
	sram_mem[108282] = 16'b0000000000000000;
	sram_mem[108283] = 16'b0000000000000000;
	sram_mem[108284] = 16'b0000000000000000;
	sram_mem[108285] = 16'b0000000000000000;
	sram_mem[108286] = 16'b0000000000000000;
	sram_mem[108287] = 16'b0000000000000000;
	sram_mem[108288] = 16'b0000000000000000;
	sram_mem[108289] = 16'b0000000000000000;
	sram_mem[108290] = 16'b0000000000000000;
	sram_mem[108291] = 16'b0000000000000000;
	sram_mem[108292] = 16'b0000000000000000;
	sram_mem[108293] = 16'b0000000000000000;
	sram_mem[108294] = 16'b0000000000000000;
	sram_mem[108295] = 16'b0000000000000000;
	sram_mem[108296] = 16'b0000000000000000;
	sram_mem[108297] = 16'b0000000000000000;
	sram_mem[108298] = 16'b0000000000000000;
	sram_mem[108299] = 16'b0000000000000000;
	sram_mem[108300] = 16'b0000000000000000;
	sram_mem[108301] = 16'b0000000000000000;
	sram_mem[108302] = 16'b0000000000000000;
	sram_mem[108303] = 16'b0000000000000000;
	sram_mem[108304] = 16'b0000000000000000;
	sram_mem[108305] = 16'b0000000000000000;
	sram_mem[108306] = 16'b0000000000000000;
	sram_mem[108307] = 16'b0000000000000000;
	sram_mem[108308] = 16'b0000000000000000;
	sram_mem[108309] = 16'b0000000000000000;
	sram_mem[108310] = 16'b0000000000000000;
	sram_mem[108311] = 16'b0000000000000000;
	sram_mem[108312] = 16'b0000000000000000;
	sram_mem[108313] = 16'b0000000000000000;
	sram_mem[108314] = 16'b0000000000000000;
	sram_mem[108315] = 16'b0000000000000000;
	sram_mem[108316] = 16'b0000000000000000;
	sram_mem[108317] = 16'b0000000000000000;
	sram_mem[108318] = 16'b0000000000000000;
	sram_mem[108319] = 16'b0000000000000000;
	sram_mem[108320] = 16'b0000000000000000;
	sram_mem[108321] = 16'b0000000000000000;
	sram_mem[108322] = 16'b0000000000000000;
	sram_mem[108323] = 16'b0000000000000000;
	sram_mem[108324] = 16'b0000000000000000;
	sram_mem[108325] = 16'b0000000000000000;
	sram_mem[108326] = 16'b0000000000000000;
	sram_mem[108327] = 16'b0000000000000000;
	sram_mem[108328] = 16'b0000000000000000;
	sram_mem[108329] = 16'b0000000000000000;
	sram_mem[108330] = 16'b0000000000000000;
	sram_mem[108331] = 16'b0000000000000000;
	sram_mem[108332] = 16'b0000000000000000;
	sram_mem[108333] = 16'b0000000000000000;
	sram_mem[108334] = 16'b0000000000000000;
	sram_mem[108335] = 16'b0000000000000000;
	sram_mem[108336] = 16'b0000000000000000;
	sram_mem[108337] = 16'b0000000000000000;
	sram_mem[108338] = 16'b0000000000000000;
	sram_mem[108339] = 16'b0000000000000000;
	sram_mem[108340] = 16'b0000000000000000;
	sram_mem[108341] = 16'b0000000000000000;
	sram_mem[108342] = 16'b0000000000000000;
	sram_mem[108343] = 16'b0000000000000000;
	sram_mem[108344] = 16'b0000000000000000;
	sram_mem[108345] = 16'b0000000000000000;
	sram_mem[108346] = 16'b0000000000000000;
	sram_mem[108347] = 16'b0000000000000000;
	sram_mem[108348] = 16'b0000000000000000;
	sram_mem[108349] = 16'b0000000000000000;
	sram_mem[108350] = 16'b0000000000000000;
	sram_mem[108351] = 16'b0000000000000000;
	sram_mem[108352] = 16'b0000000000000000;
	sram_mem[108353] = 16'b0000000000000000;
	sram_mem[108354] = 16'b0000000000000000;
	sram_mem[108355] = 16'b0000000000000000;
	sram_mem[108356] = 16'b0000000000000000;
	sram_mem[108357] = 16'b0000000000000000;
	sram_mem[108358] = 16'b0000000000000000;
	sram_mem[108359] = 16'b0000000000000000;
	sram_mem[108360] = 16'b0000000000000000;
	sram_mem[108361] = 16'b0000000000000000;
	sram_mem[108362] = 16'b0000000000000000;
	sram_mem[108363] = 16'b0000000000000000;
	sram_mem[108364] = 16'b0000000000000000;
	sram_mem[108365] = 16'b0000000000000000;
	sram_mem[108366] = 16'b0000000000000000;
	sram_mem[108367] = 16'b0000000000000000;
	sram_mem[108368] = 16'b0000000000000000;
	sram_mem[108369] = 16'b0000000000000000;
	sram_mem[108370] = 16'b0000000000000000;
	sram_mem[108371] = 16'b0000000000000000;
	sram_mem[108372] = 16'b0000000000000000;
	sram_mem[108373] = 16'b0000000000000000;
	sram_mem[108374] = 16'b0000000000000000;
	sram_mem[108375] = 16'b0000000000000000;
	sram_mem[108376] = 16'b0000000000000000;
	sram_mem[108377] = 16'b0000000000000000;
	sram_mem[108378] = 16'b0000000000000000;
	sram_mem[108379] = 16'b0000000000000000;
	sram_mem[108380] = 16'b0000000000000000;
	sram_mem[108381] = 16'b0000000000000000;
	sram_mem[108382] = 16'b0000000000000000;
	sram_mem[108383] = 16'b0000000000000000;
	sram_mem[108384] = 16'b0000000000000000;
	sram_mem[108385] = 16'b0000000000000000;
	sram_mem[108386] = 16'b0000000000000000;
	sram_mem[108387] = 16'b0000000000000000;
	sram_mem[108388] = 16'b0000000000000000;
	sram_mem[108389] = 16'b0000000000000000;
	sram_mem[108390] = 16'b0000000000000000;
	sram_mem[108391] = 16'b0000000000000000;
	sram_mem[108392] = 16'b0000000000000000;
	sram_mem[108393] = 16'b0000000000000000;
	sram_mem[108394] = 16'b0000000000000000;
	sram_mem[108395] = 16'b0000000000000000;
	sram_mem[108396] = 16'b0000000000000000;
	sram_mem[108397] = 16'b0000000000000000;
	sram_mem[108398] = 16'b0000000000000000;
	sram_mem[108399] = 16'b0000000000000000;
	sram_mem[108400] = 16'b0000000000000000;
	sram_mem[108401] = 16'b0000000000000000;
	sram_mem[108402] = 16'b0000000000000000;
	sram_mem[108403] = 16'b0000000000000000;
	sram_mem[108404] = 16'b0000000000000000;
	sram_mem[108405] = 16'b0000000000000000;
	sram_mem[108406] = 16'b0000000000000000;
	sram_mem[108407] = 16'b0000000000000000;
	sram_mem[108408] = 16'b0000000000000000;
	sram_mem[108409] = 16'b0000000000000000;
	sram_mem[108410] = 16'b0000000000000000;
	sram_mem[108411] = 16'b0000000000000000;
	sram_mem[108412] = 16'b0000000000000000;
	sram_mem[108413] = 16'b0000000000000000;
	sram_mem[108414] = 16'b0000000000000000;
	sram_mem[108415] = 16'b0000000000000000;
	sram_mem[108416] = 16'b0000000000000000;
	sram_mem[108417] = 16'b0000000000000000;
	sram_mem[108418] = 16'b0000000000000000;
	sram_mem[108419] = 16'b0000000000000000;
	sram_mem[108420] = 16'b0000000000000000;
	sram_mem[108421] = 16'b0000000000000000;
	sram_mem[108422] = 16'b0000000000000000;
	sram_mem[108423] = 16'b0000000000000000;
	sram_mem[108424] = 16'b0000000000000000;
	sram_mem[108425] = 16'b0000000000000000;
	sram_mem[108426] = 16'b0000000000000000;
	sram_mem[108427] = 16'b0000000000000000;
	sram_mem[108428] = 16'b0000000000000000;
	sram_mem[108429] = 16'b0000000000000000;
	sram_mem[108430] = 16'b0000000000000000;
	sram_mem[108431] = 16'b0000000000000000;
	sram_mem[108432] = 16'b0000000000000000;
	sram_mem[108433] = 16'b0000000000000000;
	sram_mem[108434] = 16'b0000000000000000;
	sram_mem[108435] = 16'b0000000000000000;
	sram_mem[108436] = 16'b0000000000000000;
	sram_mem[108437] = 16'b0000000000000000;
	sram_mem[108438] = 16'b0000000000000000;
	sram_mem[108439] = 16'b0000000000000000;
	sram_mem[108440] = 16'b0000000000000000;
	sram_mem[108441] = 16'b0000000000000000;
	sram_mem[108442] = 16'b0000000000000000;
	sram_mem[108443] = 16'b0000000000000000;
	sram_mem[108444] = 16'b0000000000000000;
	sram_mem[108445] = 16'b0000000000000000;
	sram_mem[108446] = 16'b0000000000000000;
	sram_mem[108447] = 16'b0000000000000000;
	sram_mem[108448] = 16'b0000000000000000;
	sram_mem[108449] = 16'b0000000000000000;
	sram_mem[108450] = 16'b0000000000000000;
	sram_mem[108451] = 16'b0000000000000000;
	sram_mem[108452] = 16'b0000000000000000;
	sram_mem[108453] = 16'b0000000000000000;
	sram_mem[108454] = 16'b0000000000000000;
	sram_mem[108455] = 16'b0000000000000000;
	sram_mem[108456] = 16'b0000000000000000;
	sram_mem[108457] = 16'b0000000000000000;
	sram_mem[108458] = 16'b0000000000000000;
	sram_mem[108459] = 16'b0000000000000000;
	sram_mem[108460] = 16'b0000000000000000;
	sram_mem[108461] = 16'b0000000000000000;
	sram_mem[108462] = 16'b0000000000000000;
	sram_mem[108463] = 16'b0000000000000000;
	sram_mem[108464] = 16'b0000000000000000;
	sram_mem[108465] = 16'b0000000000000000;
	sram_mem[108466] = 16'b0000000000000000;
	sram_mem[108467] = 16'b0000000000000000;
	sram_mem[108468] = 16'b0000000000000000;
	sram_mem[108469] = 16'b0000000000000000;
	sram_mem[108470] = 16'b0000000000000000;
	sram_mem[108471] = 16'b0000000000000000;
	sram_mem[108472] = 16'b0000000000000000;
	sram_mem[108473] = 16'b0000000000000000;
	sram_mem[108474] = 16'b0000000000000000;
	sram_mem[108475] = 16'b0000000000000000;
	sram_mem[108476] = 16'b0000000000000000;
	sram_mem[108477] = 16'b0000000000000000;
	sram_mem[108478] = 16'b0000000000000000;
	sram_mem[108479] = 16'b0000000000000000;
	sram_mem[108480] = 16'b0000000000000000;
	sram_mem[108481] = 16'b0000000000000000;
	sram_mem[108482] = 16'b0000000000000000;
	sram_mem[108483] = 16'b0000000000000000;
	sram_mem[108484] = 16'b0000000000000000;
	sram_mem[108485] = 16'b0000000000000000;
	sram_mem[108486] = 16'b0000000000000000;
	sram_mem[108487] = 16'b0000000000000000;
	sram_mem[108488] = 16'b0000000000000000;
	sram_mem[108489] = 16'b0000000000000000;
	sram_mem[108490] = 16'b0000000000000000;
	sram_mem[108491] = 16'b0000000000000000;
	sram_mem[108492] = 16'b0000000000000000;
	sram_mem[108493] = 16'b0000000000000000;
	sram_mem[108494] = 16'b0000000000000000;
	sram_mem[108495] = 16'b0000000000000000;
	sram_mem[108496] = 16'b0000000000000000;
	sram_mem[108497] = 16'b0000000000000000;
	sram_mem[108498] = 16'b0000000000000000;
	sram_mem[108499] = 16'b0000000000000000;
	sram_mem[108500] = 16'b0000000000000000;
	sram_mem[108501] = 16'b0000000000000000;
	sram_mem[108502] = 16'b0000000000000000;
	sram_mem[108503] = 16'b0000000000000000;
	sram_mem[108504] = 16'b0000000000000000;
	sram_mem[108505] = 16'b0000000000000000;
	sram_mem[108506] = 16'b0000000000000000;
	sram_mem[108507] = 16'b0000000000000000;
	sram_mem[108508] = 16'b0000000000000000;
	sram_mem[108509] = 16'b0000000000000000;
	sram_mem[108510] = 16'b0000000000000000;
	sram_mem[108511] = 16'b0000000000000000;
	sram_mem[108512] = 16'b0000000000000000;
	sram_mem[108513] = 16'b0000000000000000;
	sram_mem[108514] = 16'b0000000000000000;
	sram_mem[108515] = 16'b0000000000000000;
	sram_mem[108516] = 16'b0000000000000000;
	sram_mem[108517] = 16'b0000000000000000;
	sram_mem[108518] = 16'b0000000000000000;
	sram_mem[108519] = 16'b0000000000000000;
	sram_mem[108520] = 16'b0000000000000000;
	sram_mem[108521] = 16'b0000000000000000;
	sram_mem[108522] = 16'b0000000000000000;
	sram_mem[108523] = 16'b0000000000000000;
	sram_mem[108524] = 16'b0000000000000000;
	sram_mem[108525] = 16'b0000000000000000;
	sram_mem[108526] = 16'b0000000000000000;
	sram_mem[108527] = 16'b0000000000000000;
	sram_mem[108528] = 16'b0000000000000000;
	sram_mem[108529] = 16'b0000000000000000;
	sram_mem[108530] = 16'b0000000000000000;
	sram_mem[108531] = 16'b0000000000000000;
	sram_mem[108532] = 16'b0000000000000000;
	sram_mem[108533] = 16'b0000000000000000;
	sram_mem[108534] = 16'b0000000000000000;
	sram_mem[108535] = 16'b0000000000000000;
	sram_mem[108536] = 16'b0000000000000000;
	sram_mem[108537] = 16'b0000000000000000;
	sram_mem[108538] = 16'b0000000000000000;
	sram_mem[108539] = 16'b0000000000000000;
	sram_mem[108540] = 16'b0000000000000000;
	sram_mem[108541] = 16'b0000000000000000;
	sram_mem[108542] = 16'b0000000000000000;
	sram_mem[108543] = 16'b0000000000000000;
	sram_mem[108544] = 16'b0000000000000000;
	sram_mem[108545] = 16'b0000000000000000;
	sram_mem[108546] = 16'b0000000000000000;
	sram_mem[108547] = 16'b0000000000000000;
	sram_mem[108548] = 16'b0000000000000000;
	sram_mem[108549] = 16'b0000000000000000;
	sram_mem[108550] = 16'b0000000000000000;
	sram_mem[108551] = 16'b0000000000000000;
	sram_mem[108552] = 16'b0000000000000000;
	sram_mem[108553] = 16'b0000000000000000;
	sram_mem[108554] = 16'b0000000000000000;
	sram_mem[108555] = 16'b0000000000000000;
	sram_mem[108556] = 16'b0000000000000000;
	sram_mem[108557] = 16'b0000000000000000;
	sram_mem[108558] = 16'b0000000000000000;
	sram_mem[108559] = 16'b0000000000000000;
	sram_mem[108560] = 16'b0000000000000000;
	sram_mem[108561] = 16'b0000000000000000;
	sram_mem[108562] = 16'b0000000000000000;
	sram_mem[108563] = 16'b0000000000000000;
	sram_mem[108564] = 16'b0000000000000000;
	sram_mem[108565] = 16'b0000000000000000;
	sram_mem[108566] = 16'b0000000000000000;
	sram_mem[108567] = 16'b0000000000000000;
	sram_mem[108568] = 16'b0000000000000000;
	sram_mem[108569] = 16'b0000000000000000;
	sram_mem[108570] = 16'b0000000000000000;
	sram_mem[108571] = 16'b0000000000000000;
	sram_mem[108572] = 16'b0000000000000000;
	sram_mem[108573] = 16'b0000000000000000;
	sram_mem[108574] = 16'b0000000000000000;
	sram_mem[108575] = 16'b0000000000000000;
	sram_mem[108576] = 16'b0000000000000000;
	sram_mem[108577] = 16'b0000000000000000;
	sram_mem[108578] = 16'b0000000000000000;
	sram_mem[108579] = 16'b0000000000000000;
	sram_mem[108580] = 16'b0000000000000000;
	sram_mem[108581] = 16'b0000000000000000;
	sram_mem[108582] = 16'b0000000000000000;
	sram_mem[108583] = 16'b0000000000000000;
	sram_mem[108584] = 16'b0000000000000000;
	sram_mem[108585] = 16'b0000000000000000;
	sram_mem[108586] = 16'b0000000000000000;
	sram_mem[108587] = 16'b0000000000000000;
	sram_mem[108588] = 16'b0000000000000000;
	sram_mem[108589] = 16'b0000000000000000;
	sram_mem[108590] = 16'b0000000000000000;
	sram_mem[108591] = 16'b0000000000000000;
	sram_mem[108592] = 16'b0000000000000000;
	sram_mem[108593] = 16'b0000000000000000;
	sram_mem[108594] = 16'b0000000000000000;
	sram_mem[108595] = 16'b0000000000000000;
	sram_mem[108596] = 16'b0000000000000000;
	sram_mem[108597] = 16'b0000000000000000;
	sram_mem[108598] = 16'b0000000000000000;
	sram_mem[108599] = 16'b0000000000000000;
	sram_mem[108600] = 16'b0000000000000000;
	sram_mem[108601] = 16'b0000000000000000;
	sram_mem[108602] = 16'b0000000000000000;
	sram_mem[108603] = 16'b0000000000000000;
	sram_mem[108604] = 16'b0000000000000000;
	sram_mem[108605] = 16'b0000000000000000;
	sram_mem[108606] = 16'b0000000000000000;
	sram_mem[108607] = 16'b0000000000000000;
	sram_mem[108608] = 16'b0000000000000000;
	sram_mem[108609] = 16'b0000000000000000;
	sram_mem[108610] = 16'b0000000000000000;
	sram_mem[108611] = 16'b0000000000000000;
	sram_mem[108612] = 16'b0000000000000000;
	sram_mem[108613] = 16'b0000000000000000;
	sram_mem[108614] = 16'b0000000000000000;
	sram_mem[108615] = 16'b0000000000000000;
	sram_mem[108616] = 16'b0000000000000000;
	sram_mem[108617] = 16'b0000000000000000;
	sram_mem[108618] = 16'b0000000000000000;
	sram_mem[108619] = 16'b0000000000000000;
	sram_mem[108620] = 16'b0000000000000000;
	sram_mem[108621] = 16'b0000000000000000;
	sram_mem[108622] = 16'b0000000000000000;
	sram_mem[108623] = 16'b0000000000000000;
	sram_mem[108624] = 16'b0000000000000000;
	sram_mem[108625] = 16'b0000000000000000;
	sram_mem[108626] = 16'b0000000000000000;
	sram_mem[108627] = 16'b0000000000000000;
	sram_mem[108628] = 16'b0000000000000000;
	sram_mem[108629] = 16'b0000000000000000;
	sram_mem[108630] = 16'b0000000000000000;
	sram_mem[108631] = 16'b0000000000000000;
	sram_mem[108632] = 16'b0000000000000000;
	sram_mem[108633] = 16'b0000000000000000;
	sram_mem[108634] = 16'b0000000000000000;
	sram_mem[108635] = 16'b0000000000000000;
	sram_mem[108636] = 16'b0000000000000000;
	sram_mem[108637] = 16'b0000000000000000;
	sram_mem[108638] = 16'b0000000000000000;
	sram_mem[108639] = 16'b0000000000000000;
	sram_mem[108640] = 16'b0000000000000000;
	sram_mem[108641] = 16'b0000000000000000;
	sram_mem[108642] = 16'b0000000000000000;
	sram_mem[108643] = 16'b0000000000000000;
	sram_mem[108644] = 16'b0000000000000000;
	sram_mem[108645] = 16'b0000000000000000;
	sram_mem[108646] = 16'b0000000000000000;
	sram_mem[108647] = 16'b0000000000000000;
	sram_mem[108648] = 16'b0000000000000000;
	sram_mem[108649] = 16'b0000000000000000;
	sram_mem[108650] = 16'b0000000000000000;
	sram_mem[108651] = 16'b0000000000000000;
	sram_mem[108652] = 16'b0000000000000000;
	sram_mem[108653] = 16'b0000000000000000;
	sram_mem[108654] = 16'b0000000000000000;
	sram_mem[108655] = 16'b0000000000000000;
	sram_mem[108656] = 16'b0000000000000000;
	sram_mem[108657] = 16'b0000000000000000;
	sram_mem[108658] = 16'b0000000000000000;
	sram_mem[108659] = 16'b0000000000000000;
	sram_mem[108660] = 16'b0000000000000000;
	sram_mem[108661] = 16'b0000000000000000;
	sram_mem[108662] = 16'b0000000000000000;
	sram_mem[108663] = 16'b0000000000000000;
	sram_mem[108664] = 16'b0000000000000000;
	sram_mem[108665] = 16'b0000000000000000;
	sram_mem[108666] = 16'b0000000000000000;
	sram_mem[108667] = 16'b0000000000000000;
	sram_mem[108668] = 16'b0000000000000000;
	sram_mem[108669] = 16'b0000000000000000;
	sram_mem[108670] = 16'b0000000000000000;
	sram_mem[108671] = 16'b0000000000000000;
	sram_mem[108672] = 16'b0000000000000000;
	sram_mem[108673] = 16'b0000000000000000;
	sram_mem[108674] = 16'b0000000000000000;
	sram_mem[108675] = 16'b0000000000000000;
	sram_mem[108676] = 16'b0000000000000000;
	sram_mem[108677] = 16'b0000000000000000;
	sram_mem[108678] = 16'b0000000000000000;
	sram_mem[108679] = 16'b0000000000000000;
	sram_mem[108680] = 16'b0000000000000000;
	sram_mem[108681] = 16'b0000000000000000;
	sram_mem[108682] = 16'b0000000000000000;
	sram_mem[108683] = 16'b0000000000000000;
	sram_mem[108684] = 16'b0000000000000000;
	sram_mem[108685] = 16'b0000000000000000;
	sram_mem[108686] = 16'b0000000000000000;
	sram_mem[108687] = 16'b0000000000000000;
	sram_mem[108688] = 16'b0000000000000000;
	sram_mem[108689] = 16'b0000000000000000;
	sram_mem[108690] = 16'b0000000000000000;
	sram_mem[108691] = 16'b0000000000000000;
	sram_mem[108692] = 16'b0000000000000000;
	sram_mem[108693] = 16'b0000000000000000;
	sram_mem[108694] = 16'b0000000000000000;
	sram_mem[108695] = 16'b0000000000000000;
	sram_mem[108696] = 16'b0000000000000000;
	sram_mem[108697] = 16'b0000000000000000;
	sram_mem[108698] = 16'b0000000000000000;
	sram_mem[108699] = 16'b0000000000000000;
	sram_mem[108700] = 16'b0000000000000000;
	sram_mem[108701] = 16'b0000000000000000;
	sram_mem[108702] = 16'b0000000000000000;
	sram_mem[108703] = 16'b0000000000000000;
	sram_mem[108704] = 16'b0000000000000000;
	sram_mem[108705] = 16'b0000000000000000;
	sram_mem[108706] = 16'b0000000000000000;
	sram_mem[108707] = 16'b0000000000000000;
	sram_mem[108708] = 16'b0000000000000000;
	sram_mem[108709] = 16'b0000000000000000;
	sram_mem[108710] = 16'b0000000000000000;
	sram_mem[108711] = 16'b0000000000000000;
	sram_mem[108712] = 16'b0000000000000000;
	sram_mem[108713] = 16'b0000000000000000;
	sram_mem[108714] = 16'b0000000000000000;
	sram_mem[108715] = 16'b0000000000000000;
	sram_mem[108716] = 16'b0000000000000000;
	sram_mem[108717] = 16'b0000000000000000;
	sram_mem[108718] = 16'b0000000000000000;
	sram_mem[108719] = 16'b0000000000000000;
	sram_mem[108720] = 16'b0000000000000000;
	sram_mem[108721] = 16'b0000000000000000;
	sram_mem[108722] = 16'b0000000000000000;
	sram_mem[108723] = 16'b0000000000000000;
	sram_mem[108724] = 16'b0000000000000000;
	sram_mem[108725] = 16'b0000000000000000;
	sram_mem[108726] = 16'b0000000000000000;
	sram_mem[108727] = 16'b0000000000000000;
	sram_mem[108728] = 16'b0000000000000000;
	sram_mem[108729] = 16'b0000000000000000;
	sram_mem[108730] = 16'b0000000000000000;
	sram_mem[108731] = 16'b0000000000000000;
	sram_mem[108732] = 16'b0000000000000000;
	sram_mem[108733] = 16'b0000000000000000;
	sram_mem[108734] = 16'b0000000000000000;
	sram_mem[108735] = 16'b0000000000000000;
	sram_mem[108736] = 16'b0000000000000000;
	sram_mem[108737] = 16'b0000000000000000;
	sram_mem[108738] = 16'b0000000000000000;
	sram_mem[108739] = 16'b0000000000000000;
	sram_mem[108740] = 16'b0000000000000000;
	sram_mem[108741] = 16'b0000000000000000;
	sram_mem[108742] = 16'b0000000000000000;
	sram_mem[108743] = 16'b0000000000000000;
	sram_mem[108744] = 16'b0000000000000000;
	sram_mem[108745] = 16'b0000000000000000;
	sram_mem[108746] = 16'b0000000000000000;
	sram_mem[108747] = 16'b0000000000000000;
	sram_mem[108748] = 16'b0000000000000000;
	sram_mem[108749] = 16'b0000000000000000;
	sram_mem[108750] = 16'b0000000000000000;
	sram_mem[108751] = 16'b0000000000000000;
	sram_mem[108752] = 16'b0000000000000000;
	sram_mem[108753] = 16'b0000000000000000;
	sram_mem[108754] = 16'b0000000000000000;
	sram_mem[108755] = 16'b0000000000000000;
	sram_mem[108756] = 16'b0000000000000000;
	sram_mem[108757] = 16'b0000000000000000;
	sram_mem[108758] = 16'b0000000000000000;
	sram_mem[108759] = 16'b0000000000000000;
	sram_mem[108760] = 16'b0000000000000000;
	sram_mem[108761] = 16'b0000000000000000;
	sram_mem[108762] = 16'b0000000000000000;
	sram_mem[108763] = 16'b0000000000000000;
	sram_mem[108764] = 16'b0000000000000000;
	sram_mem[108765] = 16'b0000000000000000;
	sram_mem[108766] = 16'b0000000000000000;
	sram_mem[108767] = 16'b0000000000000000;
	sram_mem[108768] = 16'b0000000000000000;
	sram_mem[108769] = 16'b0000000000000000;
	sram_mem[108770] = 16'b0000000000000000;
	sram_mem[108771] = 16'b0000000000000000;
	sram_mem[108772] = 16'b0000000000000000;
	sram_mem[108773] = 16'b0000000000000000;
	sram_mem[108774] = 16'b0000000000000000;
	sram_mem[108775] = 16'b0000000000000000;
	sram_mem[108776] = 16'b0000000000000000;
	sram_mem[108777] = 16'b0000000000000000;
	sram_mem[108778] = 16'b0000000000000000;
	sram_mem[108779] = 16'b0000000000000000;
	sram_mem[108780] = 16'b0000000000000000;
	sram_mem[108781] = 16'b0000000000000000;
	sram_mem[108782] = 16'b0000000000000000;
	sram_mem[108783] = 16'b0000000000000000;
	sram_mem[108784] = 16'b0000000000000000;
	sram_mem[108785] = 16'b0000000000000000;
	sram_mem[108786] = 16'b0000000000000000;
	sram_mem[108787] = 16'b0000000000000000;
	sram_mem[108788] = 16'b0000000000000000;
	sram_mem[108789] = 16'b0000000000000000;
	sram_mem[108790] = 16'b0000000000000000;
	sram_mem[108791] = 16'b0000000000000000;
	sram_mem[108792] = 16'b0000000000000000;
	sram_mem[108793] = 16'b0000000000000000;
	sram_mem[108794] = 16'b0000000000000000;
	sram_mem[108795] = 16'b0000000000000000;
	sram_mem[108796] = 16'b0000000000000000;
	sram_mem[108797] = 16'b0000000000000000;
	sram_mem[108798] = 16'b0000000000000000;
	sram_mem[108799] = 16'b0000000000000000;
	sram_mem[108800] = 16'b0000000000000000;
	sram_mem[108801] = 16'b0000000000000000;
	sram_mem[108802] = 16'b0000000000000000;
	sram_mem[108803] = 16'b0000000000000000;
	sram_mem[108804] = 16'b0000000000000000;
	sram_mem[108805] = 16'b0000000000000000;
	sram_mem[108806] = 16'b0000000000000000;
	sram_mem[108807] = 16'b0000000000000000;
	sram_mem[108808] = 16'b0000000000000000;
	sram_mem[108809] = 16'b0000000000000000;
	sram_mem[108810] = 16'b0000000000000000;
	sram_mem[108811] = 16'b0000000000000000;
	sram_mem[108812] = 16'b0000000000000000;
	sram_mem[108813] = 16'b0000000000000000;
	sram_mem[108814] = 16'b0000000000000000;
	sram_mem[108815] = 16'b0000000000000000;
	sram_mem[108816] = 16'b0000000000000000;
	sram_mem[108817] = 16'b0000000000000000;
	sram_mem[108818] = 16'b0000000000000000;
	sram_mem[108819] = 16'b0000000000000000;
	sram_mem[108820] = 16'b0000000000000000;
	sram_mem[108821] = 16'b0000000000000000;
	sram_mem[108822] = 16'b0000000000000000;
	sram_mem[108823] = 16'b0000000000000000;
	sram_mem[108824] = 16'b0000000000000000;
	sram_mem[108825] = 16'b0000000000000000;
	sram_mem[108826] = 16'b0000000000000000;
	sram_mem[108827] = 16'b0000000000000000;
	sram_mem[108828] = 16'b0000000000000000;
	sram_mem[108829] = 16'b0000000000000000;
	sram_mem[108830] = 16'b0000000000000000;
	sram_mem[108831] = 16'b0000000000000000;
	sram_mem[108832] = 16'b0000000000000000;
	sram_mem[108833] = 16'b0000000000000000;
	sram_mem[108834] = 16'b0000000000000000;
	sram_mem[108835] = 16'b0000000000000000;
	sram_mem[108836] = 16'b0000000000000000;
	sram_mem[108837] = 16'b0000000000000000;
	sram_mem[108838] = 16'b0000000000000000;
	sram_mem[108839] = 16'b0000000000000000;
	sram_mem[108840] = 16'b0000000000000000;
	sram_mem[108841] = 16'b0000000000000000;
	sram_mem[108842] = 16'b0000000000000000;
	sram_mem[108843] = 16'b0000000000000000;
	sram_mem[108844] = 16'b0000000000000000;
	sram_mem[108845] = 16'b0000000000000000;
	sram_mem[108846] = 16'b0000000000000000;
	sram_mem[108847] = 16'b0000000000000000;
	sram_mem[108848] = 16'b0000000000000000;
	sram_mem[108849] = 16'b0000000000000000;
	sram_mem[108850] = 16'b0000000000000000;
	sram_mem[108851] = 16'b0000000000000000;
	sram_mem[108852] = 16'b0000000000000000;
	sram_mem[108853] = 16'b0000000000000000;
	sram_mem[108854] = 16'b0000000000000000;
	sram_mem[108855] = 16'b0000000000000000;
	sram_mem[108856] = 16'b0000000000000000;
	sram_mem[108857] = 16'b0000000000000000;
	sram_mem[108858] = 16'b0000000000000000;
	sram_mem[108859] = 16'b0000000000000000;
	sram_mem[108860] = 16'b0000000000000000;
	sram_mem[108861] = 16'b0000000000000000;
	sram_mem[108862] = 16'b0000000000000000;
	sram_mem[108863] = 16'b0000000000000000;
	sram_mem[108864] = 16'b0000000000000000;
	sram_mem[108865] = 16'b0000000000000000;
	sram_mem[108866] = 16'b0000000000000000;
	sram_mem[108867] = 16'b0000000000000000;
	sram_mem[108868] = 16'b0000000000000000;
	sram_mem[108869] = 16'b0000000000000000;
	sram_mem[108870] = 16'b0000000000000000;
	sram_mem[108871] = 16'b0000000000000000;
	sram_mem[108872] = 16'b0000000000000000;
	sram_mem[108873] = 16'b0000000000000000;
	sram_mem[108874] = 16'b0000000000000000;
	sram_mem[108875] = 16'b0000000000000000;
	sram_mem[108876] = 16'b0000000000000000;
	sram_mem[108877] = 16'b0000000000000000;
	sram_mem[108878] = 16'b0000000000000000;
	sram_mem[108879] = 16'b0000000000000000;
	sram_mem[108880] = 16'b0000000000000000;
	sram_mem[108881] = 16'b0000000000000000;
	sram_mem[108882] = 16'b0000000000000000;
	sram_mem[108883] = 16'b0000000000000000;
	sram_mem[108884] = 16'b0000000000000000;
	sram_mem[108885] = 16'b0000000000000000;
	sram_mem[108886] = 16'b0000000000000000;
	sram_mem[108887] = 16'b0000000000000000;
	sram_mem[108888] = 16'b0000000000000000;
	sram_mem[108889] = 16'b0000000000000000;
	sram_mem[108890] = 16'b0000000000000000;
	sram_mem[108891] = 16'b0000000000000000;
	sram_mem[108892] = 16'b0000000000000000;
	sram_mem[108893] = 16'b0000000000000000;
	sram_mem[108894] = 16'b0000000000000000;
	sram_mem[108895] = 16'b0000000000000000;
	sram_mem[108896] = 16'b0000000000000000;
	sram_mem[108897] = 16'b0000000000000000;
	sram_mem[108898] = 16'b0000000000000000;
	sram_mem[108899] = 16'b0000000000000000;
	sram_mem[108900] = 16'b0000000000000000;
	sram_mem[108901] = 16'b0000000000000000;
	sram_mem[108902] = 16'b0000000000000000;
	sram_mem[108903] = 16'b0000000000000000;
	sram_mem[108904] = 16'b0000000000000000;
	sram_mem[108905] = 16'b0000000000000000;
	sram_mem[108906] = 16'b0000000000000000;
	sram_mem[108907] = 16'b0000000000000000;
	sram_mem[108908] = 16'b0000000000000000;
	sram_mem[108909] = 16'b0000000000000000;
	sram_mem[108910] = 16'b0000000000000000;
	sram_mem[108911] = 16'b0000000000000000;
	sram_mem[108912] = 16'b0000000000000000;
	sram_mem[108913] = 16'b0000000000000000;
	sram_mem[108914] = 16'b0000000000000000;
	sram_mem[108915] = 16'b0000000000000000;
	sram_mem[108916] = 16'b0000000000000000;
	sram_mem[108917] = 16'b0000000000000000;
	sram_mem[108918] = 16'b0000000000000000;
	sram_mem[108919] = 16'b0000000000000000;
	sram_mem[108920] = 16'b0000000000000000;
	sram_mem[108921] = 16'b0000000000000000;
	sram_mem[108922] = 16'b0000000000000000;
	sram_mem[108923] = 16'b0000000000000000;
	sram_mem[108924] = 16'b0000000000000000;
	sram_mem[108925] = 16'b0000000000000000;
	sram_mem[108926] = 16'b0000000000000000;
	sram_mem[108927] = 16'b0000000000000000;
	sram_mem[108928] = 16'b0000000000000000;
	sram_mem[108929] = 16'b0000000000000000;
	sram_mem[108930] = 16'b0000000000000000;
	sram_mem[108931] = 16'b0000000000000000;
	sram_mem[108932] = 16'b0000000000000000;
	sram_mem[108933] = 16'b0000000000000000;
	sram_mem[108934] = 16'b0000000000000000;
	sram_mem[108935] = 16'b0000000000000000;
	sram_mem[108936] = 16'b0000000000000000;
	sram_mem[108937] = 16'b0000000000000000;
	sram_mem[108938] = 16'b0000000000000000;
	sram_mem[108939] = 16'b0000000000000000;
	sram_mem[108940] = 16'b0000000000000000;
	sram_mem[108941] = 16'b0000000000000000;
	sram_mem[108942] = 16'b0000000000000000;
	sram_mem[108943] = 16'b0000000000000000;
	sram_mem[108944] = 16'b0000000000000000;
	sram_mem[108945] = 16'b0000000000000000;
	sram_mem[108946] = 16'b0000000000000000;
	sram_mem[108947] = 16'b0000000000000000;
	sram_mem[108948] = 16'b0000000000000000;
	sram_mem[108949] = 16'b0000000000000000;
	sram_mem[108950] = 16'b0000000000000000;
	sram_mem[108951] = 16'b0000000000000000;
	sram_mem[108952] = 16'b0000000000000000;
	sram_mem[108953] = 16'b0000000000000000;
	sram_mem[108954] = 16'b0000000000000000;
	sram_mem[108955] = 16'b0000000000000000;
	sram_mem[108956] = 16'b0000000000000000;
	sram_mem[108957] = 16'b0000000000000000;
	sram_mem[108958] = 16'b0000000000000000;
	sram_mem[108959] = 16'b0000000000000000;
	sram_mem[108960] = 16'b0000000000000000;
	sram_mem[108961] = 16'b0000000000000000;
	sram_mem[108962] = 16'b0000000000000000;
	sram_mem[108963] = 16'b0000000000000000;
	sram_mem[108964] = 16'b0000000000000000;
	sram_mem[108965] = 16'b0000000000000000;
	sram_mem[108966] = 16'b0000000000000000;
	sram_mem[108967] = 16'b0000000000000000;
	sram_mem[108968] = 16'b0000000000000000;
	sram_mem[108969] = 16'b0000000000000000;
	sram_mem[108970] = 16'b0000000000000000;
	sram_mem[108971] = 16'b0000000000000000;
	sram_mem[108972] = 16'b0000000000000000;
	sram_mem[108973] = 16'b0000000000000000;
	sram_mem[108974] = 16'b0000000000000000;
	sram_mem[108975] = 16'b0000000000000000;
	sram_mem[108976] = 16'b0000000000000000;
	sram_mem[108977] = 16'b0000000000000000;
	sram_mem[108978] = 16'b0000000000000000;
	sram_mem[108979] = 16'b0000000000000000;
	sram_mem[108980] = 16'b0000000000000000;
	sram_mem[108981] = 16'b0000000000000000;
	sram_mem[108982] = 16'b0000000000000000;
	sram_mem[108983] = 16'b0000000000000000;
	sram_mem[108984] = 16'b0000000000000000;
	sram_mem[108985] = 16'b0000000000000000;
	sram_mem[108986] = 16'b0000000000000000;
	sram_mem[108987] = 16'b0000000000000000;
	sram_mem[108988] = 16'b0000000000000000;
	sram_mem[108989] = 16'b0000000000000000;
	sram_mem[108990] = 16'b0000000000000000;
	sram_mem[108991] = 16'b0000000000000000;
	sram_mem[108992] = 16'b0000000000000000;
	sram_mem[108993] = 16'b0000000000000000;
	sram_mem[108994] = 16'b0000000000000000;
	sram_mem[108995] = 16'b0000000000000000;
	sram_mem[108996] = 16'b0000000000000000;
	sram_mem[108997] = 16'b0000000000000000;
	sram_mem[108998] = 16'b0000000000000000;
	sram_mem[108999] = 16'b0000000000000000;
	sram_mem[109000] = 16'b0000000000000000;
	sram_mem[109001] = 16'b0000000000000000;
	sram_mem[109002] = 16'b0000000000000000;
	sram_mem[109003] = 16'b0000000000000000;
	sram_mem[109004] = 16'b0000000000000000;
	sram_mem[109005] = 16'b0000000000000000;
	sram_mem[109006] = 16'b0000000000000000;
	sram_mem[109007] = 16'b0000000000000000;
	sram_mem[109008] = 16'b0000000000000000;
	sram_mem[109009] = 16'b0000000000000000;
	sram_mem[109010] = 16'b0000000000000000;
	sram_mem[109011] = 16'b0000000000000000;
	sram_mem[109012] = 16'b0000000000000000;
	sram_mem[109013] = 16'b0000000000000000;
	sram_mem[109014] = 16'b0000000000000000;
	sram_mem[109015] = 16'b0000000000000000;
	sram_mem[109016] = 16'b0000000000000000;
	sram_mem[109017] = 16'b0000000000000000;
	sram_mem[109018] = 16'b0000000000000000;
	sram_mem[109019] = 16'b0000000000000000;
	sram_mem[109020] = 16'b0000000000000000;
	sram_mem[109021] = 16'b0000000000000000;
	sram_mem[109022] = 16'b0000000000000000;
	sram_mem[109023] = 16'b0000000000000000;
	sram_mem[109024] = 16'b0000000000000000;
	sram_mem[109025] = 16'b0000000000000000;
	sram_mem[109026] = 16'b0000000000000000;
	sram_mem[109027] = 16'b0000000000000000;
	sram_mem[109028] = 16'b0000000000000000;
	sram_mem[109029] = 16'b0000000000000000;
	sram_mem[109030] = 16'b0000000000000000;
	sram_mem[109031] = 16'b0000000000000000;
	sram_mem[109032] = 16'b0000000000000000;
	sram_mem[109033] = 16'b0000000000000000;
	sram_mem[109034] = 16'b0000000000000000;
	sram_mem[109035] = 16'b0000000000000000;
	sram_mem[109036] = 16'b0000000000000000;
	sram_mem[109037] = 16'b0000000000000000;
	sram_mem[109038] = 16'b0000000000000000;
	sram_mem[109039] = 16'b0000000000000000;
	sram_mem[109040] = 16'b0000000000000000;
	sram_mem[109041] = 16'b0000000000000000;
	sram_mem[109042] = 16'b0000000000000000;
	sram_mem[109043] = 16'b0000000000000000;
	sram_mem[109044] = 16'b0000000000000000;
	sram_mem[109045] = 16'b0000000000000000;
	sram_mem[109046] = 16'b0000000000000000;
	sram_mem[109047] = 16'b0000000000000000;
	sram_mem[109048] = 16'b0000000000000000;
	sram_mem[109049] = 16'b0000000000000000;
	sram_mem[109050] = 16'b0000000000000000;
	sram_mem[109051] = 16'b0000000000000000;
	sram_mem[109052] = 16'b0000000000000000;
	sram_mem[109053] = 16'b0000000000000000;
	sram_mem[109054] = 16'b0000000000000000;
	sram_mem[109055] = 16'b0000000000000000;
	sram_mem[109056] = 16'b0000000000000000;
	sram_mem[109057] = 16'b0000000000000000;
	sram_mem[109058] = 16'b0000000000000000;
	sram_mem[109059] = 16'b0000000000000000;
	sram_mem[109060] = 16'b0000000000000000;
	sram_mem[109061] = 16'b0000000000000000;
	sram_mem[109062] = 16'b0000000000000000;
	sram_mem[109063] = 16'b0000000000000000;
	sram_mem[109064] = 16'b0000000000000000;
	sram_mem[109065] = 16'b0000000000000000;
	sram_mem[109066] = 16'b0000000000000000;
	sram_mem[109067] = 16'b0000000000000000;
	sram_mem[109068] = 16'b0000000000000000;
	sram_mem[109069] = 16'b0000000000000000;
	sram_mem[109070] = 16'b0000000000000000;
	sram_mem[109071] = 16'b0000000000000000;
	sram_mem[109072] = 16'b0000000000000000;
	sram_mem[109073] = 16'b0000000000000000;
	sram_mem[109074] = 16'b0000000000000000;
	sram_mem[109075] = 16'b0000000000000000;
	sram_mem[109076] = 16'b0000000000000000;
	sram_mem[109077] = 16'b0000000000000000;
	sram_mem[109078] = 16'b0000000000000000;
	sram_mem[109079] = 16'b0000000000000000;
	sram_mem[109080] = 16'b0000000000000000;
	sram_mem[109081] = 16'b0000000000000000;
	sram_mem[109082] = 16'b0000000000000000;
	sram_mem[109083] = 16'b0000000000000000;
	sram_mem[109084] = 16'b0000000000000000;
	sram_mem[109085] = 16'b0000000000000000;
	sram_mem[109086] = 16'b0000000000000000;
	sram_mem[109087] = 16'b0000000000000000;
	sram_mem[109088] = 16'b0000000000000000;
	sram_mem[109089] = 16'b0000000000000000;
	sram_mem[109090] = 16'b0000000000000000;
	sram_mem[109091] = 16'b0000000000000000;
	sram_mem[109092] = 16'b0000000000000000;
	sram_mem[109093] = 16'b0000000000000000;
	sram_mem[109094] = 16'b0000000000000000;
	sram_mem[109095] = 16'b0000000000000000;
	sram_mem[109096] = 16'b0000000000000000;
	sram_mem[109097] = 16'b0000000000000000;
	sram_mem[109098] = 16'b0000000000000000;
	sram_mem[109099] = 16'b0000000000000000;
	sram_mem[109100] = 16'b0000000000000000;
	sram_mem[109101] = 16'b0000000000000000;
	sram_mem[109102] = 16'b0000000000000000;
	sram_mem[109103] = 16'b0000000000000000;
	sram_mem[109104] = 16'b0000000000000000;
	sram_mem[109105] = 16'b0000000000000000;
	sram_mem[109106] = 16'b0000000000000000;
	sram_mem[109107] = 16'b0000000000000000;
	sram_mem[109108] = 16'b0000000000000000;
	sram_mem[109109] = 16'b0000000000000000;
	sram_mem[109110] = 16'b0000000000000000;
	sram_mem[109111] = 16'b0000000000000000;
	sram_mem[109112] = 16'b0000000000000000;
	sram_mem[109113] = 16'b0000000000000000;
	sram_mem[109114] = 16'b0000000000000000;
	sram_mem[109115] = 16'b0000000000000000;
	sram_mem[109116] = 16'b0000000000000000;
	sram_mem[109117] = 16'b0000000000000000;
	sram_mem[109118] = 16'b0000000000000000;
	sram_mem[109119] = 16'b0000000000000000;
	sram_mem[109120] = 16'b0000000000000000;
	sram_mem[109121] = 16'b0000000000000000;
	sram_mem[109122] = 16'b0000000000000000;
	sram_mem[109123] = 16'b0000000000000000;
	sram_mem[109124] = 16'b0000000000000000;
	sram_mem[109125] = 16'b0000000000000000;
	sram_mem[109126] = 16'b0000000000000000;
	sram_mem[109127] = 16'b0000000000000000;
	sram_mem[109128] = 16'b0000000000000000;
	sram_mem[109129] = 16'b0000000000000000;
	sram_mem[109130] = 16'b0000000000000000;
	sram_mem[109131] = 16'b0000000000000000;
	sram_mem[109132] = 16'b0000000000000000;
	sram_mem[109133] = 16'b0000000000000000;
	sram_mem[109134] = 16'b0000000000000000;
	sram_mem[109135] = 16'b0000000000000000;
	sram_mem[109136] = 16'b0000000000000000;
	sram_mem[109137] = 16'b0000000000000000;
	sram_mem[109138] = 16'b0000000000000000;
	sram_mem[109139] = 16'b0000000000000000;
	sram_mem[109140] = 16'b0000000000000000;
	sram_mem[109141] = 16'b0000000000000000;
	sram_mem[109142] = 16'b0000000000000000;
	sram_mem[109143] = 16'b0000000000000000;
	sram_mem[109144] = 16'b0000000000000000;
	sram_mem[109145] = 16'b0000000000000000;
	sram_mem[109146] = 16'b0000000000000000;
	sram_mem[109147] = 16'b0000000000000000;
	sram_mem[109148] = 16'b0000000000000000;
	sram_mem[109149] = 16'b0000000000000000;
	sram_mem[109150] = 16'b0000000000000000;
	sram_mem[109151] = 16'b0000000000000000;
	sram_mem[109152] = 16'b0000000000000000;
	sram_mem[109153] = 16'b0000000000000000;
	sram_mem[109154] = 16'b0000000000000000;
	sram_mem[109155] = 16'b0000000000000000;
	sram_mem[109156] = 16'b0000000000000000;
	sram_mem[109157] = 16'b0000000000000000;
	sram_mem[109158] = 16'b0000000000000000;
	sram_mem[109159] = 16'b0000000000000000;
	sram_mem[109160] = 16'b0000000000000000;
	sram_mem[109161] = 16'b0000000000000000;
	sram_mem[109162] = 16'b0000000000000000;
	sram_mem[109163] = 16'b0000000000000000;
	sram_mem[109164] = 16'b0000000000000000;
	sram_mem[109165] = 16'b0000000000000000;
	sram_mem[109166] = 16'b0000000000000000;
	sram_mem[109167] = 16'b0000000000000000;
	sram_mem[109168] = 16'b0000000000000000;
	sram_mem[109169] = 16'b0000000000000000;
	sram_mem[109170] = 16'b0000000000000000;
	sram_mem[109171] = 16'b0000000000000000;
	sram_mem[109172] = 16'b0000000000000000;
	sram_mem[109173] = 16'b0000000000000000;
	sram_mem[109174] = 16'b0000000000000000;
	sram_mem[109175] = 16'b0000000000000000;
	sram_mem[109176] = 16'b0000000000000000;
	sram_mem[109177] = 16'b0000000000000000;
	sram_mem[109178] = 16'b0000000000000000;
	sram_mem[109179] = 16'b0000000000000000;
	sram_mem[109180] = 16'b0000000000000000;
	sram_mem[109181] = 16'b0000000000000000;
	sram_mem[109182] = 16'b0000000000000000;
	sram_mem[109183] = 16'b0000000000000000;
	sram_mem[109184] = 16'b0000000000000000;
	sram_mem[109185] = 16'b0000000000000000;
	sram_mem[109186] = 16'b0000000000000000;
	sram_mem[109187] = 16'b0000000000000000;
	sram_mem[109188] = 16'b0000000000000000;
	sram_mem[109189] = 16'b0000000000000000;
	sram_mem[109190] = 16'b0000000000000000;
	sram_mem[109191] = 16'b0000000000000000;
	sram_mem[109192] = 16'b0000000000000000;
	sram_mem[109193] = 16'b0000000000000000;
	sram_mem[109194] = 16'b0000000000000000;
	sram_mem[109195] = 16'b0000000000000000;
	sram_mem[109196] = 16'b0000000000000000;
	sram_mem[109197] = 16'b0000000000000000;
	sram_mem[109198] = 16'b0000000000000000;
	sram_mem[109199] = 16'b0000000000000000;
	sram_mem[109200] = 16'b0000000000000000;
	sram_mem[109201] = 16'b0000000000000000;
	sram_mem[109202] = 16'b0000000000000000;
	sram_mem[109203] = 16'b0000000000000000;
	sram_mem[109204] = 16'b0000000000000000;
	sram_mem[109205] = 16'b0000000000000000;
	sram_mem[109206] = 16'b0000000000000000;
	sram_mem[109207] = 16'b0000000000000000;
	sram_mem[109208] = 16'b0000000000000000;
	sram_mem[109209] = 16'b0000000000000000;
	sram_mem[109210] = 16'b0000000000000000;
	sram_mem[109211] = 16'b0000000000000000;
	sram_mem[109212] = 16'b0000000000000000;
	sram_mem[109213] = 16'b0000000000000000;
	sram_mem[109214] = 16'b0000000000000000;
	sram_mem[109215] = 16'b0000000000000000;
	sram_mem[109216] = 16'b0000000000000000;
	sram_mem[109217] = 16'b0000000000000000;
	sram_mem[109218] = 16'b0000000000000000;
	sram_mem[109219] = 16'b0000000000000000;
	sram_mem[109220] = 16'b0000000000000000;
	sram_mem[109221] = 16'b0000000000000000;
	sram_mem[109222] = 16'b0000000000000000;
	sram_mem[109223] = 16'b0000000000000000;
	sram_mem[109224] = 16'b0000000000000000;
	sram_mem[109225] = 16'b0000000000000000;
	sram_mem[109226] = 16'b0000000000000000;
	sram_mem[109227] = 16'b0000000000000000;
	sram_mem[109228] = 16'b0000000000000000;
	sram_mem[109229] = 16'b0000000000000000;
	sram_mem[109230] = 16'b0000000000000000;
	sram_mem[109231] = 16'b0000000000000000;
	sram_mem[109232] = 16'b0000000000000000;
	sram_mem[109233] = 16'b0000000000000000;
	sram_mem[109234] = 16'b0000000000000000;
	sram_mem[109235] = 16'b0000000000000000;
	sram_mem[109236] = 16'b0000000000000000;
	sram_mem[109237] = 16'b0000000000000000;
	sram_mem[109238] = 16'b0000000000000000;
	sram_mem[109239] = 16'b0000000000000000;
	sram_mem[109240] = 16'b0000000000000000;
	sram_mem[109241] = 16'b0000000000000000;
	sram_mem[109242] = 16'b0000000000000000;
	sram_mem[109243] = 16'b0000000000000000;
	sram_mem[109244] = 16'b0000000000000000;
	sram_mem[109245] = 16'b0000000000000000;
	sram_mem[109246] = 16'b0000000000000000;
	sram_mem[109247] = 16'b0000000000000000;
	sram_mem[109248] = 16'b0000000000000000;
	sram_mem[109249] = 16'b0000000000000000;
	sram_mem[109250] = 16'b0000000000000000;
	sram_mem[109251] = 16'b0000000000000000;
	sram_mem[109252] = 16'b0000000000000000;
	sram_mem[109253] = 16'b0000000000000000;
	sram_mem[109254] = 16'b0000000000000000;
	sram_mem[109255] = 16'b0000000000000000;
	sram_mem[109256] = 16'b0000000000000000;
	sram_mem[109257] = 16'b0000000000000000;
	sram_mem[109258] = 16'b0000000000000000;
	sram_mem[109259] = 16'b0000000000000000;
	sram_mem[109260] = 16'b0000000000000000;
	sram_mem[109261] = 16'b0000000000000000;
	sram_mem[109262] = 16'b0000000000000000;
	sram_mem[109263] = 16'b0000000000000000;
	sram_mem[109264] = 16'b0000000000000000;
	sram_mem[109265] = 16'b0000000000000000;
	sram_mem[109266] = 16'b0000000000000000;
	sram_mem[109267] = 16'b0000000000000000;
	sram_mem[109268] = 16'b0000000000000000;
	sram_mem[109269] = 16'b0000000000000000;
	sram_mem[109270] = 16'b0000000000000000;
	sram_mem[109271] = 16'b0000000000000000;
	sram_mem[109272] = 16'b0000000000000000;
	sram_mem[109273] = 16'b0000000000000000;
	sram_mem[109274] = 16'b0000000000000000;
	sram_mem[109275] = 16'b0000000000000000;
	sram_mem[109276] = 16'b0000000000000000;
	sram_mem[109277] = 16'b0000000000000000;
	sram_mem[109278] = 16'b0000000000000000;
	sram_mem[109279] = 16'b0000000000000000;
	sram_mem[109280] = 16'b0000000000000000;
	sram_mem[109281] = 16'b0000000000000000;
	sram_mem[109282] = 16'b0000000000000000;
	sram_mem[109283] = 16'b0000000000000000;
	sram_mem[109284] = 16'b0000000000000000;
	sram_mem[109285] = 16'b0000000000000000;
	sram_mem[109286] = 16'b0000000000000000;
	sram_mem[109287] = 16'b0000000000000000;
	sram_mem[109288] = 16'b0000000000000000;
	sram_mem[109289] = 16'b0000000000000000;
	sram_mem[109290] = 16'b0000000000000000;
	sram_mem[109291] = 16'b0000000000000000;
	sram_mem[109292] = 16'b0000000000000000;
	sram_mem[109293] = 16'b0000000000000000;
	sram_mem[109294] = 16'b0000000000000000;
	sram_mem[109295] = 16'b0000000000000000;
	sram_mem[109296] = 16'b0000000000000000;
	sram_mem[109297] = 16'b0000000000000000;
	sram_mem[109298] = 16'b0000000000000000;
	sram_mem[109299] = 16'b0000000000000000;
	sram_mem[109300] = 16'b0000000000000000;
	sram_mem[109301] = 16'b0000000000000000;
	sram_mem[109302] = 16'b0000000000000000;
	sram_mem[109303] = 16'b0000000000000000;
	sram_mem[109304] = 16'b0000000000000000;
	sram_mem[109305] = 16'b0000000000000000;
	sram_mem[109306] = 16'b0000000000000000;
	sram_mem[109307] = 16'b0000000000000000;
	sram_mem[109308] = 16'b0000000000000000;
	sram_mem[109309] = 16'b0000000000000000;
	sram_mem[109310] = 16'b0000000000000000;
	sram_mem[109311] = 16'b0000000000000000;
	sram_mem[109312] = 16'b0000000000000000;
	sram_mem[109313] = 16'b0000000000000000;
	sram_mem[109314] = 16'b0000000000000000;
	sram_mem[109315] = 16'b0000000000000000;
	sram_mem[109316] = 16'b0000000000000000;
	sram_mem[109317] = 16'b0000000000000000;
	sram_mem[109318] = 16'b0000000000000000;
	sram_mem[109319] = 16'b0000000000000000;
	sram_mem[109320] = 16'b0000000000000000;
	sram_mem[109321] = 16'b0000000000000000;
	sram_mem[109322] = 16'b0000000000000000;
	sram_mem[109323] = 16'b0000000000000000;
	sram_mem[109324] = 16'b0000000000000000;
	sram_mem[109325] = 16'b0000000000000000;
	sram_mem[109326] = 16'b0000000000000000;
	sram_mem[109327] = 16'b0000000000000000;
	sram_mem[109328] = 16'b0000000000000000;
	sram_mem[109329] = 16'b0000000000000000;
	sram_mem[109330] = 16'b0000000000000000;
	sram_mem[109331] = 16'b0000000000000000;
	sram_mem[109332] = 16'b0000000000000000;
	sram_mem[109333] = 16'b0000000000000000;
	sram_mem[109334] = 16'b0000000000000000;
	sram_mem[109335] = 16'b0000000000000000;
	sram_mem[109336] = 16'b0000000000000000;
	sram_mem[109337] = 16'b0000000000000000;
	sram_mem[109338] = 16'b0000000000000000;
	sram_mem[109339] = 16'b0000000000000000;
	sram_mem[109340] = 16'b0000000000000000;
	sram_mem[109341] = 16'b0000000000000000;
	sram_mem[109342] = 16'b0000000000000000;
	sram_mem[109343] = 16'b0000000000000000;
	sram_mem[109344] = 16'b0000000000000000;
	sram_mem[109345] = 16'b0000000000000000;
	sram_mem[109346] = 16'b0000000000000000;
	sram_mem[109347] = 16'b0000000000000000;
	sram_mem[109348] = 16'b0000000000000000;
	sram_mem[109349] = 16'b0000000000000000;
	sram_mem[109350] = 16'b0000000000000000;
	sram_mem[109351] = 16'b0000000000000000;
	sram_mem[109352] = 16'b0000000000000000;
	sram_mem[109353] = 16'b0000000000000000;
	sram_mem[109354] = 16'b0000000000000000;
	sram_mem[109355] = 16'b0000000000000000;
	sram_mem[109356] = 16'b0000000000000000;
	sram_mem[109357] = 16'b0000000000000000;
	sram_mem[109358] = 16'b0000000000000000;
	sram_mem[109359] = 16'b0000000000000000;
	sram_mem[109360] = 16'b0000000000000000;
	sram_mem[109361] = 16'b0000000000000000;
	sram_mem[109362] = 16'b0000000000000000;
	sram_mem[109363] = 16'b0000000000000000;
	sram_mem[109364] = 16'b0000000000000000;
	sram_mem[109365] = 16'b0000000000000000;
	sram_mem[109366] = 16'b0000000000000000;
	sram_mem[109367] = 16'b0000000000000000;
	sram_mem[109368] = 16'b0000000000000000;
	sram_mem[109369] = 16'b0000000000000000;
	sram_mem[109370] = 16'b0000000000000000;
	sram_mem[109371] = 16'b0000000000000000;
	sram_mem[109372] = 16'b0000000000000000;
	sram_mem[109373] = 16'b0000000000000000;
	sram_mem[109374] = 16'b0000000000000000;
	sram_mem[109375] = 16'b0000000000000000;
	sram_mem[109376] = 16'b0000000000000000;
	sram_mem[109377] = 16'b0000000000000000;
	sram_mem[109378] = 16'b0000000000000000;
	sram_mem[109379] = 16'b0000000000000000;
	sram_mem[109380] = 16'b0000000000000000;
	sram_mem[109381] = 16'b0000000000000000;
	sram_mem[109382] = 16'b0000000000000000;
	sram_mem[109383] = 16'b0000000000000000;
	sram_mem[109384] = 16'b0000000000000000;
	sram_mem[109385] = 16'b0000000000000000;
	sram_mem[109386] = 16'b0000000000000000;
	sram_mem[109387] = 16'b0000000000000000;
	sram_mem[109388] = 16'b0000000000000000;
	sram_mem[109389] = 16'b0000000000000000;
	sram_mem[109390] = 16'b0000000000000000;
	sram_mem[109391] = 16'b0000000000000000;
	sram_mem[109392] = 16'b0000000000000000;
	sram_mem[109393] = 16'b0000000000000000;
	sram_mem[109394] = 16'b0000000000000000;
	sram_mem[109395] = 16'b0000000000000000;
	sram_mem[109396] = 16'b0000000000000000;
	sram_mem[109397] = 16'b0000000000000000;
	sram_mem[109398] = 16'b0000000000000000;
	sram_mem[109399] = 16'b0000000000000000;
	sram_mem[109400] = 16'b0000000000000000;
	sram_mem[109401] = 16'b0000000000000000;
	sram_mem[109402] = 16'b0000000000000000;
	sram_mem[109403] = 16'b0000000000000000;
	sram_mem[109404] = 16'b0000000000000000;
	sram_mem[109405] = 16'b0000000000000000;
	sram_mem[109406] = 16'b0000000000000000;
	sram_mem[109407] = 16'b0000000000000000;
	sram_mem[109408] = 16'b0000000000000000;
	sram_mem[109409] = 16'b0000000000000000;
	sram_mem[109410] = 16'b0000000000000000;
	sram_mem[109411] = 16'b0000000000000000;
	sram_mem[109412] = 16'b0000000000000000;
	sram_mem[109413] = 16'b0000000000000000;
	sram_mem[109414] = 16'b0000000000000000;
	sram_mem[109415] = 16'b0000000000000000;
	sram_mem[109416] = 16'b0000000000000000;
	sram_mem[109417] = 16'b0000000000000000;
	sram_mem[109418] = 16'b0000000000000000;
	sram_mem[109419] = 16'b0000000000000000;
	sram_mem[109420] = 16'b0000000000000000;
	sram_mem[109421] = 16'b0000000000000000;
	sram_mem[109422] = 16'b0000000000000000;
	sram_mem[109423] = 16'b0000000000000000;
	sram_mem[109424] = 16'b0000000000000000;
	sram_mem[109425] = 16'b0000000000000000;
	sram_mem[109426] = 16'b0000000000000000;
	sram_mem[109427] = 16'b0000000000000000;
	sram_mem[109428] = 16'b0000000000000000;
	sram_mem[109429] = 16'b0000000000000000;
	sram_mem[109430] = 16'b0000000000000000;
	sram_mem[109431] = 16'b0000000000000000;
	sram_mem[109432] = 16'b0000000000000000;
	sram_mem[109433] = 16'b0000000000000000;
	sram_mem[109434] = 16'b0000000000000000;
	sram_mem[109435] = 16'b0000000000000000;
	sram_mem[109436] = 16'b0000000000000000;
	sram_mem[109437] = 16'b0000000000000000;
	sram_mem[109438] = 16'b0000000000000000;
	sram_mem[109439] = 16'b0000000000000000;
	sram_mem[109440] = 16'b0000000000000000;
	sram_mem[109441] = 16'b0000000000000000;
	sram_mem[109442] = 16'b0000000000000000;
	sram_mem[109443] = 16'b0000000000000000;
	sram_mem[109444] = 16'b0000000000000000;
	sram_mem[109445] = 16'b0000000000000000;
	sram_mem[109446] = 16'b0000000000000000;
	sram_mem[109447] = 16'b0000000000000000;
	sram_mem[109448] = 16'b0000000000000000;
	sram_mem[109449] = 16'b0000000000000000;
	sram_mem[109450] = 16'b0000000000000000;
	sram_mem[109451] = 16'b0000000000000000;
	sram_mem[109452] = 16'b0000000000000000;
	sram_mem[109453] = 16'b0000000000000000;
	sram_mem[109454] = 16'b0000000000000000;
	sram_mem[109455] = 16'b0000000000000000;
	sram_mem[109456] = 16'b0000000000000000;
	sram_mem[109457] = 16'b0000000000000000;
	sram_mem[109458] = 16'b0000000000000000;
	sram_mem[109459] = 16'b0000000000000000;
	sram_mem[109460] = 16'b0000000000000000;
	sram_mem[109461] = 16'b0000000000000000;
	sram_mem[109462] = 16'b0000000000000000;
	sram_mem[109463] = 16'b0000000000000000;
	sram_mem[109464] = 16'b0000000000000000;
	sram_mem[109465] = 16'b0000000000000000;
	sram_mem[109466] = 16'b0000000000000000;
	sram_mem[109467] = 16'b0000000000000000;
	sram_mem[109468] = 16'b0000000000000000;
	sram_mem[109469] = 16'b0000000000000000;
	sram_mem[109470] = 16'b0000000000000000;
	sram_mem[109471] = 16'b0000000000000000;
	sram_mem[109472] = 16'b0000000000000000;
	sram_mem[109473] = 16'b0000000000000000;
	sram_mem[109474] = 16'b0000000000000000;
	sram_mem[109475] = 16'b0000000000000000;
	sram_mem[109476] = 16'b0000000000000000;
	sram_mem[109477] = 16'b0000000000000000;
	sram_mem[109478] = 16'b0000000000000000;
	sram_mem[109479] = 16'b0000000000000000;
	sram_mem[109480] = 16'b0000000000000000;
	sram_mem[109481] = 16'b0000000000000000;
	sram_mem[109482] = 16'b0000000000000000;
	sram_mem[109483] = 16'b0000000000000000;
	sram_mem[109484] = 16'b0000000000000000;
	sram_mem[109485] = 16'b0000000000000000;
	sram_mem[109486] = 16'b0000000000000000;
	sram_mem[109487] = 16'b0000000000000000;
	sram_mem[109488] = 16'b0000000000000000;
	sram_mem[109489] = 16'b0000000000000000;
	sram_mem[109490] = 16'b0000000000000000;
	sram_mem[109491] = 16'b0000000000000000;
	sram_mem[109492] = 16'b0000000000000000;
	sram_mem[109493] = 16'b0000000000000000;
	sram_mem[109494] = 16'b0000000000000000;
	sram_mem[109495] = 16'b0000000000000000;
	sram_mem[109496] = 16'b0000000000000000;
	sram_mem[109497] = 16'b0000000000000000;
	sram_mem[109498] = 16'b0000000000000000;
	sram_mem[109499] = 16'b0000000000000000;
	sram_mem[109500] = 16'b0000000000000000;
	sram_mem[109501] = 16'b0000000000000000;
	sram_mem[109502] = 16'b0000000000000000;
	sram_mem[109503] = 16'b0000000000000000;
	sram_mem[109504] = 16'b0000000000000000;
	sram_mem[109505] = 16'b0000000000000000;
	sram_mem[109506] = 16'b0000000000000000;
	sram_mem[109507] = 16'b0000000000000000;
	sram_mem[109508] = 16'b0000000000000000;
	sram_mem[109509] = 16'b0000000000000000;
	sram_mem[109510] = 16'b0000000000000000;
	sram_mem[109511] = 16'b0000000000000000;
	sram_mem[109512] = 16'b0000000000000000;
	sram_mem[109513] = 16'b0000000000000000;
	sram_mem[109514] = 16'b0000000000000000;
	sram_mem[109515] = 16'b0000000000000000;
	sram_mem[109516] = 16'b0000000000000000;
	sram_mem[109517] = 16'b0000000000000000;
	sram_mem[109518] = 16'b0000000000000000;
	sram_mem[109519] = 16'b0000000000000000;
	sram_mem[109520] = 16'b0000000000000000;
	sram_mem[109521] = 16'b0000000000000000;
	sram_mem[109522] = 16'b0000000000000000;
	sram_mem[109523] = 16'b0000000000000000;
	sram_mem[109524] = 16'b0000000000000000;
	sram_mem[109525] = 16'b0000000000000000;
	sram_mem[109526] = 16'b0000000000000000;
	sram_mem[109527] = 16'b0000000000000000;
	sram_mem[109528] = 16'b0000000000000000;
	sram_mem[109529] = 16'b0000000000000000;
	sram_mem[109530] = 16'b0000000000000000;
	sram_mem[109531] = 16'b0000000000000000;
	sram_mem[109532] = 16'b0000000000000000;
	sram_mem[109533] = 16'b0000000000000000;
	sram_mem[109534] = 16'b0000000000000000;
	sram_mem[109535] = 16'b0000000000000000;
	sram_mem[109536] = 16'b0000000000000000;
	sram_mem[109537] = 16'b0000000000000000;
	sram_mem[109538] = 16'b0000000000000000;
	sram_mem[109539] = 16'b0000000000000000;
	sram_mem[109540] = 16'b0000000000000000;
	sram_mem[109541] = 16'b0000000000000000;
	sram_mem[109542] = 16'b0000000000000000;
	sram_mem[109543] = 16'b0000000000000000;
	sram_mem[109544] = 16'b0000000000000000;
	sram_mem[109545] = 16'b0000000000000000;
	sram_mem[109546] = 16'b0000000000000000;
	sram_mem[109547] = 16'b0000000000000000;
	sram_mem[109548] = 16'b0000000000000000;
	sram_mem[109549] = 16'b0000000000000000;
	sram_mem[109550] = 16'b0000000000000000;
	sram_mem[109551] = 16'b0000000000000000;
	sram_mem[109552] = 16'b0000000000000000;
	sram_mem[109553] = 16'b0000000000000000;
	sram_mem[109554] = 16'b0000000000000000;
	sram_mem[109555] = 16'b0000000000000000;
	sram_mem[109556] = 16'b0000000000000000;
	sram_mem[109557] = 16'b0000000000000000;
	sram_mem[109558] = 16'b0000000000000000;
	sram_mem[109559] = 16'b0000000000000000;
	sram_mem[109560] = 16'b0000000000000000;
	sram_mem[109561] = 16'b0000000000000000;
	sram_mem[109562] = 16'b0000000000000000;
	sram_mem[109563] = 16'b0000000000000000;
	sram_mem[109564] = 16'b0000000000000000;
	sram_mem[109565] = 16'b0000000000000000;
	sram_mem[109566] = 16'b0000000000000000;
	sram_mem[109567] = 16'b0000000000000000;
	sram_mem[109568] = 16'b0000000000000000;
	sram_mem[109569] = 16'b0000000000000000;
	sram_mem[109570] = 16'b0000000000000000;
	sram_mem[109571] = 16'b0000000000000000;
	sram_mem[109572] = 16'b0000000000000000;
	sram_mem[109573] = 16'b0000000000000000;
	sram_mem[109574] = 16'b0000000000000000;
	sram_mem[109575] = 16'b0000000000000000;
	sram_mem[109576] = 16'b0000000000000000;
	sram_mem[109577] = 16'b0000000000000000;
	sram_mem[109578] = 16'b0000000000000000;
	sram_mem[109579] = 16'b0000000000000000;
	sram_mem[109580] = 16'b0000000000000000;
	sram_mem[109581] = 16'b0000000000000000;
	sram_mem[109582] = 16'b0000000000000000;
	sram_mem[109583] = 16'b0000000000000000;
	sram_mem[109584] = 16'b0000000000000000;
	sram_mem[109585] = 16'b0000000000000000;
	sram_mem[109586] = 16'b0000000000000000;
	sram_mem[109587] = 16'b0000000000000000;
	sram_mem[109588] = 16'b0000000000000000;
	sram_mem[109589] = 16'b0000000000000000;
	sram_mem[109590] = 16'b0000000000000000;
	sram_mem[109591] = 16'b0000000000000000;
	sram_mem[109592] = 16'b0000000000000000;
	sram_mem[109593] = 16'b0000000000000000;
	sram_mem[109594] = 16'b0000000000000000;
	sram_mem[109595] = 16'b0000000000000000;
	sram_mem[109596] = 16'b0000000000000000;
	sram_mem[109597] = 16'b0000000000000000;
	sram_mem[109598] = 16'b0000000000000000;
	sram_mem[109599] = 16'b0000000000000000;
	sram_mem[109600] = 16'b0000000000000000;
	sram_mem[109601] = 16'b0000000000000000;
	sram_mem[109602] = 16'b0000000000000000;
	sram_mem[109603] = 16'b0000000000000000;
	sram_mem[109604] = 16'b0000000000000000;
	sram_mem[109605] = 16'b0000000000000000;
	sram_mem[109606] = 16'b0000000000000000;
	sram_mem[109607] = 16'b0000000000000000;
	sram_mem[109608] = 16'b0000000000000000;
	sram_mem[109609] = 16'b0000000000000000;
	sram_mem[109610] = 16'b0000000000000000;
	sram_mem[109611] = 16'b0000000000000000;
	sram_mem[109612] = 16'b0000000000000000;
	sram_mem[109613] = 16'b0000000000000000;
	sram_mem[109614] = 16'b0000000000000000;
	sram_mem[109615] = 16'b0000000000000000;
	sram_mem[109616] = 16'b0000000000000000;
	sram_mem[109617] = 16'b0000000000000000;
	sram_mem[109618] = 16'b0000000000000000;
	sram_mem[109619] = 16'b0000000000000000;
	sram_mem[109620] = 16'b0000000000000000;
	sram_mem[109621] = 16'b0000000000000000;
	sram_mem[109622] = 16'b0000000000000000;
	sram_mem[109623] = 16'b0000000000000000;
	sram_mem[109624] = 16'b0000000000000000;
	sram_mem[109625] = 16'b0000000000000000;
	sram_mem[109626] = 16'b0000000000000000;
	sram_mem[109627] = 16'b0000000000000000;
	sram_mem[109628] = 16'b0000000000000000;
	sram_mem[109629] = 16'b0000000000000000;
	sram_mem[109630] = 16'b0000000000000000;
	sram_mem[109631] = 16'b0000000000000000;
	sram_mem[109632] = 16'b0000000000000000;
	sram_mem[109633] = 16'b0000000000000000;
	sram_mem[109634] = 16'b0000000000000000;
	sram_mem[109635] = 16'b0000000000000000;
	sram_mem[109636] = 16'b0000000000000000;
	sram_mem[109637] = 16'b0000000000000000;
	sram_mem[109638] = 16'b0000000000000000;
	sram_mem[109639] = 16'b0000000000000000;
	sram_mem[109640] = 16'b0000000000000000;
	sram_mem[109641] = 16'b0000000000000000;
	sram_mem[109642] = 16'b0000000000000000;
	sram_mem[109643] = 16'b0000000000000000;
	sram_mem[109644] = 16'b0000000000000000;
	sram_mem[109645] = 16'b0000000000000000;
	sram_mem[109646] = 16'b0000000000000000;
	sram_mem[109647] = 16'b0000000000000000;
	sram_mem[109648] = 16'b0000000000000000;
	sram_mem[109649] = 16'b0000000000000000;
	sram_mem[109650] = 16'b0000000000000000;
	sram_mem[109651] = 16'b0000000000000000;
	sram_mem[109652] = 16'b0000000000000000;
	sram_mem[109653] = 16'b0000000000000000;
	sram_mem[109654] = 16'b0000000000000000;
	sram_mem[109655] = 16'b0000000000000000;
	sram_mem[109656] = 16'b0000000000000000;
	sram_mem[109657] = 16'b0000000000000000;
	sram_mem[109658] = 16'b0000000000000000;
	sram_mem[109659] = 16'b0000000000000000;
	sram_mem[109660] = 16'b0000000000000000;
	sram_mem[109661] = 16'b0000000000000000;
	sram_mem[109662] = 16'b0000000000000000;
	sram_mem[109663] = 16'b0000000000000000;
	sram_mem[109664] = 16'b0000000000000000;
	sram_mem[109665] = 16'b0000000000000000;
	sram_mem[109666] = 16'b0000000000000000;
	sram_mem[109667] = 16'b0000000000000000;
	sram_mem[109668] = 16'b0000000000000000;
	sram_mem[109669] = 16'b0000000000000000;
	sram_mem[109670] = 16'b0000000000000000;
	sram_mem[109671] = 16'b0000000000000000;
	sram_mem[109672] = 16'b0000000000000000;
	sram_mem[109673] = 16'b0000000000000000;
	sram_mem[109674] = 16'b0000000000000000;
	sram_mem[109675] = 16'b0000000000000000;
	sram_mem[109676] = 16'b0000000000000000;
	sram_mem[109677] = 16'b0000000000000000;
	sram_mem[109678] = 16'b0000000000000000;
	sram_mem[109679] = 16'b0000000000000000;
	sram_mem[109680] = 16'b0000000000000000;
	sram_mem[109681] = 16'b0000000000000000;
	sram_mem[109682] = 16'b0000000000000000;
	sram_mem[109683] = 16'b0000000000000000;
	sram_mem[109684] = 16'b0000000000000000;
	sram_mem[109685] = 16'b0000000000000000;
	sram_mem[109686] = 16'b0000000000000000;
	sram_mem[109687] = 16'b0000000000000000;
	sram_mem[109688] = 16'b0000000000000000;
	sram_mem[109689] = 16'b0000000000000000;
	sram_mem[109690] = 16'b0000000000000000;
	sram_mem[109691] = 16'b0000000000000000;
	sram_mem[109692] = 16'b0000000000000000;
	sram_mem[109693] = 16'b0000000000000000;
	sram_mem[109694] = 16'b0000000000000000;
	sram_mem[109695] = 16'b0000000000000000;
	sram_mem[109696] = 16'b0000000000000000;
	sram_mem[109697] = 16'b0000000000000000;
	sram_mem[109698] = 16'b0000000000000000;
	sram_mem[109699] = 16'b0000000000000000;
	sram_mem[109700] = 16'b0000000000000000;
	sram_mem[109701] = 16'b0000000000000000;
	sram_mem[109702] = 16'b0000000000000000;
	sram_mem[109703] = 16'b0000000000000000;
	sram_mem[109704] = 16'b0000000000000000;
	sram_mem[109705] = 16'b0000000000000000;
	sram_mem[109706] = 16'b0000000000000000;
	sram_mem[109707] = 16'b0000000000000000;
	sram_mem[109708] = 16'b0000000000000000;
	sram_mem[109709] = 16'b0000000000000000;
	sram_mem[109710] = 16'b0000000000000000;
	sram_mem[109711] = 16'b0000000000000000;
	sram_mem[109712] = 16'b0000000000000000;
	sram_mem[109713] = 16'b0000000000000000;
	sram_mem[109714] = 16'b0000000000000000;
	sram_mem[109715] = 16'b0000000000000000;
	sram_mem[109716] = 16'b0000000000000000;
	sram_mem[109717] = 16'b0000000000000000;
	sram_mem[109718] = 16'b0000000000000000;
	sram_mem[109719] = 16'b0000000000000000;
	sram_mem[109720] = 16'b0000000000000000;
	sram_mem[109721] = 16'b0000000000000000;
	sram_mem[109722] = 16'b0000000000000000;
	sram_mem[109723] = 16'b0000000000000000;
	sram_mem[109724] = 16'b0000000000000000;
	sram_mem[109725] = 16'b0000000000000000;
	sram_mem[109726] = 16'b0000000000000000;
	sram_mem[109727] = 16'b0000000000000000;
	sram_mem[109728] = 16'b0000000000000000;
	sram_mem[109729] = 16'b0000000000000000;
	sram_mem[109730] = 16'b0000000000000000;
	sram_mem[109731] = 16'b0000000000000000;
	sram_mem[109732] = 16'b0000000000000000;
	sram_mem[109733] = 16'b0000000000000000;
	sram_mem[109734] = 16'b0000000000000000;
	sram_mem[109735] = 16'b0000000000000000;
	sram_mem[109736] = 16'b0000000000000000;
	sram_mem[109737] = 16'b0000000000000000;
	sram_mem[109738] = 16'b0000000000000000;
	sram_mem[109739] = 16'b0000000000000000;
	sram_mem[109740] = 16'b0000000000000000;
	sram_mem[109741] = 16'b0000000000000000;
	sram_mem[109742] = 16'b0000000000000000;
	sram_mem[109743] = 16'b0000000000000000;
	sram_mem[109744] = 16'b0000000000000000;
	sram_mem[109745] = 16'b0000000000000000;
	sram_mem[109746] = 16'b0000000000000000;
	sram_mem[109747] = 16'b0000000000000000;
	sram_mem[109748] = 16'b0000000000000000;
	sram_mem[109749] = 16'b0000000000000000;
	sram_mem[109750] = 16'b0000000000000000;
	sram_mem[109751] = 16'b0000000000000000;
	sram_mem[109752] = 16'b0000000000000000;
	sram_mem[109753] = 16'b0000000000000000;
	sram_mem[109754] = 16'b0000000000000000;
	sram_mem[109755] = 16'b0000000000000000;
	sram_mem[109756] = 16'b0000000000000000;
	sram_mem[109757] = 16'b0000000000000000;
	sram_mem[109758] = 16'b0000000000000000;
	sram_mem[109759] = 16'b0000000000000000;
	sram_mem[109760] = 16'b0000000000000000;
	sram_mem[109761] = 16'b0000000000000000;
	sram_mem[109762] = 16'b0000000000000000;
	sram_mem[109763] = 16'b0000000000000000;
	sram_mem[109764] = 16'b0000000000000000;
	sram_mem[109765] = 16'b0000000000000000;
	sram_mem[109766] = 16'b0000000000000000;
	sram_mem[109767] = 16'b0000000000000000;
	sram_mem[109768] = 16'b0000000000000000;
	sram_mem[109769] = 16'b0000000000000000;
	sram_mem[109770] = 16'b0000000000000000;
	sram_mem[109771] = 16'b0000000000000000;
	sram_mem[109772] = 16'b0000000000000000;
	sram_mem[109773] = 16'b0000000000000000;
	sram_mem[109774] = 16'b0000000000000000;
	sram_mem[109775] = 16'b0000000000000000;
	sram_mem[109776] = 16'b0000000000000000;
	sram_mem[109777] = 16'b0000000000000000;
	sram_mem[109778] = 16'b0000000000000000;
	sram_mem[109779] = 16'b0000000000000000;
	sram_mem[109780] = 16'b0000000000000000;
	sram_mem[109781] = 16'b0000000000000000;
	sram_mem[109782] = 16'b0000000000000000;
	sram_mem[109783] = 16'b0000000000000000;
	sram_mem[109784] = 16'b0000000000000000;
	sram_mem[109785] = 16'b0000000000000000;
	sram_mem[109786] = 16'b0000000000000000;
	sram_mem[109787] = 16'b0000000000000000;
	sram_mem[109788] = 16'b0000000000000000;
	sram_mem[109789] = 16'b0000000000000000;
	sram_mem[109790] = 16'b0000000000000000;
	sram_mem[109791] = 16'b0000000000000000;
	sram_mem[109792] = 16'b0000000000000000;
	sram_mem[109793] = 16'b0000000000000000;
	sram_mem[109794] = 16'b0000000000000000;
	sram_mem[109795] = 16'b0000000000000000;
	sram_mem[109796] = 16'b0000000000000000;
	sram_mem[109797] = 16'b0000000000000000;
	sram_mem[109798] = 16'b0000000000000000;
	sram_mem[109799] = 16'b0000000000000000;
	sram_mem[109800] = 16'b0000000000000000;
	sram_mem[109801] = 16'b0000000000000000;
	sram_mem[109802] = 16'b0000000000000000;
	sram_mem[109803] = 16'b0000000000000000;
	sram_mem[109804] = 16'b0000000000000000;
	sram_mem[109805] = 16'b0000000000000000;
	sram_mem[109806] = 16'b0000000000000000;
	sram_mem[109807] = 16'b0000000000000000;
	sram_mem[109808] = 16'b0000000000000000;
	sram_mem[109809] = 16'b0000000000000000;
	sram_mem[109810] = 16'b0000000000000000;
	sram_mem[109811] = 16'b0000000000000000;
	sram_mem[109812] = 16'b0000000000000000;
	sram_mem[109813] = 16'b0000000000000000;
	sram_mem[109814] = 16'b0000000000000000;
	sram_mem[109815] = 16'b0000000000000000;
	sram_mem[109816] = 16'b0000000000000000;
	sram_mem[109817] = 16'b0000000000000000;
	sram_mem[109818] = 16'b0000000000000000;
	sram_mem[109819] = 16'b0000000000000000;
	sram_mem[109820] = 16'b0000000000000000;
	sram_mem[109821] = 16'b0000000000000000;
	sram_mem[109822] = 16'b0000000000000000;
	sram_mem[109823] = 16'b0000000000000000;
	sram_mem[109824] = 16'b0000000000000000;
	sram_mem[109825] = 16'b0000000000000000;
	sram_mem[109826] = 16'b0000000000000000;
	sram_mem[109827] = 16'b0000000000000000;
	sram_mem[109828] = 16'b0000000000000000;
	sram_mem[109829] = 16'b0000000000000000;
	sram_mem[109830] = 16'b0000000000000000;
	sram_mem[109831] = 16'b0000000000000000;
	sram_mem[109832] = 16'b0000000000000000;
	sram_mem[109833] = 16'b0000000000000000;
	sram_mem[109834] = 16'b0000000000000000;
	sram_mem[109835] = 16'b0000000000000000;
	sram_mem[109836] = 16'b0000000000000000;
	sram_mem[109837] = 16'b0000000000000000;
	sram_mem[109838] = 16'b0000000000000000;
	sram_mem[109839] = 16'b0000000000000000;
	sram_mem[109840] = 16'b0000000000000000;
	sram_mem[109841] = 16'b0000000000000000;
	sram_mem[109842] = 16'b0000000000000000;
	sram_mem[109843] = 16'b0000000000000000;
	sram_mem[109844] = 16'b0000000000000000;
	sram_mem[109845] = 16'b0000000000000000;
	sram_mem[109846] = 16'b0000000000000000;
	sram_mem[109847] = 16'b0000000000000000;
	sram_mem[109848] = 16'b0000000000000000;
	sram_mem[109849] = 16'b0000000000000000;
	sram_mem[109850] = 16'b0000000000000000;
	sram_mem[109851] = 16'b0000000000000000;
	sram_mem[109852] = 16'b0000000000000000;
	sram_mem[109853] = 16'b0000000000000000;
	sram_mem[109854] = 16'b0000000000000000;
	sram_mem[109855] = 16'b0000000000000000;
	sram_mem[109856] = 16'b0000000000000000;
	sram_mem[109857] = 16'b0000000000000000;
	sram_mem[109858] = 16'b0000000000000000;
	sram_mem[109859] = 16'b0000000000000000;
	sram_mem[109860] = 16'b0000000000000000;
	sram_mem[109861] = 16'b0000000000000000;
	sram_mem[109862] = 16'b0000000000000000;
	sram_mem[109863] = 16'b0000000000000000;
	sram_mem[109864] = 16'b0000000000000000;
	sram_mem[109865] = 16'b0000000000000000;
	sram_mem[109866] = 16'b0000000000000000;
	sram_mem[109867] = 16'b0000000000000000;
	sram_mem[109868] = 16'b0000000000000000;
	sram_mem[109869] = 16'b0000000000000000;
	sram_mem[109870] = 16'b0000000000000000;
	sram_mem[109871] = 16'b0000000000000000;
	sram_mem[109872] = 16'b0000000000000000;
	sram_mem[109873] = 16'b0000000000000000;
	sram_mem[109874] = 16'b0000000000000000;
	sram_mem[109875] = 16'b0000000000000000;
	sram_mem[109876] = 16'b0000000000000000;
	sram_mem[109877] = 16'b0000000000000000;
	sram_mem[109878] = 16'b0000000000000000;
	sram_mem[109879] = 16'b0000000000000000;
	sram_mem[109880] = 16'b0000000000000000;
	sram_mem[109881] = 16'b0000000000000000;
	sram_mem[109882] = 16'b0000000000000000;
	sram_mem[109883] = 16'b0000000000000000;
	sram_mem[109884] = 16'b0000000000000000;
	sram_mem[109885] = 16'b0000000000000000;
	sram_mem[109886] = 16'b0000000000000000;
	sram_mem[109887] = 16'b0000000000000000;
	sram_mem[109888] = 16'b0000000000000000;
	sram_mem[109889] = 16'b0000000000000000;
	sram_mem[109890] = 16'b0000000000000000;
	sram_mem[109891] = 16'b0000000000000000;
	sram_mem[109892] = 16'b0000000000000000;
	sram_mem[109893] = 16'b0000000000000000;
	sram_mem[109894] = 16'b0000000000000000;
	sram_mem[109895] = 16'b0000000000000000;
	sram_mem[109896] = 16'b0000000000000000;
	sram_mem[109897] = 16'b0000000000000000;
	sram_mem[109898] = 16'b0000000000000000;
	sram_mem[109899] = 16'b0000000000000000;
	sram_mem[109900] = 16'b0000000000000000;
	sram_mem[109901] = 16'b0000000000000000;
	sram_mem[109902] = 16'b0000000000000000;
	sram_mem[109903] = 16'b0000000000000000;
	sram_mem[109904] = 16'b0000000000000000;
	sram_mem[109905] = 16'b0000000000000000;
	sram_mem[109906] = 16'b0000000000000000;
	sram_mem[109907] = 16'b0000000000000000;
	sram_mem[109908] = 16'b0000000000000000;
	sram_mem[109909] = 16'b0000000000000000;
	sram_mem[109910] = 16'b0000000000000000;
	sram_mem[109911] = 16'b0000000000000000;
	sram_mem[109912] = 16'b0000000000000000;
	sram_mem[109913] = 16'b0000000000000000;
	sram_mem[109914] = 16'b0000000000000000;
	sram_mem[109915] = 16'b0000000000000000;
	sram_mem[109916] = 16'b0000000000000000;
	sram_mem[109917] = 16'b0000000000000000;
	sram_mem[109918] = 16'b0000000000000000;
	sram_mem[109919] = 16'b0000000000000000;
	sram_mem[109920] = 16'b0000000000000000;
	sram_mem[109921] = 16'b0000000000000000;
	sram_mem[109922] = 16'b0000000000000000;
	sram_mem[109923] = 16'b0000000000000000;
	sram_mem[109924] = 16'b0000000000000000;
	sram_mem[109925] = 16'b0000000000000000;
	sram_mem[109926] = 16'b0000000000000000;
	sram_mem[109927] = 16'b0000000000000000;
	sram_mem[109928] = 16'b0000000000000000;
	sram_mem[109929] = 16'b0000000000000000;
	sram_mem[109930] = 16'b0000000000000000;
	sram_mem[109931] = 16'b0000000000000000;
	sram_mem[109932] = 16'b0000000000000000;
	sram_mem[109933] = 16'b0000000000000000;
	sram_mem[109934] = 16'b0000000000000000;
	sram_mem[109935] = 16'b0000000000000000;
	sram_mem[109936] = 16'b0000000000000000;
	sram_mem[109937] = 16'b0000000000000000;
	sram_mem[109938] = 16'b0000000000000000;
	sram_mem[109939] = 16'b0000000000000000;
	sram_mem[109940] = 16'b0000000000000000;
	sram_mem[109941] = 16'b0000000000000000;
	sram_mem[109942] = 16'b0000000000000000;
	sram_mem[109943] = 16'b0000000000000000;
	sram_mem[109944] = 16'b0000000000000000;
	sram_mem[109945] = 16'b0000000000000000;
	sram_mem[109946] = 16'b0000000000000000;
	sram_mem[109947] = 16'b0000000000000000;
	sram_mem[109948] = 16'b0000000000000000;
	sram_mem[109949] = 16'b0000000000000000;
	sram_mem[109950] = 16'b0000000000000000;
	sram_mem[109951] = 16'b0000000000000000;
	sram_mem[109952] = 16'b0000000000000000;
	sram_mem[109953] = 16'b0000000000000000;
	sram_mem[109954] = 16'b0000000000000000;
	sram_mem[109955] = 16'b0000000000000000;
	sram_mem[109956] = 16'b0000000000000000;
	sram_mem[109957] = 16'b0000000000000000;
	sram_mem[109958] = 16'b0000000000000000;
	sram_mem[109959] = 16'b0000000000000000;
	sram_mem[109960] = 16'b0000000000000000;
	sram_mem[109961] = 16'b0000000000000000;
	sram_mem[109962] = 16'b0000000000000000;
	sram_mem[109963] = 16'b0000000000000000;
	sram_mem[109964] = 16'b0000000000000000;
	sram_mem[109965] = 16'b0000000000000000;
	sram_mem[109966] = 16'b0000000000000000;
	sram_mem[109967] = 16'b0000000000000000;
	sram_mem[109968] = 16'b0000000000000000;
	sram_mem[109969] = 16'b0000000000000000;
	sram_mem[109970] = 16'b0000000000000000;
	sram_mem[109971] = 16'b0000000000000000;
	sram_mem[109972] = 16'b0000000000000000;
	sram_mem[109973] = 16'b0000000000000000;
	sram_mem[109974] = 16'b0000000000000000;
	sram_mem[109975] = 16'b0000000000000000;
	sram_mem[109976] = 16'b0000000000000000;
	sram_mem[109977] = 16'b0000000000000000;
	sram_mem[109978] = 16'b0000000000000000;
	sram_mem[109979] = 16'b0000000000000000;
	sram_mem[109980] = 16'b0000000000000000;
	sram_mem[109981] = 16'b0000000000000000;
	sram_mem[109982] = 16'b0000000000000000;
	sram_mem[109983] = 16'b0000000000000000;
	sram_mem[109984] = 16'b0000000000000000;
	sram_mem[109985] = 16'b0000000000000000;
	sram_mem[109986] = 16'b0000000000000000;
	sram_mem[109987] = 16'b0000000000000000;
	sram_mem[109988] = 16'b0000000000000000;
	sram_mem[109989] = 16'b0000000000000000;
	sram_mem[109990] = 16'b0000000000000000;
	sram_mem[109991] = 16'b0000000000000000;
	sram_mem[109992] = 16'b0000000000000000;
	sram_mem[109993] = 16'b0000000000000000;
	sram_mem[109994] = 16'b0000000000000000;
	sram_mem[109995] = 16'b0000000000000000;
	sram_mem[109996] = 16'b0000000000000000;
	sram_mem[109997] = 16'b0000000000000000;
	sram_mem[109998] = 16'b0000000000000000;
	sram_mem[109999] = 16'b0000000000000000;
	sram_mem[110000] = 16'b0000000000000000;
	sram_mem[110001] = 16'b0000000000000000;
	sram_mem[110002] = 16'b0000000000000000;
	sram_mem[110003] = 16'b0000000000000000;
	sram_mem[110004] = 16'b0000000000000000;
	sram_mem[110005] = 16'b0000000000000000;
	sram_mem[110006] = 16'b0000000000000000;
	sram_mem[110007] = 16'b0000000000000000;
	sram_mem[110008] = 16'b0000000000000000;
	sram_mem[110009] = 16'b0000000000000000;
	sram_mem[110010] = 16'b0000000000000000;
	sram_mem[110011] = 16'b0000000000000000;
	sram_mem[110012] = 16'b0000000000000000;
	sram_mem[110013] = 16'b0000000000000000;
	sram_mem[110014] = 16'b0000000000000000;
	sram_mem[110015] = 16'b0000000000000000;
	sram_mem[110016] = 16'b0000000000000000;
	sram_mem[110017] = 16'b0000000000000000;
	sram_mem[110018] = 16'b0000000000000000;
	sram_mem[110019] = 16'b0000000000000000;
	sram_mem[110020] = 16'b0000000000000000;
	sram_mem[110021] = 16'b0000000000000000;
	sram_mem[110022] = 16'b0000000000000000;
	sram_mem[110023] = 16'b0000000000000000;
	sram_mem[110024] = 16'b0000000000000000;
	sram_mem[110025] = 16'b0000000000000000;
	sram_mem[110026] = 16'b0000000000000000;
	sram_mem[110027] = 16'b0000000000000000;
	sram_mem[110028] = 16'b0000000000000000;
	sram_mem[110029] = 16'b0000000000000000;
	sram_mem[110030] = 16'b0000000000000000;
	sram_mem[110031] = 16'b0000000000000000;
	sram_mem[110032] = 16'b0000000000000000;
	sram_mem[110033] = 16'b0000000000000000;
	sram_mem[110034] = 16'b0000000000000000;
	sram_mem[110035] = 16'b0000000000000000;
	sram_mem[110036] = 16'b0000000000000000;
	sram_mem[110037] = 16'b0000000000000000;
	sram_mem[110038] = 16'b0000000000000000;
	sram_mem[110039] = 16'b0000000000000000;
	sram_mem[110040] = 16'b0000000000000000;
	sram_mem[110041] = 16'b0000000000000000;
	sram_mem[110042] = 16'b0000000000000000;
	sram_mem[110043] = 16'b0000000000000000;
	sram_mem[110044] = 16'b0000000000000000;
	sram_mem[110045] = 16'b0000000000000000;
	sram_mem[110046] = 16'b0000000000000000;
	sram_mem[110047] = 16'b0000000000000000;
	sram_mem[110048] = 16'b0000000000000000;
	sram_mem[110049] = 16'b0000000000000000;
	sram_mem[110050] = 16'b0000000000000000;
	sram_mem[110051] = 16'b0000000000000000;
	sram_mem[110052] = 16'b0000000000000000;
	sram_mem[110053] = 16'b0000000000000000;
	sram_mem[110054] = 16'b0000000000000000;
	sram_mem[110055] = 16'b0000000000000000;
	sram_mem[110056] = 16'b0000000000000000;
	sram_mem[110057] = 16'b0000000000000000;
	sram_mem[110058] = 16'b0000000000000000;
	sram_mem[110059] = 16'b0000000000000000;
	sram_mem[110060] = 16'b0000000000000000;
	sram_mem[110061] = 16'b0000000000000000;
	sram_mem[110062] = 16'b0000000000000000;
	sram_mem[110063] = 16'b0000000000000000;
	sram_mem[110064] = 16'b0000000000000000;
	sram_mem[110065] = 16'b0000000000000000;
	sram_mem[110066] = 16'b0000000000000000;
	sram_mem[110067] = 16'b0000000000000000;
	sram_mem[110068] = 16'b0000000000000000;
	sram_mem[110069] = 16'b0000000000000000;
	sram_mem[110070] = 16'b0000000000000000;
	sram_mem[110071] = 16'b0000000000000000;
	sram_mem[110072] = 16'b0000000000000000;
	sram_mem[110073] = 16'b0000000000000000;
	sram_mem[110074] = 16'b0000000000000000;
	sram_mem[110075] = 16'b0000000000000000;
	sram_mem[110076] = 16'b0000000000000000;
	sram_mem[110077] = 16'b0000000000000000;
	sram_mem[110078] = 16'b0000000000000000;
	sram_mem[110079] = 16'b0000000000000000;
	sram_mem[110080] = 16'b0000000000000000;
	sram_mem[110081] = 16'b0000000000000000;
	sram_mem[110082] = 16'b0000000000000000;
	sram_mem[110083] = 16'b0000000000000000;
	sram_mem[110084] = 16'b0000000000000000;
	sram_mem[110085] = 16'b0000000000000000;
	sram_mem[110086] = 16'b0000000000000000;
	sram_mem[110087] = 16'b0000000000000000;
	sram_mem[110088] = 16'b0000000000000000;
	sram_mem[110089] = 16'b0000000000000000;
	sram_mem[110090] = 16'b0000000000000000;
	sram_mem[110091] = 16'b0000000000000000;
	sram_mem[110092] = 16'b0000000000000000;
	sram_mem[110093] = 16'b0000000000000000;
	sram_mem[110094] = 16'b0000000000000000;
	sram_mem[110095] = 16'b0000000000000000;
	sram_mem[110096] = 16'b0000000000000000;
	sram_mem[110097] = 16'b0000000000000000;
	sram_mem[110098] = 16'b0000000000000000;
	sram_mem[110099] = 16'b0000000000000000;
	sram_mem[110100] = 16'b0000000000000000;
	sram_mem[110101] = 16'b0000000000000000;
	sram_mem[110102] = 16'b0000000000000000;
	sram_mem[110103] = 16'b0000000000000000;
	sram_mem[110104] = 16'b0000000000000000;
	sram_mem[110105] = 16'b0000000000000000;
	sram_mem[110106] = 16'b0000000000000000;
	sram_mem[110107] = 16'b0000000000000000;
	sram_mem[110108] = 16'b0000000000000000;
	sram_mem[110109] = 16'b0000000000000000;
	sram_mem[110110] = 16'b0000000000000000;
	sram_mem[110111] = 16'b0000000000000000;
	sram_mem[110112] = 16'b0000000000000000;
	sram_mem[110113] = 16'b0000000000000000;
	sram_mem[110114] = 16'b0000000000000000;
	sram_mem[110115] = 16'b0000000000000000;
	sram_mem[110116] = 16'b0000000000000000;
	sram_mem[110117] = 16'b0000000000000000;
	sram_mem[110118] = 16'b0000000000000000;
	sram_mem[110119] = 16'b0000000000000000;
	sram_mem[110120] = 16'b0000000000000000;
	sram_mem[110121] = 16'b0000000000000000;
	sram_mem[110122] = 16'b0000000000000000;
	sram_mem[110123] = 16'b0000000000000000;
	sram_mem[110124] = 16'b0000000000000000;
	sram_mem[110125] = 16'b0000000000000000;
	sram_mem[110126] = 16'b0000000000000000;
	sram_mem[110127] = 16'b0000000000000000;
	sram_mem[110128] = 16'b0000000000000000;
	sram_mem[110129] = 16'b0000000000000000;
	sram_mem[110130] = 16'b0000000000000000;
	sram_mem[110131] = 16'b0000000000000000;
	sram_mem[110132] = 16'b0000000000000000;
	sram_mem[110133] = 16'b0000000000000000;
	sram_mem[110134] = 16'b0000000000000000;
	sram_mem[110135] = 16'b0000000000000000;
	sram_mem[110136] = 16'b0000000000000000;
	sram_mem[110137] = 16'b0000000000000000;
	sram_mem[110138] = 16'b0000000000000000;
	sram_mem[110139] = 16'b0000000000000000;
	sram_mem[110140] = 16'b0000000000000000;
	sram_mem[110141] = 16'b0000000000000000;
	sram_mem[110142] = 16'b0000000000000000;
	sram_mem[110143] = 16'b0000000000000000;
	sram_mem[110144] = 16'b0000000000000000;
	sram_mem[110145] = 16'b0000000000000000;
	sram_mem[110146] = 16'b0000000000000000;
	sram_mem[110147] = 16'b0000000000000000;
	sram_mem[110148] = 16'b0000000000000000;
	sram_mem[110149] = 16'b0000000000000000;
	sram_mem[110150] = 16'b0000000000000000;
	sram_mem[110151] = 16'b0000000000000000;
	sram_mem[110152] = 16'b0000000000000000;
	sram_mem[110153] = 16'b0000000000000000;
	sram_mem[110154] = 16'b0000000000000000;
	sram_mem[110155] = 16'b0000000000000000;
	sram_mem[110156] = 16'b0000000000000000;
	sram_mem[110157] = 16'b0000000000000000;
	sram_mem[110158] = 16'b0000000000000000;
	sram_mem[110159] = 16'b0000000000000000;
	sram_mem[110160] = 16'b0000000000000000;
	sram_mem[110161] = 16'b0000000000000000;
	sram_mem[110162] = 16'b0000000000000000;
	sram_mem[110163] = 16'b0000000000000000;
	sram_mem[110164] = 16'b0000000000000000;
	sram_mem[110165] = 16'b0000000000000000;
	sram_mem[110166] = 16'b0000000000000000;
	sram_mem[110167] = 16'b0000000000000000;
	sram_mem[110168] = 16'b0000000000000000;
	sram_mem[110169] = 16'b0000000000000000;
	sram_mem[110170] = 16'b0000000000000000;
	sram_mem[110171] = 16'b0000000000000000;
	sram_mem[110172] = 16'b0000000000000000;
	sram_mem[110173] = 16'b0000000000000000;
	sram_mem[110174] = 16'b0000000000000000;
	sram_mem[110175] = 16'b0000000000000000;
	sram_mem[110176] = 16'b0000000000000000;
	sram_mem[110177] = 16'b0000000000000000;
	sram_mem[110178] = 16'b0000000000000000;
	sram_mem[110179] = 16'b0000000000000000;
	sram_mem[110180] = 16'b0000000000000000;
	sram_mem[110181] = 16'b0000000000000000;
	sram_mem[110182] = 16'b0000000000000000;
	sram_mem[110183] = 16'b0000000000000000;
	sram_mem[110184] = 16'b0000000000000000;
	sram_mem[110185] = 16'b0000000000000000;
	sram_mem[110186] = 16'b0000000000000000;
	sram_mem[110187] = 16'b0000000000000000;
	sram_mem[110188] = 16'b0000000000000000;
	sram_mem[110189] = 16'b0000000000000000;
	sram_mem[110190] = 16'b0000000000000000;
	sram_mem[110191] = 16'b0000000000000000;
	sram_mem[110192] = 16'b0000000000000000;
	sram_mem[110193] = 16'b0000000000000000;
	sram_mem[110194] = 16'b0000000000000000;
	sram_mem[110195] = 16'b0000000000000000;
	sram_mem[110196] = 16'b0000000000000000;
	sram_mem[110197] = 16'b0000000000000000;
	sram_mem[110198] = 16'b0000000000000000;
	sram_mem[110199] = 16'b0000000000000000;
	sram_mem[110200] = 16'b0000000000000000;
	sram_mem[110201] = 16'b0000000000000000;
	sram_mem[110202] = 16'b0000000000000000;
	sram_mem[110203] = 16'b0000000000000000;
	sram_mem[110204] = 16'b0000000000000000;
	sram_mem[110205] = 16'b0000000000000000;
	sram_mem[110206] = 16'b0000000000000000;
	sram_mem[110207] = 16'b0000000000000000;
	sram_mem[110208] = 16'b0000000000000000;
	sram_mem[110209] = 16'b0000000000000000;
	sram_mem[110210] = 16'b0000000000000000;
	sram_mem[110211] = 16'b0000000000000000;
	sram_mem[110212] = 16'b0000000000000000;
	sram_mem[110213] = 16'b0000000000000000;
	sram_mem[110214] = 16'b0000000000000000;
	sram_mem[110215] = 16'b0000000000000000;
	sram_mem[110216] = 16'b0000000000000000;
	sram_mem[110217] = 16'b0000000000000000;
	sram_mem[110218] = 16'b0000000000000000;
	sram_mem[110219] = 16'b0000000000000000;
	sram_mem[110220] = 16'b0000000000000000;
	sram_mem[110221] = 16'b0000000000000000;
	sram_mem[110222] = 16'b0000000000000000;
	sram_mem[110223] = 16'b0000000000000000;
	sram_mem[110224] = 16'b0000000000000000;
	sram_mem[110225] = 16'b0000000000000000;
	sram_mem[110226] = 16'b0000000000000000;
	sram_mem[110227] = 16'b0000000000000000;
	sram_mem[110228] = 16'b0000000000000000;
	sram_mem[110229] = 16'b0000000000000000;
	sram_mem[110230] = 16'b0000000000000000;
	sram_mem[110231] = 16'b0000000000000000;
	sram_mem[110232] = 16'b0000000000000000;
	sram_mem[110233] = 16'b0000000000000000;
	sram_mem[110234] = 16'b0000000000000000;
	sram_mem[110235] = 16'b0000000000000000;
	sram_mem[110236] = 16'b0000000000000000;
	sram_mem[110237] = 16'b0000000000000000;
	sram_mem[110238] = 16'b0000000000000000;
	sram_mem[110239] = 16'b0000000000000000;
	sram_mem[110240] = 16'b0000000000000000;
	sram_mem[110241] = 16'b0000000000000000;
	sram_mem[110242] = 16'b0000000000000000;
	sram_mem[110243] = 16'b0000000000000000;
	sram_mem[110244] = 16'b0000000000000000;
	sram_mem[110245] = 16'b0000000000000000;
	sram_mem[110246] = 16'b0000000000000000;
	sram_mem[110247] = 16'b0000000000000000;
	sram_mem[110248] = 16'b0000000000000000;
	sram_mem[110249] = 16'b0000000000000000;
	sram_mem[110250] = 16'b0000000000000000;
	sram_mem[110251] = 16'b0000000000000000;
	sram_mem[110252] = 16'b0000000000000000;
	sram_mem[110253] = 16'b0000000000000000;
	sram_mem[110254] = 16'b0000000000000000;
	sram_mem[110255] = 16'b0000000000000000;
	sram_mem[110256] = 16'b0000000000000000;
	sram_mem[110257] = 16'b0000000000000000;
	sram_mem[110258] = 16'b0000000000000000;
	sram_mem[110259] = 16'b0000000000000000;
	sram_mem[110260] = 16'b0000000000000000;
	sram_mem[110261] = 16'b0000000000000000;
	sram_mem[110262] = 16'b0000000000000000;
	sram_mem[110263] = 16'b0000000000000000;
	sram_mem[110264] = 16'b0000000000000000;
	sram_mem[110265] = 16'b0000000000000000;
	sram_mem[110266] = 16'b0000000000000000;
	sram_mem[110267] = 16'b0000000000000000;
	sram_mem[110268] = 16'b0000000000000000;
	sram_mem[110269] = 16'b0000000000000000;
	sram_mem[110270] = 16'b0000000000000000;
	sram_mem[110271] = 16'b0000000000000000;
	sram_mem[110272] = 16'b0000000000000000;
	sram_mem[110273] = 16'b0000000000000000;
	sram_mem[110274] = 16'b0000000000000000;
	sram_mem[110275] = 16'b0000000000000000;
	sram_mem[110276] = 16'b0000000000000000;
	sram_mem[110277] = 16'b0000000000000000;
	sram_mem[110278] = 16'b0000000000000000;
	sram_mem[110279] = 16'b0000000000000000;
	sram_mem[110280] = 16'b0000000000000000;
	sram_mem[110281] = 16'b0000000000000000;
	sram_mem[110282] = 16'b0000000000000000;
	sram_mem[110283] = 16'b0000000000000000;
	sram_mem[110284] = 16'b0000000000000000;
	sram_mem[110285] = 16'b0000000000000000;
	sram_mem[110286] = 16'b0000000000000000;
	sram_mem[110287] = 16'b0000000000000000;
	sram_mem[110288] = 16'b0000000000000000;
	sram_mem[110289] = 16'b0000000000000000;
	sram_mem[110290] = 16'b0000000000000000;
	sram_mem[110291] = 16'b0000000000000000;
	sram_mem[110292] = 16'b0000000000000000;
	sram_mem[110293] = 16'b0000000000000000;
	sram_mem[110294] = 16'b0000000000000000;
	sram_mem[110295] = 16'b0000000000000000;
	sram_mem[110296] = 16'b0000000000000000;
	sram_mem[110297] = 16'b0000000000000000;
	sram_mem[110298] = 16'b0000000000000000;
	sram_mem[110299] = 16'b0000000000000000;
	sram_mem[110300] = 16'b0000000000000000;
	sram_mem[110301] = 16'b0000000000000000;
	sram_mem[110302] = 16'b0000000000000000;
	sram_mem[110303] = 16'b0000000000000000;
	sram_mem[110304] = 16'b0000000000000000;
	sram_mem[110305] = 16'b0000000000000000;
	sram_mem[110306] = 16'b0000000000000000;
	sram_mem[110307] = 16'b0000000000000000;
	sram_mem[110308] = 16'b0000000000000000;
	sram_mem[110309] = 16'b0000000000000000;
	sram_mem[110310] = 16'b0000000000000000;
	sram_mem[110311] = 16'b0000000000000000;
	sram_mem[110312] = 16'b0000000000000000;
	sram_mem[110313] = 16'b0000000000000000;
	sram_mem[110314] = 16'b0000000000000000;
	sram_mem[110315] = 16'b0000000000000000;
	sram_mem[110316] = 16'b0000000000000000;
	sram_mem[110317] = 16'b0000000000000000;
	sram_mem[110318] = 16'b0000000000000000;
	sram_mem[110319] = 16'b0000000000000000;
	sram_mem[110320] = 16'b0000000000000000;
	sram_mem[110321] = 16'b0000000000000000;
	sram_mem[110322] = 16'b0000000000000000;
	sram_mem[110323] = 16'b0000000000000000;
	sram_mem[110324] = 16'b0000000000000000;
	sram_mem[110325] = 16'b0000000000000000;
	sram_mem[110326] = 16'b0000000000000000;
	sram_mem[110327] = 16'b0000000000000000;
	sram_mem[110328] = 16'b0000000000000000;
	sram_mem[110329] = 16'b0000000000000000;
	sram_mem[110330] = 16'b0000000000000000;
	sram_mem[110331] = 16'b0000000000000000;
	sram_mem[110332] = 16'b0000000000000000;
	sram_mem[110333] = 16'b0000000000000000;
	sram_mem[110334] = 16'b0000000000000000;
	sram_mem[110335] = 16'b0000000000000000;
	sram_mem[110336] = 16'b0000000000000000;
	sram_mem[110337] = 16'b0000000000000000;
	sram_mem[110338] = 16'b0000000000000000;
	sram_mem[110339] = 16'b0000000000000000;
	sram_mem[110340] = 16'b0000000000000000;
	sram_mem[110341] = 16'b0000000000000000;
	sram_mem[110342] = 16'b0000000000000000;
	sram_mem[110343] = 16'b0000000000000000;
	sram_mem[110344] = 16'b0000000000000000;
	sram_mem[110345] = 16'b0000000000000000;
	sram_mem[110346] = 16'b0000000000000000;
	sram_mem[110347] = 16'b0000000000000000;
	sram_mem[110348] = 16'b0000000000000000;
	sram_mem[110349] = 16'b0000000000000000;
	sram_mem[110350] = 16'b0000000000000000;
	sram_mem[110351] = 16'b0000000000000000;
	sram_mem[110352] = 16'b0000000000000000;
	sram_mem[110353] = 16'b0000000000000000;
	sram_mem[110354] = 16'b0000000000000000;
	sram_mem[110355] = 16'b0000000000000000;
	sram_mem[110356] = 16'b0000000000000000;
	sram_mem[110357] = 16'b0000000000000000;
	sram_mem[110358] = 16'b0000000000000000;
	sram_mem[110359] = 16'b0000000000000000;
	sram_mem[110360] = 16'b0000000000000000;
	sram_mem[110361] = 16'b0000000000000000;
	sram_mem[110362] = 16'b0000000000000000;
	sram_mem[110363] = 16'b0000000000000000;
	sram_mem[110364] = 16'b0000000000000000;
	sram_mem[110365] = 16'b0000000000000000;
	sram_mem[110366] = 16'b0000000000000000;
	sram_mem[110367] = 16'b0000000000000000;
	sram_mem[110368] = 16'b0000000000000000;
	sram_mem[110369] = 16'b0000000000000000;
	sram_mem[110370] = 16'b0000000000000000;
	sram_mem[110371] = 16'b0000000000000000;
	sram_mem[110372] = 16'b0000000000000000;
	sram_mem[110373] = 16'b0000000000000000;
	sram_mem[110374] = 16'b0000000000000000;
	sram_mem[110375] = 16'b0000000000000000;
	sram_mem[110376] = 16'b0000000000000000;
	sram_mem[110377] = 16'b0000000000000000;
	sram_mem[110378] = 16'b0000000000000000;
	sram_mem[110379] = 16'b0000000000000000;
	sram_mem[110380] = 16'b0000000000000000;
	sram_mem[110381] = 16'b0000000000000000;
	sram_mem[110382] = 16'b0000000000000000;
	sram_mem[110383] = 16'b0000000000000000;
	sram_mem[110384] = 16'b0000000000000000;
	sram_mem[110385] = 16'b0000000000000000;
	sram_mem[110386] = 16'b0000000000000000;
	sram_mem[110387] = 16'b0000000000000000;
	sram_mem[110388] = 16'b0000000000000000;
	sram_mem[110389] = 16'b0000000000000000;
	sram_mem[110390] = 16'b0000000000000000;
	sram_mem[110391] = 16'b0000000000000000;
	sram_mem[110392] = 16'b0000000000000000;
	sram_mem[110393] = 16'b0000000000000000;
	sram_mem[110394] = 16'b0000000000000000;
	sram_mem[110395] = 16'b0000000000000000;
	sram_mem[110396] = 16'b0000000000000000;
	sram_mem[110397] = 16'b0000000000000000;
	sram_mem[110398] = 16'b0000000000000000;
	sram_mem[110399] = 16'b0000000000000000;
	sram_mem[110400] = 16'b0000000000000000;
	sram_mem[110401] = 16'b0000000000000000;
	sram_mem[110402] = 16'b0000000000000000;
	sram_mem[110403] = 16'b0000000000000000;
	sram_mem[110404] = 16'b0000000000000000;
	sram_mem[110405] = 16'b0000000000000000;
	sram_mem[110406] = 16'b0000000000000000;
	sram_mem[110407] = 16'b0000000000000000;
	sram_mem[110408] = 16'b0000000000000000;
	sram_mem[110409] = 16'b0000000000000000;
	sram_mem[110410] = 16'b0000000000000000;
	sram_mem[110411] = 16'b0000000000000000;
	sram_mem[110412] = 16'b0000000000000000;
	sram_mem[110413] = 16'b0000000000000000;
	sram_mem[110414] = 16'b0000000000000000;
	sram_mem[110415] = 16'b0000000000000000;
	sram_mem[110416] = 16'b0000000000000000;
	sram_mem[110417] = 16'b0000000000000000;
	sram_mem[110418] = 16'b0000000000000000;
	sram_mem[110419] = 16'b0000000000000000;
	sram_mem[110420] = 16'b0000000000000000;
	sram_mem[110421] = 16'b0000000000000000;
	sram_mem[110422] = 16'b0000000000000000;
	sram_mem[110423] = 16'b0000000000000000;
	sram_mem[110424] = 16'b0000000000000000;
	sram_mem[110425] = 16'b0000000000000000;
	sram_mem[110426] = 16'b0000000000000000;
	sram_mem[110427] = 16'b0000000000000000;
	sram_mem[110428] = 16'b0000000000000000;
	sram_mem[110429] = 16'b0000000000000000;
	sram_mem[110430] = 16'b0000000000000000;
	sram_mem[110431] = 16'b0000000000000000;
	sram_mem[110432] = 16'b0000000000000000;
	sram_mem[110433] = 16'b0000000000000000;
	sram_mem[110434] = 16'b0000000000000000;
	sram_mem[110435] = 16'b0000000000000000;
	sram_mem[110436] = 16'b0000000000000000;
	sram_mem[110437] = 16'b0000000000000000;
	sram_mem[110438] = 16'b0000000000000000;
	sram_mem[110439] = 16'b0000000000000000;
	sram_mem[110440] = 16'b0000000000000000;
	sram_mem[110441] = 16'b0000000000000000;
	sram_mem[110442] = 16'b0000000000000000;
	sram_mem[110443] = 16'b0000000000000000;
	sram_mem[110444] = 16'b0000000000000000;
	sram_mem[110445] = 16'b0000000000000000;
	sram_mem[110446] = 16'b0000000000000000;
	sram_mem[110447] = 16'b0000000000000000;
	sram_mem[110448] = 16'b0000000000000000;
	sram_mem[110449] = 16'b0000000000000000;
	sram_mem[110450] = 16'b0000000000000000;
	sram_mem[110451] = 16'b0000000000000000;
	sram_mem[110452] = 16'b0000000000000000;
	sram_mem[110453] = 16'b0000000000000000;
	sram_mem[110454] = 16'b0000000000000000;
	sram_mem[110455] = 16'b0000000000000000;
	sram_mem[110456] = 16'b0000000000000000;
	sram_mem[110457] = 16'b0000000000000000;
	sram_mem[110458] = 16'b0000000000000000;
	sram_mem[110459] = 16'b0000000000000000;
	sram_mem[110460] = 16'b0000000000000000;
	sram_mem[110461] = 16'b0000000000000000;
	sram_mem[110462] = 16'b0000000000000000;
	sram_mem[110463] = 16'b0000000000000000;
	sram_mem[110464] = 16'b0000000000000000;
	sram_mem[110465] = 16'b0000000000000000;
	sram_mem[110466] = 16'b0000000000000000;
	sram_mem[110467] = 16'b0000000000000000;
	sram_mem[110468] = 16'b0000000000000000;
	sram_mem[110469] = 16'b0000000000000000;
	sram_mem[110470] = 16'b0000000000000000;
	sram_mem[110471] = 16'b0000000000000000;
	sram_mem[110472] = 16'b0000000000000000;
	sram_mem[110473] = 16'b0000000000000000;
	sram_mem[110474] = 16'b0000000000000000;
	sram_mem[110475] = 16'b0000000000000000;
	sram_mem[110476] = 16'b0000000000000000;
	sram_mem[110477] = 16'b0000000000000000;
	sram_mem[110478] = 16'b0000000000000000;
	sram_mem[110479] = 16'b0000000000000000;
	sram_mem[110480] = 16'b0000000000000000;
	sram_mem[110481] = 16'b0000000000000000;
	sram_mem[110482] = 16'b0000000000000000;
	sram_mem[110483] = 16'b0000000000000000;
	sram_mem[110484] = 16'b0000000000000000;
	sram_mem[110485] = 16'b0000000000000000;
	sram_mem[110486] = 16'b0000000000000000;
	sram_mem[110487] = 16'b0000000000000000;
	sram_mem[110488] = 16'b0000000000000000;
	sram_mem[110489] = 16'b0000000000000000;
	sram_mem[110490] = 16'b0000000000000000;
	sram_mem[110491] = 16'b0000000000000000;
	sram_mem[110492] = 16'b0000000000000000;
	sram_mem[110493] = 16'b0000000000000000;
	sram_mem[110494] = 16'b0000000000000000;
	sram_mem[110495] = 16'b0000000000000000;
	sram_mem[110496] = 16'b0000000000000000;
	sram_mem[110497] = 16'b0000000000000000;
	sram_mem[110498] = 16'b0000000000000000;
	sram_mem[110499] = 16'b0000000000000000;
	sram_mem[110500] = 16'b0000000000000000;
	sram_mem[110501] = 16'b0000000000000000;
	sram_mem[110502] = 16'b0000000000000000;
	sram_mem[110503] = 16'b0000000000000000;
	sram_mem[110504] = 16'b0000000000000000;
	sram_mem[110505] = 16'b0000000000000000;
	sram_mem[110506] = 16'b0000000000000000;
	sram_mem[110507] = 16'b0000000000000000;
	sram_mem[110508] = 16'b0000000000000000;
	sram_mem[110509] = 16'b0000000000000000;
	sram_mem[110510] = 16'b0000000000000000;
	sram_mem[110511] = 16'b0000000000000000;
	sram_mem[110512] = 16'b0000000000000000;
	sram_mem[110513] = 16'b0000000000000000;
	sram_mem[110514] = 16'b0000000000000000;
	sram_mem[110515] = 16'b0000000000000000;
	sram_mem[110516] = 16'b0000000000000000;
	sram_mem[110517] = 16'b0000000000000000;
	sram_mem[110518] = 16'b0000000000000000;
	sram_mem[110519] = 16'b0000000000000000;
	sram_mem[110520] = 16'b0000000000000000;
	sram_mem[110521] = 16'b0000000000000000;
	sram_mem[110522] = 16'b0000000000000000;
	sram_mem[110523] = 16'b0000000000000000;
	sram_mem[110524] = 16'b0000000000000000;
	sram_mem[110525] = 16'b0000000000000000;
	sram_mem[110526] = 16'b0000000000000000;
	sram_mem[110527] = 16'b0000000000000000;
	sram_mem[110528] = 16'b0000000000000000;
	sram_mem[110529] = 16'b0000000000000000;
	sram_mem[110530] = 16'b0000000000000000;
	sram_mem[110531] = 16'b0000000000000000;
	sram_mem[110532] = 16'b0000000000000000;
	sram_mem[110533] = 16'b0000000000000000;
	sram_mem[110534] = 16'b0000000000000000;
	sram_mem[110535] = 16'b0000000000000000;
	sram_mem[110536] = 16'b0000000000000000;
	sram_mem[110537] = 16'b0000000000000000;
	sram_mem[110538] = 16'b0000000000000000;
	sram_mem[110539] = 16'b0000000000000000;
	sram_mem[110540] = 16'b0000000000000000;
	sram_mem[110541] = 16'b0000000000000000;
	sram_mem[110542] = 16'b0000000000000000;
	sram_mem[110543] = 16'b0000000000000000;
	sram_mem[110544] = 16'b0000000000000000;
	sram_mem[110545] = 16'b0000000000000000;
	sram_mem[110546] = 16'b0000000000000000;
	sram_mem[110547] = 16'b0000000000000000;
	sram_mem[110548] = 16'b0000000000000000;
	sram_mem[110549] = 16'b0000000000000000;
	sram_mem[110550] = 16'b0000000000000000;
	sram_mem[110551] = 16'b0000000000000000;
	sram_mem[110552] = 16'b0000000000000000;
	sram_mem[110553] = 16'b0000000000000000;
	sram_mem[110554] = 16'b0000000000000000;
	sram_mem[110555] = 16'b0000000000000000;
	sram_mem[110556] = 16'b0000000000000000;
	sram_mem[110557] = 16'b0000000000000000;
	sram_mem[110558] = 16'b0000000000000000;
	sram_mem[110559] = 16'b0000000000000000;
	sram_mem[110560] = 16'b0000000000000000;
	sram_mem[110561] = 16'b0000000000000000;
	sram_mem[110562] = 16'b0000000000000000;
	sram_mem[110563] = 16'b0000000000000000;
	sram_mem[110564] = 16'b0000000000000000;
	sram_mem[110565] = 16'b0000000000000000;
	sram_mem[110566] = 16'b0000000000000000;
	sram_mem[110567] = 16'b0000000000000000;
	sram_mem[110568] = 16'b0000000000000000;
	sram_mem[110569] = 16'b0000000000000000;
	sram_mem[110570] = 16'b0000000000000000;
	sram_mem[110571] = 16'b0000000000000000;
	sram_mem[110572] = 16'b0000000000000000;
	sram_mem[110573] = 16'b0000000000000000;
	sram_mem[110574] = 16'b0000000000000000;
	sram_mem[110575] = 16'b0000000000000000;
	sram_mem[110576] = 16'b0000000000000000;
	sram_mem[110577] = 16'b0000000000000000;
	sram_mem[110578] = 16'b0000000000000000;
	sram_mem[110579] = 16'b0000000000000000;
	sram_mem[110580] = 16'b0000000000000000;
	sram_mem[110581] = 16'b0000000000000000;
	sram_mem[110582] = 16'b0000000000000000;
	sram_mem[110583] = 16'b0000000000000000;
	sram_mem[110584] = 16'b0000000000000000;
	sram_mem[110585] = 16'b0000000000000000;
	sram_mem[110586] = 16'b0000000000000000;
	sram_mem[110587] = 16'b0000000000000000;
	sram_mem[110588] = 16'b0000000000000000;
	sram_mem[110589] = 16'b0000000000000000;
	sram_mem[110590] = 16'b0000000000000000;
	sram_mem[110591] = 16'b0000000000000000;
	sram_mem[110592] = 16'b0000000000000000;
	sram_mem[110593] = 16'b0000000000000000;
	sram_mem[110594] = 16'b0000000000000000;
	sram_mem[110595] = 16'b0000000000000000;
	sram_mem[110596] = 16'b0000000000000000;
	sram_mem[110597] = 16'b0000000000000000;
	sram_mem[110598] = 16'b0000000000000000;
	sram_mem[110599] = 16'b0000000000000000;
	sram_mem[110600] = 16'b0000000000000000;
	sram_mem[110601] = 16'b0000000000000000;
	sram_mem[110602] = 16'b0000000000000000;
	sram_mem[110603] = 16'b0000000000000000;
	sram_mem[110604] = 16'b0000000000000000;
	sram_mem[110605] = 16'b0000000000000000;
	sram_mem[110606] = 16'b0000000000000000;
	sram_mem[110607] = 16'b0000000000000000;
	sram_mem[110608] = 16'b0000000000000000;
	sram_mem[110609] = 16'b0000000000000000;
	sram_mem[110610] = 16'b0000000000000000;
	sram_mem[110611] = 16'b0000000000000000;
	sram_mem[110612] = 16'b0000000000000000;
	sram_mem[110613] = 16'b0000000000000000;
	sram_mem[110614] = 16'b0000000000000000;
	sram_mem[110615] = 16'b0000000000000000;
	sram_mem[110616] = 16'b0000000000000000;
	sram_mem[110617] = 16'b0000000000000000;
	sram_mem[110618] = 16'b0000000000000000;
	sram_mem[110619] = 16'b0000000000000000;
	sram_mem[110620] = 16'b0000000000000000;
	sram_mem[110621] = 16'b0000000000000000;
	sram_mem[110622] = 16'b0000000000000000;
	sram_mem[110623] = 16'b0000000000000000;
	sram_mem[110624] = 16'b0000000000000000;
	sram_mem[110625] = 16'b0000000000000000;
	sram_mem[110626] = 16'b0000000000000000;
	sram_mem[110627] = 16'b0000000000000000;
	sram_mem[110628] = 16'b0000000000000000;
	sram_mem[110629] = 16'b0000000000000000;
	sram_mem[110630] = 16'b0000000000000000;
	sram_mem[110631] = 16'b0000000000000000;
	sram_mem[110632] = 16'b0000000000000000;
	sram_mem[110633] = 16'b0000000000000000;
	sram_mem[110634] = 16'b0000000000000000;
	sram_mem[110635] = 16'b0000000000000000;
	sram_mem[110636] = 16'b0000000000000000;
	sram_mem[110637] = 16'b0000000000000000;
	sram_mem[110638] = 16'b0000000000000000;
	sram_mem[110639] = 16'b0000000000000000;
	sram_mem[110640] = 16'b0000000000000000;
	sram_mem[110641] = 16'b0000000000000000;
	sram_mem[110642] = 16'b0000000000000000;
	sram_mem[110643] = 16'b0000000000000000;
	sram_mem[110644] = 16'b0000000000000000;
	sram_mem[110645] = 16'b0000000000000000;
	sram_mem[110646] = 16'b0000000000000000;
	sram_mem[110647] = 16'b0000000000000000;
	sram_mem[110648] = 16'b0000000000000000;
	sram_mem[110649] = 16'b0000000000000000;
	sram_mem[110650] = 16'b0000000000000000;
	sram_mem[110651] = 16'b0000000000000000;
	sram_mem[110652] = 16'b0000000000000000;
	sram_mem[110653] = 16'b0000000000000000;
	sram_mem[110654] = 16'b0000000000000000;
	sram_mem[110655] = 16'b0000000000000000;
	sram_mem[110656] = 16'b0000000000000000;
	sram_mem[110657] = 16'b0000000000000000;
	sram_mem[110658] = 16'b0000000000000000;
	sram_mem[110659] = 16'b0000000000000000;
	sram_mem[110660] = 16'b0000000000000000;
	sram_mem[110661] = 16'b0000000000000000;
	sram_mem[110662] = 16'b0000000000000000;
	sram_mem[110663] = 16'b0000000000000000;
	sram_mem[110664] = 16'b0000000000000000;
	sram_mem[110665] = 16'b0000000000000000;
	sram_mem[110666] = 16'b0000000000000000;
	sram_mem[110667] = 16'b0000000000000000;
	sram_mem[110668] = 16'b0000000000000000;
	sram_mem[110669] = 16'b0000000000000000;
	sram_mem[110670] = 16'b0000000000000000;
	sram_mem[110671] = 16'b0000000000000000;
	sram_mem[110672] = 16'b0000000000000000;
	sram_mem[110673] = 16'b0000000000000000;
	sram_mem[110674] = 16'b0000000000000000;
	sram_mem[110675] = 16'b0000000000000000;
	sram_mem[110676] = 16'b0000000000000000;
	sram_mem[110677] = 16'b0000000000000000;
	sram_mem[110678] = 16'b0000000000000000;
	sram_mem[110679] = 16'b0000000000000000;
	sram_mem[110680] = 16'b0000000000000000;
	sram_mem[110681] = 16'b0000000000000000;
	sram_mem[110682] = 16'b0000000000000000;
	sram_mem[110683] = 16'b0000000000000000;
	sram_mem[110684] = 16'b0000000000000000;
	sram_mem[110685] = 16'b0000000000000000;
	sram_mem[110686] = 16'b0000000000000000;
	sram_mem[110687] = 16'b0000000000000000;
	sram_mem[110688] = 16'b0000000000000000;
	sram_mem[110689] = 16'b0000000000000000;
	sram_mem[110690] = 16'b0000000000000000;
	sram_mem[110691] = 16'b0000000000000000;
	sram_mem[110692] = 16'b0000000000000000;
	sram_mem[110693] = 16'b0000000000000000;
	sram_mem[110694] = 16'b0000000000000000;
	sram_mem[110695] = 16'b0000000000000000;
	sram_mem[110696] = 16'b0000000000000000;
	sram_mem[110697] = 16'b0000000000000000;
	sram_mem[110698] = 16'b0000000000000000;
	sram_mem[110699] = 16'b0000000000000000;
	sram_mem[110700] = 16'b0000000000000000;
	sram_mem[110701] = 16'b0000000000000000;
	sram_mem[110702] = 16'b0000000000000000;
	sram_mem[110703] = 16'b0000000000000000;
	sram_mem[110704] = 16'b0000000000000000;
	sram_mem[110705] = 16'b0000000000000000;
	sram_mem[110706] = 16'b0000000000000000;
	sram_mem[110707] = 16'b0000000000000000;
	sram_mem[110708] = 16'b0000000000000000;
	sram_mem[110709] = 16'b0000000000000000;
	sram_mem[110710] = 16'b0000000000000000;
	sram_mem[110711] = 16'b0000000000000000;
	sram_mem[110712] = 16'b0000000000000000;
	sram_mem[110713] = 16'b0000000000000000;
	sram_mem[110714] = 16'b0000000000000000;
	sram_mem[110715] = 16'b0000000000000000;
	sram_mem[110716] = 16'b0000000000000000;
	sram_mem[110717] = 16'b0000000000000000;
	sram_mem[110718] = 16'b0000000000000000;
	sram_mem[110719] = 16'b0000000000000000;
	sram_mem[110720] = 16'b0000000000000000;
	sram_mem[110721] = 16'b0000000000000000;
	sram_mem[110722] = 16'b0000000000000000;
	sram_mem[110723] = 16'b0000000000000000;
	sram_mem[110724] = 16'b0000000000000000;
	sram_mem[110725] = 16'b0000000000000000;
	sram_mem[110726] = 16'b0000000000000000;
	sram_mem[110727] = 16'b0000000000000000;
	sram_mem[110728] = 16'b0000000000000000;
	sram_mem[110729] = 16'b0000000000000000;
	sram_mem[110730] = 16'b0000000000000000;
	sram_mem[110731] = 16'b0000000000000000;
	sram_mem[110732] = 16'b0000000000000000;
	sram_mem[110733] = 16'b0000000000000000;
	sram_mem[110734] = 16'b0000000000000000;
	sram_mem[110735] = 16'b0000000000000000;
	sram_mem[110736] = 16'b0000000000000000;
	sram_mem[110737] = 16'b0000000000000000;
	sram_mem[110738] = 16'b0000000000000000;
	sram_mem[110739] = 16'b0000000000000000;
	sram_mem[110740] = 16'b0000000000000000;
	sram_mem[110741] = 16'b0000000000000000;
	sram_mem[110742] = 16'b0000000000000000;
	sram_mem[110743] = 16'b0000000000000000;
	sram_mem[110744] = 16'b0000000000000000;
	sram_mem[110745] = 16'b0000000000000000;
	sram_mem[110746] = 16'b0000000000000000;
	sram_mem[110747] = 16'b0000000000000000;
	sram_mem[110748] = 16'b0000000000000000;
	sram_mem[110749] = 16'b0000000000000000;
	sram_mem[110750] = 16'b0000000000000000;
	sram_mem[110751] = 16'b0000000000000000;
	sram_mem[110752] = 16'b0000000000000000;
	sram_mem[110753] = 16'b0000000000000000;
	sram_mem[110754] = 16'b0000000000000000;
	sram_mem[110755] = 16'b0000000000000000;
	sram_mem[110756] = 16'b0000000000000000;
	sram_mem[110757] = 16'b0000000000000000;
	sram_mem[110758] = 16'b0000000000000000;
	sram_mem[110759] = 16'b0000000000000000;
	sram_mem[110760] = 16'b0000000000000000;
	sram_mem[110761] = 16'b0000000000000000;
	sram_mem[110762] = 16'b0000000000000000;
	sram_mem[110763] = 16'b0000000000000000;
	sram_mem[110764] = 16'b0000000000000000;
	sram_mem[110765] = 16'b0000000000000000;
	sram_mem[110766] = 16'b0000000000000000;
	sram_mem[110767] = 16'b0000000000000000;
	sram_mem[110768] = 16'b0000000000000000;
	sram_mem[110769] = 16'b0000000000000000;
	sram_mem[110770] = 16'b0000000000000000;
	sram_mem[110771] = 16'b0000000000000000;
	sram_mem[110772] = 16'b0000000000000000;
	sram_mem[110773] = 16'b0000000000000000;
	sram_mem[110774] = 16'b0000000000000000;
	sram_mem[110775] = 16'b0000000000000000;
	sram_mem[110776] = 16'b0000000000000000;
	sram_mem[110777] = 16'b0000000000000000;
	sram_mem[110778] = 16'b0000000000000000;
	sram_mem[110779] = 16'b0000000000000000;
	sram_mem[110780] = 16'b0000000000000000;
	sram_mem[110781] = 16'b0000000000000000;
	sram_mem[110782] = 16'b0000000000000000;
	sram_mem[110783] = 16'b0000000000000000;
	sram_mem[110784] = 16'b0000000000000000;
	sram_mem[110785] = 16'b0000000000000000;
	sram_mem[110786] = 16'b0000000000000000;
	sram_mem[110787] = 16'b0000000000000000;
	sram_mem[110788] = 16'b0000000000000000;
	sram_mem[110789] = 16'b0000000000000000;
	sram_mem[110790] = 16'b0000000000000000;
	sram_mem[110791] = 16'b0000000000000000;
	sram_mem[110792] = 16'b0000000000000000;
	sram_mem[110793] = 16'b0000000000000000;
	sram_mem[110794] = 16'b0000000000000000;
	sram_mem[110795] = 16'b0000000000000000;
	sram_mem[110796] = 16'b0000000000000000;
	sram_mem[110797] = 16'b0000000000000000;
	sram_mem[110798] = 16'b0000000000000000;
	sram_mem[110799] = 16'b0000000000000000;
	sram_mem[110800] = 16'b0000000000000000;
	sram_mem[110801] = 16'b0000000000000000;
	sram_mem[110802] = 16'b0000000000000000;
	sram_mem[110803] = 16'b0000000000000000;
	sram_mem[110804] = 16'b0000000000000000;
	sram_mem[110805] = 16'b0000000000000000;
	sram_mem[110806] = 16'b0000000000000000;
	sram_mem[110807] = 16'b0000000000000000;
	sram_mem[110808] = 16'b0000000000000000;
	sram_mem[110809] = 16'b0000000000000000;
	sram_mem[110810] = 16'b0000000000000000;
	sram_mem[110811] = 16'b0000000000000000;
	sram_mem[110812] = 16'b0000000000000000;
	sram_mem[110813] = 16'b0000000000000000;
	sram_mem[110814] = 16'b0000000000000000;
	sram_mem[110815] = 16'b0000000000000000;
	sram_mem[110816] = 16'b0000000000000000;
	sram_mem[110817] = 16'b0000000000000000;
	sram_mem[110818] = 16'b0000000000000000;
	sram_mem[110819] = 16'b0000000000000000;
	sram_mem[110820] = 16'b0000000000000000;
	sram_mem[110821] = 16'b0000000000000000;
	sram_mem[110822] = 16'b0000000000000000;
	sram_mem[110823] = 16'b0000000000000000;
	sram_mem[110824] = 16'b0000000000000000;
	sram_mem[110825] = 16'b0000000000000000;
	sram_mem[110826] = 16'b0000000000000000;
	sram_mem[110827] = 16'b0000000000000000;
	sram_mem[110828] = 16'b0000000000000000;
	sram_mem[110829] = 16'b0000000000000000;
	sram_mem[110830] = 16'b0000000000000000;
	sram_mem[110831] = 16'b0000000000000000;
	sram_mem[110832] = 16'b0000000000000000;
	sram_mem[110833] = 16'b0000000000000000;
	sram_mem[110834] = 16'b0000000000000000;
	sram_mem[110835] = 16'b0000000000000000;
	sram_mem[110836] = 16'b0000000000000000;
	sram_mem[110837] = 16'b0000000000000000;
	sram_mem[110838] = 16'b0000000000000000;
	sram_mem[110839] = 16'b0000000000000000;
	sram_mem[110840] = 16'b0000000000000000;
	sram_mem[110841] = 16'b0000000000000000;
	sram_mem[110842] = 16'b0000000000000000;
	sram_mem[110843] = 16'b0000000000000000;
	sram_mem[110844] = 16'b0000000000000000;
	sram_mem[110845] = 16'b0000000000000000;
	sram_mem[110846] = 16'b0000000000000000;
	sram_mem[110847] = 16'b0000000000000000;
	sram_mem[110848] = 16'b0000000000000000;
	sram_mem[110849] = 16'b0000000000000000;
	sram_mem[110850] = 16'b0000000000000000;
	sram_mem[110851] = 16'b0000000000000000;
	sram_mem[110852] = 16'b0000000000000000;
	sram_mem[110853] = 16'b0000000000000000;
	sram_mem[110854] = 16'b0000000000000000;
	sram_mem[110855] = 16'b0000000000000000;
	sram_mem[110856] = 16'b0000000000000000;
	sram_mem[110857] = 16'b0000000000000000;
	sram_mem[110858] = 16'b0000000000000000;
	sram_mem[110859] = 16'b0000000000000000;
	sram_mem[110860] = 16'b0000000000000000;
	sram_mem[110861] = 16'b0000000000000000;
	sram_mem[110862] = 16'b0000000000000000;
	sram_mem[110863] = 16'b0000000000000000;
	sram_mem[110864] = 16'b0000000000000000;
	sram_mem[110865] = 16'b0000000000000000;
	sram_mem[110866] = 16'b0000000000000000;
	sram_mem[110867] = 16'b0000000000000000;
	sram_mem[110868] = 16'b0000000000000000;
	sram_mem[110869] = 16'b0000000000000000;
	sram_mem[110870] = 16'b0000000000000000;
	sram_mem[110871] = 16'b0000000000000000;
	sram_mem[110872] = 16'b0000000000000000;
	sram_mem[110873] = 16'b0000000000000000;
	sram_mem[110874] = 16'b0000000000000000;
	sram_mem[110875] = 16'b0000000000000000;
	sram_mem[110876] = 16'b0000000000000000;
	sram_mem[110877] = 16'b0000000000000000;
	sram_mem[110878] = 16'b0000000000000000;
	sram_mem[110879] = 16'b0000000000000000;
	sram_mem[110880] = 16'b0000000000000000;
	sram_mem[110881] = 16'b0000000000000000;
	sram_mem[110882] = 16'b0000000000000000;
	sram_mem[110883] = 16'b0000000000000000;
	sram_mem[110884] = 16'b0000000000000000;
	sram_mem[110885] = 16'b0000000000000000;
	sram_mem[110886] = 16'b0000000000000000;
	sram_mem[110887] = 16'b0000000000000000;
	sram_mem[110888] = 16'b0000000000000000;
	sram_mem[110889] = 16'b0000000000000000;
	sram_mem[110890] = 16'b0000000000000000;
	sram_mem[110891] = 16'b0000000000000000;
	sram_mem[110892] = 16'b0000000000000000;
	sram_mem[110893] = 16'b0000000000000000;
	sram_mem[110894] = 16'b0000000000000000;
	sram_mem[110895] = 16'b0000000000000000;
	sram_mem[110896] = 16'b0000000000000000;
	sram_mem[110897] = 16'b0000000000000000;
	sram_mem[110898] = 16'b0000000000000000;
	sram_mem[110899] = 16'b0000000000000000;
	sram_mem[110900] = 16'b0000000000000000;
	sram_mem[110901] = 16'b0000000000000000;
	sram_mem[110902] = 16'b0000000000000000;
	sram_mem[110903] = 16'b0000000000000000;
	sram_mem[110904] = 16'b0000000000000000;
	sram_mem[110905] = 16'b0000000000000000;
	sram_mem[110906] = 16'b0000000000000000;
	sram_mem[110907] = 16'b0000000000000000;
	sram_mem[110908] = 16'b0000000000000000;
	sram_mem[110909] = 16'b0000000000000000;
	sram_mem[110910] = 16'b0000000000000000;
	sram_mem[110911] = 16'b0000000000000000;
	sram_mem[110912] = 16'b0000000000000000;
	sram_mem[110913] = 16'b0000000000000000;
	sram_mem[110914] = 16'b0000000000000000;
	sram_mem[110915] = 16'b0000000000000000;
	sram_mem[110916] = 16'b0000000000000000;
	sram_mem[110917] = 16'b0000000000000000;
	sram_mem[110918] = 16'b0000000000000000;
	sram_mem[110919] = 16'b0000000000000000;
	sram_mem[110920] = 16'b0000000000000000;
	sram_mem[110921] = 16'b0000000000000000;
	sram_mem[110922] = 16'b0000000000000000;
	sram_mem[110923] = 16'b0000000000000000;
	sram_mem[110924] = 16'b0000000000000000;
	sram_mem[110925] = 16'b0000000000000000;
	sram_mem[110926] = 16'b0000000000000000;
	sram_mem[110927] = 16'b0000000000000000;
	sram_mem[110928] = 16'b0000000000000000;
	sram_mem[110929] = 16'b0000000000000000;
	sram_mem[110930] = 16'b0000000000000000;
	sram_mem[110931] = 16'b0000000000000000;
	sram_mem[110932] = 16'b0000000000000000;
	sram_mem[110933] = 16'b0000000000000000;
	sram_mem[110934] = 16'b0000000000000000;
	sram_mem[110935] = 16'b0000000000000000;
	sram_mem[110936] = 16'b0000000000000000;
	sram_mem[110937] = 16'b0000000000000000;
	sram_mem[110938] = 16'b0000000000000000;
	sram_mem[110939] = 16'b0000000000000000;
	sram_mem[110940] = 16'b0000000000000000;
	sram_mem[110941] = 16'b0000000000000000;
	sram_mem[110942] = 16'b0000000000000000;
	sram_mem[110943] = 16'b0000000000000000;
	sram_mem[110944] = 16'b0000000000000000;
	sram_mem[110945] = 16'b0000000000000000;
	sram_mem[110946] = 16'b0000000000000000;
	sram_mem[110947] = 16'b0000000000000000;
	sram_mem[110948] = 16'b0000000000000000;
	sram_mem[110949] = 16'b0000000000000000;
	sram_mem[110950] = 16'b0000000000000000;
	sram_mem[110951] = 16'b0000000000000000;
	sram_mem[110952] = 16'b0000000000000000;
	sram_mem[110953] = 16'b0000000000000000;
	sram_mem[110954] = 16'b0000000000000000;
	sram_mem[110955] = 16'b0000000000000000;
	sram_mem[110956] = 16'b0000000000000000;
	sram_mem[110957] = 16'b0000000000000000;
	sram_mem[110958] = 16'b0000000000000000;
	sram_mem[110959] = 16'b0000000000000000;
	sram_mem[110960] = 16'b0000000000000000;
	sram_mem[110961] = 16'b0000000000000000;
	sram_mem[110962] = 16'b0000000000000000;
	sram_mem[110963] = 16'b0000000000000000;
	sram_mem[110964] = 16'b0000000000000000;
	sram_mem[110965] = 16'b0000000000000000;
	sram_mem[110966] = 16'b0000000000000000;
	sram_mem[110967] = 16'b0000000000000000;
	sram_mem[110968] = 16'b0000000000000000;
	sram_mem[110969] = 16'b0000000000000000;
	sram_mem[110970] = 16'b0000000000000000;
	sram_mem[110971] = 16'b0000000000000000;
	sram_mem[110972] = 16'b0000000000000000;
	sram_mem[110973] = 16'b0000000000000000;
	sram_mem[110974] = 16'b0000000000000000;
	sram_mem[110975] = 16'b0000000000000000;
	sram_mem[110976] = 16'b0000000000000000;
	sram_mem[110977] = 16'b0000000000000000;
	sram_mem[110978] = 16'b0000000000000000;
	sram_mem[110979] = 16'b0000000000000000;
	sram_mem[110980] = 16'b0000000000000000;
	sram_mem[110981] = 16'b0000000000000000;
	sram_mem[110982] = 16'b0000000000000000;
	sram_mem[110983] = 16'b0000000000000000;
	sram_mem[110984] = 16'b0000000000000000;
	sram_mem[110985] = 16'b0000000000000000;
	sram_mem[110986] = 16'b0000000000000000;
	sram_mem[110987] = 16'b0000000000000000;
	sram_mem[110988] = 16'b0000000000000000;
	sram_mem[110989] = 16'b0000000000000000;
	sram_mem[110990] = 16'b0000000000000000;
	sram_mem[110991] = 16'b0000000000000000;
	sram_mem[110992] = 16'b0000000000000000;
	sram_mem[110993] = 16'b0000000000000000;
	sram_mem[110994] = 16'b0000000000000000;
	sram_mem[110995] = 16'b0000000000000000;
	sram_mem[110996] = 16'b0000000000000000;
	sram_mem[110997] = 16'b0000000000000000;
	sram_mem[110998] = 16'b0000000000000000;
	sram_mem[110999] = 16'b0000000000000000;
	sram_mem[111000] = 16'b0000000000000000;
	sram_mem[111001] = 16'b0000000000000000;
	sram_mem[111002] = 16'b0000000000000000;
	sram_mem[111003] = 16'b0000000000000000;
	sram_mem[111004] = 16'b0000000000000000;
	sram_mem[111005] = 16'b0000000000000000;
	sram_mem[111006] = 16'b0000000000000000;
	sram_mem[111007] = 16'b0000000000000000;
	sram_mem[111008] = 16'b0000000000000000;
	sram_mem[111009] = 16'b0000000000000000;
	sram_mem[111010] = 16'b0000000000000000;
	sram_mem[111011] = 16'b0000000000000000;
	sram_mem[111012] = 16'b0000000000000000;
	sram_mem[111013] = 16'b0000000000000000;
	sram_mem[111014] = 16'b0000000000000000;
	sram_mem[111015] = 16'b0000000000000000;
	sram_mem[111016] = 16'b0000000000000000;
	sram_mem[111017] = 16'b0000000000000000;
	sram_mem[111018] = 16'b0000000000000000;
	sram_mem[111019] = 16'b0000000000000000;
	sram_mem[111020] = 16'b0000000000000000;
	sram_mem[111021] = 16'b0000000000000000;
	sram_mem[111022] = 16'b0000000000000000;
	sram_mem[111023] = 16'b0000000000000000;
	sram_mem[111024] = 16'b0000000000000000;
	sram_mem[111025] = 16'b0000000000000000;
	sram_mem[111026] = 16'b0000000000000000;
	sram_mem[111027] = 16'b0000000000000000;
	sram_mem[111028] = 16'b0000000000000000;
	sram_mem[111029] = 16'b0000000000000000;
	sram_mem[111030] = 16'b0000000000000000;
	sram_mem[111031] = 16'b0000000000000000;
	sram_mem[111032] = 16'b0000000000000000;
	sram_mem[111033] = 16'b0000000000000000;
	sram_mem[111034] = 16'b0000000000000000;
	sram_mem[111035] = 16'b0000000000000000;
	sram_mem[111036] = 16'b0000000000000000;
	sram_mem[111037] = 16'b0000000000000000;
	sram_mem[111038] = 16'b0000000000000000;
	sram_mem[111039] = 16'b0000000000000000;
	sram_mem[111040] = 16'b0000000000000000;
	sram_mem[111041] = 16'b0000000000000000;
	sram_mem[111042] = 16'b0000000000000000;
	sram_mem[111043] = 16'b0000000000000000;
	sram_mem[111044] = 16'b0000000000000000;
	sram_mem[111045] = 16'b0000000000000000;
	sram_mem[111046] = 16'b0000000000000000;
	sram_mem[111047] = 16'b0000000000000000;
	sram_mem[111048] = 16'b0000000000000000;
	sram_mem[111049] = 16'b0000000000000000;
	sram_mem[111050] = 16'b0000000000000000;
	sram_mem[111051] = 16'b0000000000000000;
	sram_mem[111052] = 16'b0000000000000000;
	sram_mem[111053] = 16'b0000000000000000;
	sram_mem[111054] = 16'b0000000000000000;
	sram_mem[111055] = 16'b0000000000000000;
	sram_mem[111056] = 16'b0000000000000000;
	sram_mem[111057] = 16'b0000000000000000;
	sram_mem[111058] = 16'b0000000000000000;
	sram_mem[111059] = 16'b0000000000000000;
	sram_mem[111060] = 16'b0000000000000000;
	sram_mem[111061] = 16'b0000000000000000;
	sram_mem[111062] = 16'b0000000000000000;
	sram_mem[111063] = 16'b0000000000000000;
	sram_mem[111064] = 16'b0000000000000000;
	sram_mem[111065] = 16'b0000000000000000;
	sram_mem[111066] = 16'b0000000000000000;
	sram_mem[111067] = 16'b0000000000000000;
	sram_mem[111068] = 16'b0000000000000000;
	sram_mem[111069] = 16'b0000000000000000;
	sram_mem[111070] = 16'b0000000000000000;
	sram_mem[111071] = 16'b0000000000000000;
	sram_mem[111072] = 16'b0000000000000000;
	sram_mem[111073] = 16'b0000000000000000;
	sram_mem[111074] = 16'b0000000000000000;
	sram_mem[111075] = 16'b0000000000000000;
	sram_mem[111076] = 16'b0000000000000000;
	sram_mem[111077] = 16'b0000000000000000;
	sram_mem[111078] = 16'b0000000000000000;
	sram_mem[111079] = 16'b0000000000000000;
	sram_mem[111080] = 16'b0000000000000000;
	sram_mem[111081] = 16'b0000000000000000;
	sram_mem[111082] = 16'b0000000000000000;
	sram_mem[111083] = 16'b0000000000000000;
	sram_mem[111084] = 16'b0000000000000000;
	sram_mem[111085] = 16'b0000000000000000;
	sram_mem[111086] = 16'b0000000000000000;
	sram_mem[111087] = 16'b0000000000000000;
	sram_mem[111088] = 16'b0000000000000000;
	sram_mem[111089] = 16'b0000000000000000;
	sram_mem[111090] = 16'b0000000000000000;
	sram_mem[111091] = 16'b0000000000000000;
	sram_mem[111092] = 16'b0000000000000000;
	sram_mem[111093] = 16'b0000000000000000;
	sram_mem[111094] = 16'b0000000000000000;
	sram_mem[111095] = 16'b0000000000000000;
	sram_mem[111096] = 16'b0000000000000000;
	sram_mem[111097] = 16'b0000000000000000;
	sram_mem[111098] = 16'b0000000000000000;
	sram_mem[111099] = 16'b0000000000000000;
	sram_mem[111100] = 16'b0000000000000000;
	sram_mem[111101] = 16'b0000000000000000;
	sram_mem[111102] = 16'b0000000000000000;
	sram_mem[111103] = 16'b0000000000000000;
	sram_mem[111104] = 16'b0000000000000000;
	sram_mem[111105] = 16'b0000000000000000;
	sram_mem[111106] = 16'b0000000000000000;
	sram_mem[111107] = 16'b0000000000000000;
	sram_mem[111108] = 16'b0000000000000000;
	sram_mem[111109] = 16'b0000000000000000;
	sram_mem[111110] = 16'b0000000000000000;
	sram_mem[111111] = 16'b0000000000000000;
	sram_mem[111112] = 16'b0000000000000000;
	sram_mem[111113] = 16'b0000000000000000;
	sram_mem[111114] = 16'b0000000000000000;
	sram_mem[111115] = 16'b0000000000000000;
	sram_mem[111116] = 16'b0000000000000000;
	sram_mem[111117] = 16'b0000000000000000;
	sram_mem[111118] = 16'b0000000000000000;
	sram_mem[111119] = 16'b0000000000000000;
	sram_mem[111120] = 16'b0000000000000000;
	sram_mem[111121] = 16'b0000000000000000;
	sram_mem[111122] = 16'b0000000000000000;
	sram_mem[111123] = 16'b0000000000000000;
	sram_mem[111124] = 16'b0000000000000000;
	sram_mem[111125] = 16'b0000000000000000;
	sram_mem[111126] = 16'b0000000000000000;
	sram_mem[111127] = 16'b0000000000000000;
	sram_mem[111128] = 16'b0000000000000000;
	sram_mem[111129] = 16'b0000000000000000;
	sram_mem[111130] = 16'b0000000000000000;
	sram_mem[111131] = 16'b0000000000000000;
	sram_mem[111132] = 16'b0000000000000000;
	sram_mem[111133] = 16'b0000000000000000;
	sram_mem[111134] = 16'b0000000000000000;
	sram_mem[111135] = 16'b0000000000000000;
	sram_mem[111136] = 16'b0000000000000000;
	sram_mem[111137] = 16'b0000000000000000;
	sram_mem[111138] = 16'b0000000000000000;
	sram_mem[111139] = 16'b0000000000000000;
	sram_mem[111140] = 16'b0000000000000000;
	sram_mem[111141] = 16'b0000000000000000;
	sram_mem[111142] = 16'b0000000000000000;
	sram_mem[111143] = 16'b0000000000000000;
	sram_mem[111144] = 16'b0000000000000000;
	sram_mem[111145] = 16'b0000000000000000;
	sram_mem[111146] = 16'b0000000000000000;
	sram_mem[111147] = 16'b0000000000000000;
	sram_mem[111148] = 16'b0000000000000000;
	sram_mem[111149] = 16'b0000000000000000;
	sram_mem[111150] = 16'b0000000000000000;
	sram_mem[111151] = 16'b0000000000000000;
	sram_mem[111152] = 16'b0000000000000000;
	sram_mem[111153] = 16'b0000000000000000;
	sram_mem[111154] = 16'b0000000000000000;
	sram_mem[111155] = 16'b0000000000000000;
	sram_mem[111156] = 16'b0000000000000000;
	sram_mem[111157] = 16'b0000000000000000;
	sram_mem[111158] = 16'b0000000000000000;
	sram_mem[111159] = 16'b0000000000000000;
	sram_mem[111160] = 16'b0000000000000000;
	sram_mem[111161] = 16'b0000000000000000;
	sram_mem[111162] = 16'b0000000000000000;
	sram_mem[111163] = 16'b0000000000000000;
	sram_mem[111164] = 16'b0000000000000000;
	sram_mem[111165] = 16'b0000000000000000;
	sram_mem[111166] = 16'b0000000000000000;
	sram_mem[111167] = 16'b0000000000000000;
	sram_mem[111168] = 16'b0000000000000000;
	sram_mem[111169] = 16'b0000000000000000;
	sram_mem[111170] = 16'b0000000000000000;
	sram_mem[111171] = 16'b0000000000000000;
	sram_mem[111172] = 16'b0000000000000000;
	sram_mem[111173] = 16'b0000000000000000;
	sram_mem[111174] = 16'b0000000000000000;
	sram_mem[111175] = 16'b0000000000000000;
	sram_mem[111176] = 16'b0000000000000000;
	sram_mem[111177] = 16'b0000000000000000;
	sram_mem[111178] = 16'b0000000000000000;
	sram_mem[111179] = 16'b0000000000000000;
	sram_mem[111180] = 16'b0000000000000000;
	sram_mem[111181] = 16'b0000000000000000;
	sram_mem[111182] = 16'b0000000000000000;
	sram_mem[111183] = 16'b0000000000000000;
	sram_mem[111184] = 16'b0000000000000000;
	sram_mem[111185] = 16'b0000000000000000;
	sram_mem[111186] = 16'b0000000000000000;
	sram_mem[111187] = 16'b0000000000000000;
	sram_mem[111188] = 16'b0000000000000000;
	sram_mem[111189] = 16'b0000000000000000;
	sram_mem[111190] = 16'b0000000000000000;
	sram_mem[111191] = 16'b0000000000000000;
	sram_mem[111192] = 16'b0000000000000000;
	sram_mem[111193] = 16'b0000000000000000;
	sram_mem[111194] = 16'b0000000000000000;
	sram_mem[111195] = 16'b0000000000000000;
	sram_mem[111196] = 16'b0000000000000000;
	sram_mem[111197] = 16'b0000000000000000;
	sram_mem[111198] = 16'b0000000000000000;
	sram_mem[111199] = 16'b0000000000000000;
	sram_mem[111200] = 16'b0000000000000000;
	sram_mem[111201] = 16'b0000000000000000;
	sram_mem[111202] = 16'b0000000000000000;
	sram_mem[111203] = 16'b0000000000000000;
	sram_mem[111204] = 16'b0000000000000000;
	sram_mem[111205] = 16'b0000000000000000;
	sram_mem[111206] = 16'b0000000000000000;
	sram_mem[111207] = 16'b0000000000000000;
	sram_mem[111208] = 16'b0000000000000000;
	sram_mem[111209] = 16'b0000000000000000;
	sram_mem[111210] = 16'b0000000000000000;
	sram_mem[111211] = 16'b0000000000000000;
	sram_mem[111212] = 16'b0000000000000000;
	sram_mem[111213] = 16'b0000000000000000;
	sram_mem[111214] = 16'b0000000000000000;
	sram_mem[111215] = 16'b0000000000000000;
	sram_mem[111216] = 16'b0000000000000000;
	sram_mem[111217] = 16'b0000000000000000;
	sram_mem[111218] = 16'b0000000000000000;
	sram_mem[111219] = 16'b0000000000000000;
	sram_mem[111220] = 16'b0000000000000000;
	sram_mem[111221] = 16'b0000000000000000;
	sram_mem[111222] = 16'b0000000000000000;
	sram_mem[111223] = 16'b0000000000000000;
	sram_mem[111224] = 16'b0000000000000000;
	sram_mem[111225] = 16'b0000000000000000;
	sram_mem[111226] = 16'b0000000000000000;
	sram_mem[111227] = 16'b0000000000000000;
	sram_mem[111228] = 16'b0000000000000000;
	sram_mem[111229] = 16'b0000000000000000;
	sram_mem[111230] = 16'b0000000000000000;
	sram_mem[111231] = 16'b0000000000000000;
	sram_mem[111232] = 16'b0000000000000000;
	sram_mem[111233] = 16'b0000000000000000;
	sram_mem[111234] = 16'b0000000000000000;
	sram_mem[111235] = 16'b0000000000000000;
	sram_mem[111236] = 16'b0000000000000000;
	sram_mem[111237] = 16'b0000000000000000;
	sram_mem[111238] = 16'b0000000000000000;
	sram_mem[111239] = 16'b0000000000000000;
	sram_mem[111240] = 16'b0000000000000000;
	sram_mem[111241] = 16'b0000000000000000;
	sram_mem[111242] = 16'b0000000000000000;
	sram_mem[111243] = 16'b0000000000000000;
	sram_mem[111244] = 16'b0000000000000000;
	sram_mem[111245] = 16'b0000000000000000;
	sram_mem[111246] = 16'b0000000000000000;
	sram_mem[111247] = 16'b0000000000000000;
	sram_mem[111248] = 16'b0000000000000000;
	sram_mem[111249] = 16'b0000000000000000;
	sram_mem[111250] = 16'b0000000000000000;
	sram_mem[111251] = 16'b0000000000000000;
	sram_mem[111252] = 16'b0000000000000000;
	sram_mem[111253] = 16'b0000000000000000;
	sram_mem[111254] = 16'b0000000000000000;
	sram_mem[111255] = 16'b0000000000000000;
	sram_mem[111256] = 16'b0000000000000000;
	sram_mem[111257] = 16'b0000000000000000;
	sram_mem[111258] = 16'b0000000000000000;
	sram_mem[111259] = 16'b0000000000000000;
	sram_mem[111260] = 16'b0000000000000000;
	sram_mem[111261] = 16'b0000000000000000;
	sram_mem[111262] = 16'b0000000000000000;
	sram_mem[111263] = 16'b0000000000000000;
	sram_mem[111264] = 16'b0000000000000000;
	sram_mem[111265] = 16'b0000000000000000;
	sram_mem[111266] = 16'b0000000000000000;
	sram_mem[111267] = 16'b0000000000000000;
	sram_mem[111268] = 16'b0000000000000000;
	sram_mem[111269] = 16'b0000000000000000;
	sram_mem[111270] = 16'b0000000000000000;
	sram_mem[111271] = 16'b0000000000000000;
	sram_mem[111272] = 16'b0000000000000000;
	sram_mem[111273] = 16'b0000000000000000;
	sram_mem[111274] = 16'b0000000000000000;
	sram_mem[111275] = 16'b0000000000000000;
	sram_mem[111276] = 16'b0000000000000000;
	sram_mem[111277] = 16'b0000000000000000;
	sram_mem[111278] = 16'b0000000000000000;
	sram_mem[111279] = 16'b0000000000000000;
	sram_mem[111280] = 16'b0000000000000000;
	sram_mem[111281] = 16'b0000000000000000;
	sram_mem[111282] = 16'b0000000000000000;
	sram_mem[111283] = 16'b0000000000000000;
	sram_mem[111284] = 16'b0000000000000000;
	sram_mem[111285] = 16'b0000000000000000;
	sram_mem[111286] = 16'b0000000000000000;
	sram_mem[111287] = 16'b0000000000000000;
	sram_mem[111288] = 16'b0000000000000000;
	sram_mem[111289] = 16'b0000000000000000;
	sram_mem[111290] = 16'b0000000000000000;
	sram_mem[111291] = 16'b0000000000000000;
	sram_mem[111292] = 16'b0000000000000000;
	sram_mem[111293] = 16'b0000000000000000;
	sram_mem[111294] = 16'b0000000000000000;
	sram_mem[111295] = 16'b0000000000000000;
	sram_mem[111296] = 16'b0000000000000000;
	sram_mem[111297] = 16'b0000000000000000;
	sram_mem[111298] = 16'b0000000000000000;
	sram_mem[111299] = 16'b0000000000000000;
	sram_mem[111300] = 16'b0000000000000000;
	sram_mem[111301] = 16'b0000000000000000;
	sram_mem[111302] = 16'b0000000000000000;
	sram_mem[111303] = 16'b0000000000000000;
	sram_mem[111304] = 16'b0000000000000000;
	sram_mem[111305] = 16'b0000000000000000;
	sram_mem[111306] = 16'b0000000000000000;
	sram_mem[111307] = 16'b0000000000000000;
	sram_mem[111308] = 16'b0000000000000000;
	sram_mem[111309] = 16'b0000000000000000;
	sram_mem[111310] = 16'b0000000000000000;
	sram_mem[111311] = 16'b0000000000000000;
	sram_mem[111312] = 16'b0000000000000000;
	sram_mem[111313] = 16'b0000000000000000;
	sram_mem[111314] = 16'b0000000000000000;
	sram_mem[111315] = 16'b0000000000000000;
	sram_mem[111316] = 16'b0000000000000000;
	sram_mem[111317] = 16'b0000000000000000;
	sram_mem[111318] = 16'b0000000000000000;
	sram_mem[111319] = 16'b0000000000000000;
	sram_mem[111320] = 16'b0000000000000000;
	sram_mem[111321] = 16'b0000000000000000;
	sram_mem[111322] = 16'b0000000000000000;
	sram_mem[111323] = 16'b0000000000000000;
	sram_mem[111324] = 16'b0000000000000000;
	sram_mem[111325] = 16'b0000000000000000;
	sram_mem[111326] = 16'b0000000000000000;
	sram_mem[111327] = 16'b0000000000000000;
	sram_mem[111328] = 16'b0000000000000000;
	sram_mem[111329] = 16'b0000000000000000;
	sram_mem[111330] = 16'b0000000000000000;
	sram_mem[111331] = 16'b0000000000000000;
	sram_mem[111332] = 16'b0000000000000000;
	sram_mem[111333] = 16'b0000000000000000;
	sram_mem[111334] = 16'b0000000000000000;
	sram_mem[111335] = 16'b0000000000000000;
	sram_mem[111336] = 16'b0000000000000000;
	sram_mem[111337] = 16'b0000000000000000;
	sram_mem[111338] = 16'b0000000000000000;
	sram_mem[111339] = 16'b0000000000000000;
	sram_mem[111340] = 16'b0000000000000000;
	sram_mem[111341] = 16'b0000000000000000;
	sram_mem[111342] = 16'b0000000000000000;
	sram_mem[111343] = 16'b0000000000000000;
	sram_mem[111344] = 16'b0000000000000000;
	sram_mem[111345] = 16'b0000000000000000;
	sram_mem[111346] = 16'b0000000000000000;
	sram_mem[111347] = 16'b0000000000000000;
	sram_mem[111348] = 16'b0000000000000000;
	sram_mem[111349] = 16'b0000000000000000;
	sram_mem[111350] = 16'b0000000000000000;
	sram_mem[111351] = 16'b0000000000000000;
	sram_mem[111352] = 16'b0000000000000000;
	sram_mem[111353] = 16'b0000000000000000;
	sram_mem[111354] = 16'b0000000000000000;
	sram_mem[111355] = 16'b0000000000000000;
	sram_mem[111356] = 16'b0000000000000000;
	sram_mem[111357] = 16'b0000000000000000;
	sram_mem[111358] = 16'b0000000000000000;
	sram_mem[111359] = 16'b0000000000000000;
	sram_mem[111360] = 16'b0000000000000000;
	sram_mem[111361] = 16'b0000000000000000;
	sram_mem[111362] = 16'b0000000000000000;
	sram_mem[111363] = 16'b0000000000000000;
	sram_mem[111364] = 16'b0000000000000000;
	sram_mem[111365] = 16'b0000000000000000;
	sram_mem[111366] = 16'b0000000000000000;
	sram_mem[111367] = 16'b0000000000000000;
	sram_mem[111368] = 16'b0000000000000000;
	sram_mem[111369] = 16'b0000000000000000;
	sram_mem[111370] = 16'b0000000000000000;
	sram_mem[111371] = 16'b0000000000000000;
	sram_mem[111372] = 16'b0000000000000000;
	sram_mem[111373] = 16'b0000000000000000;
	sram_mem[111374] = 16'b0000000000000000;
	sram_mem[111375] = 16'b0000000000000000;
	sram_mem[111376] = 16'b0000000000000000;
	sram_mem[111377] = 16'b0000000000000000;
	sram_mem[111378] = 16'b0000000000000000;
	sram_mem[111379] = 16'b0000000000000000;
	sram_mem[111380] = 16'b0000000000000000;
	sram_mem[111381] = 16'b0000000000000000;
	sram_mem[111382] = 16'b0000000000000000;
	sram_mem[111383] = 16'b0000000000000000;
	sram_mem[111384] = 16'b0000000000000000;
	sram_mem[111385] = 16'b0000000000000000;
	sram_mem[111386] = 16'b0000000000000000;
	sram_mem[111387] = 16'b0000000000000000;
	sram_mem[111388] = 16'b0000000000000000;
	sram_mem[111389] = 16'b0000000000000000;
	sram_mem[111390] = 16'b0000000000000000;
	sram_mem[111391] = 16'b0000000000000000;
	sram_mem[111392] = 16'b0000000000000000;
	sram_mem[111393] = 16'b0000000000000000;
	sram_mem[111394] = 16'b0000000000000000;
	sram_mem[111395] = 16'b0000000000000000;
	sram_mem[111396] = 16'b0000000000000000;
	sram_mem[111397] = 16'b0000000000000000;
	sram_mem[111398] = 16'b0000000000000000;
	sram_mem[111399] = 16'b0000000000000000;
	sram_mem[111400] = 16'b0000000000000000;
	sram_mem[111401] = 16'b0000000000000000;
	sram_mem[111402] = 16'b0000000000000000;
	sram_mem[111403] = 16'b0000000000000000;
	sram_mem[111404] = 16'b0000000000000000;
	sram_mem[111405] = 16'b0000000000000000;
	sram_mem[111406] = 16'b0000000000000000;
	sram_mem[111407] = 16'b0000000000000000;
	sram_mem[111408] = 16'b0000000000000000;
	sram_mem[111409] = 16'b0000000000000000;
	sram_mem[111410] = 16'b0000000000000000;
	sram_mem[111411] = 16'b0000000000000000;
	sram_mem[111412] = 16'b0000000000000000;
	sram_mem[111413] = 16'b0000000000000000;
	sram_mem[111414] = 16'b0000000000000000;
	sram_mem[111415] = 16'b0000000000000000;
	sram_mem[111416] = 16'b0000000000000000;
	sram_mem[111417] = 16'b0000000000000000;
	sram_mem[111418] = 16'b0000000000000000;
	sram_mem[111419] = 16'b0000000000000000;
	sram_mem[111420] = 16'b0000000000000000;
	sram_mem[111421] = 16'b0000000000000000;
	sram_mem[111422] = 16'b0000000000000000;
	sram_mem[111423] = 16'b0000000000000000;
	sram_mem[111424] = 16'b0000000000000000;
	sram_mem[111425] = 16'b0000000000000000;
	sram_mem[111426] = 16'b0000000000000000;
	sram_mem[111427] = 16'b0000000000000000;
	sram_mem[111428] = 16'b0000000000000000;
	sram_mem[111429] = 16'b0000000000000000;
	sram_mem[111430] = 16'b0000000000000000;
	sram_mem[111431] = 16'b0000000000000000;
	sram_mem[111432] = 16'b0000000000000000;
	sram_mem[111433] = 16'b0000000000000000;
	sram_mem[111434] = 16'b0000000000000000;
	sram_mem[111435] = 16'b0000000000000000;
	sram_mem[111436] = 16'b0000000000000000;
	sram_mem[111437] = 16'b0000000000000000;
	sram_mem[111438] = 16'b0000000000000000;
	sram_mem[111439] = 16'b0000000000000000;
	sram_mem[111440] = 16'b0000000000000000;
	sram_mem[111441] = 16'b0000000000000000;
	sram_mem[111442] = 16'b0000000000000000;
	sram_mem[111443] = 16'b0000000000000000;
	sram_mem[111444] = 16'b0000000000000000;
	sram_mem[111445] = 16'b0000000000000000;
	sram_mem[111446] = 16'b0000000000000000;
	sram_mem[111447] = 16'b0000000000000000;
	sram_mem[111448] = 16'b0000000000000000;
	sram_mem[111449] = 16'b0000000000000000;
	sram_mem[111450] = 16'b0000000000000000;
	sram_mem[111451] = 16'b0000000000000000;
	sram_mem[111452] = 16'b0000000000000000;
	sram_mem[111453] = 16'b0000000000000000;
	sram_mem[111454] = 16'b0000000000000000;
	sram_mem[111455] = 16'b0000000000000000;
	sram_mem[111456] = 16'b0000000000000000;
	sram_mem[111457] = 16'b0000000000000000;
	sram_mem[111458] = 16'b0000000000000000;
	sram_mem[111459] = 16'b0000000000000000;
	sram_mem[111460] = 16'b0000000000000000;
	sram_mem[111461] = 16'b0000000000000000;
	sram_mem[111462] = 16'b0000000000000000;
	sram_mem[111463] = 16'b0000000000000000;
	sram_mem[111464] = 16'b0000000000000000;
	sram_mem[111465] = 16'b0000000000000000;
	sram_mem[111466] = 16'b0000000000000000;
	sram_mem[111467] = 16'b0000000000000000;
	sram_mem[111468] = 16'b0000000000000000;
	sram_mem[111469] = 16'b0000000000000000;
	sram_mem[111470] = 16'b0000000000000000;
	sram_mem[111471] = 16'b0000000000000000;
	sram_mem[111472] = 16'b0000000000000000;
	sram_mem[111473] = 16'b0000000000000000;
	sram_mem[111474] = 16'b0000000000000000;
	sram_mem[111475] = 16'b0000000000000000;
	sram_mem[111476] = 16'b0000000000000000;
	sram_mem[111477] = 16'b0000000000000000;
	sram_mem[111478] = 16'b0000000000000000;
	sram_mem[111479] = 16'b0000000000000000;
	sram_mem[111480] = 16'b0000000000000000;
	sram_mem[111481] = 16'b0000000000000000;
	sram_mem[111482] = 16'b0000000000000000;
	sram_mem[111483] = 16'b0000000000000000;
	sram_mem[111484] = 16'b0000000000000000;
	sram_mem[111485] = 16'b0000000000000000;
	sram_mem[111486] = 16'b0000000000000000;
	sram_mem[111487] = 16'b0000000000000000;
	sram_mem[111488] = 16'b0000000000000000;
	sram_mem[111489] = 16'b0000000000000000;
	sram_mem[111490] = 16'b0000000000000000;
	sram_mem[111491] = 16'b0000000000000000;
	sram_mem[111492] = 16'b0000000000000000;
	sram_mem[111493] = 16'b0000000000000000;
	sram_mem[111494] = 16'b0000000000000000;
	sram_mem[111495] = 16'b0000000000000000;
	sram_mem[111496] = 16'b0000000000000000;
	sram_mem[111497] = 16'b0000000000000000;
	sram_mem[111498] = 16'b0000000000000000;
	sram_mem[111499] = 16'b0000000000000000;
	sram_mem[111500] = 16'b0000000000000000;
	sram_mem[111501] = 16'b0000000000000000;
	sram_mem[111502] = 16'b0000000000000000;
	sram_mem[111503] = 16'b0000000000000000;
	sram_mem[111504] = 16'b0000000000000000;
	sram_mem[111505] = 16'b0000000000000000;
	sram_mem[111506] = 16'b0000000000000000;
	sram_mem[111507] = 16'b0000000000000000;
	sram_mem[111508] = 16'b0000000000000000;
	sram_mem[111509] = 16'b0000000000000000;
	sram_mem[111510] = 16'b0000000000000000;
	sram_mem[111511] = 16'b0000000000000000;
	sram_mem[111512] = 16'b0000000000000000;
	sram_mem[111513] = 16'b0000000000000000;
	sram_mem[111514] = 16'b0000000000000000;
	sram_mem[111515] = 16'b0000000000000000;
	sram_mem[111516] = 16'b0000000000000000;
	sram_mem[111517] = 16'b0000000000000000;
	sram_mem[111518] = 16'b0000000000000000;
	sram_mem[111519] = 16'b0000000000000000;
	sram_mem[111520] = 16'b0000000000000000;
	sram_mem[111521] = 16'b0000000000000000;
	sram_mem[111522] = 16'b0000000000000000;
	sram_mem[111523] = 16'b0000000000000000;
	sram_mem[111524] = 16'b0000000000000000;
	sram_mem[111525] = 16'b0000000000000000;
	sram_mem[111526] = 16'b0000000000000000;
	sram_mem[111527] = 16'b0000000000000000;
	sram_mem[111528] = 16'b0000000000000000;
	sram_mem[111529] = 16'b0000000000000000;
	sram_mem[111530] = 16'b0000000000000000;
	sram_mem[111531] = 16'b0000000000000000;
	sram_mem[111532] = 16'b0000000000000000;
	sram_mem[111533] = 16'b0000000000000000;
	sram_mem[111534] = 16'b0000000000000000;
	sram_mem[111535] = 16'b0000000000000000;
	sram_mem[111536] = 16'b0000000000000000;
	sram_mem[111537] = 16'b0000000000000000;
	sram_mem[111538] = 16'b0000000000000000;
	sram_mem[111539] = 16'b0000000000000000;
	sram_mem[111540] = 16'b0000000000000000;
	sram_mem[111541] = 16'b0000000000000000;
	sram_mem[111542] = 16'b0000000000000000;
	sram_mem[111543] = 16'b0000000000000000;
	sram_mem[111544] = 16'b0000000000000000;
	sram_mem[111545] = 16'b0000000000000000;
	sram_mem[111546] = 16'b0000000000000000;
	sram_mem[111547] = 16'b0000000000000000;
	sram_mem[111548] = 16'b0000000000000000;
	sram_mem[111549] = 16'b0000000000000000;
	sram_mem[111550] = 16'b0000000000000000;
	sram_mem[111551] = 16'b0000000000000000;
	sram_mem[111552] = 16'b0000000000000000;
	sram_mem[111553] = 16'b0000000000000000;
	sram_mem[111554] = 16'b0000000000000000;
	sram_mem[111555] = 16'b0000000000000000;
	sram_mem[111556] = 16'b0000000000000000;
	sram_mem[111557] = 16'b0000000000000000;
	sram_mem[111558] = 16'b0000000000000000;
	sram_mem[111559] = 16'b0000000000000000;
	sram_mem[111560] = 16'b0000000000000000;
	sram_mem[111561] = 16'b0000000000000000;
	sram_mem[111562] = 16'b0000000000000000;
	sram_mem[111563] = 16'b0000000000000000;
	sram_mem[111564] = 16'b0000000000000000;
	sram_mem[111565] = 16'b0000000000000000;
	sram_mem[111566] = 16'b0000000000000000;
	sram_mem[111567] = 16'b0000000000000000;
	sram_mem[111568] = 16'b0000000000000000;
	sram_mem[111569] = 16'b0000000000000000;
	sram_mem[111570] = 16'b0000000000000000;
	sram_mem[111571] = 16'b0000000000000000;
	sram_mem[111572] = 16'b0000000000000000;
	sram_mem[111573] = 16'b0000000000000000;
	sram_mem[111574] = 16'b0000000000000000;
	sram_mem[111575] = 16'b0000000000000000;
	sram_mem[111576] = 16'b0000000000000000;
	sram_mem[111577] = 16'b0000000000000000;
	sram_mem[111578] = 16'b0000000000000000;
	sram_mem[111579] = 16'b0000000000000000;
	sram_mem[111580] = 16'b0000000000000000;
	sram_mem[111581] = 16'b0000000000000000;
	sram_mem[111582] = 16'b0000000000000000;
	sram_mem[111583] = 16'b0000000000000000;
	sram_mem[111584] = 16'b0000000000000000;
	sram_mem[111585] = 16'b0000000000000000;
	sram_mem[111586] = 16'b0000000000000000;
	sram_mem[111587] = 16'b0000000000000000;
	sram_mem[111588] = 16'b0000000000000000;
	sram_mem[111589] = 16'b0000000000000000;
	sram_mem[111590] = 16'b0000000000000000;
	sram_mem[111591] = 16'b0000000000000000;
	sram_mem[111592] = 16'b0000000000000000;
	sram_mem[111593] = 16'b0000000000000000;
	sram_mem[111594] = 16'b0000000000000000;
	sram_mem[111595] = 16'b0000000000000000;
	sram_mem[111596] = 16'b0000000000000000;
	sram_mem[111597] = 16'b0000000000000000;
	sram_mem[111598] = 16'b0000000000000000;
	sram_mem[111599] = 16'b0000000000000000;
	sram_mem[111600] = 16'b0000000000000000;
	sram_mem[111601] = 16'b0000000000000000;
	sram_mem[111602] = 16'b0000000000000000;
	sram_mem[111603] = 16'b0000000000000000;
	sram_mem[111604] = 16'b0000000000000000;
	sram_mem[111605] = 16'b0000000000000000;
	sram_mem[111606] = 16'b0000000000000000;
	sram_mem[111607] = 16'b0000000000000000;
	sram_mem[111608] = 16'b0000000000000000;
	sram_mem[111609] = 16'b0000000000000000;
	sram_mem[111610] = 16'b0000000000000000;
	sram_mem[111611] = 16'b0000000000000000;
	sram_mem[111612] = 16'b0000000000000000;
	sram_mem[111613] = 16'b0000000000000000;
	sram_mem[111614] = 16'b0000000000000000;
	sram_mem[111615] = 16'b0000000000000000;
	sram_mem[111616] = 16'b0000000000000000;
	sram_mem[111617] = 16'b0000000000000000;
	sram_mem[111618] = 16'b0000000000000000;
	sram_mem[111619] = 16'b0000000000000000;
	sram_mem[111620] = 16'b0000000000000000;
	sram_mem[111621] = 16'b0000000000000000;
	sram_mem[111622] = 16'b0000000000000000;
	sram_mem[111623] = 16'b0000000000000000;
	sram_mem[111624] = 16'b0000000000000000;
	sram_mem[111625] = 16'b0000000000000000;
	sram_mem[111626] = 16'b0000000000000000;
	sram_mem[111627] = 16'b0000000000000000;
	sram_mem[111628] = 16'b0000000000000000;
	sram_mem[111629] = 16'b0000000000000000;
	sram_mem[111630] = 16'b0000000000000000;
	sram_mem[111631] = 16'b0000000000000000;
	sram_mem[111632] = 16'b0000000000000000;
	sram_mem[111633] = 16'b0000000000000000;
	sram_mem[111634] = 16'b0000000000000000;
	sram_mem[111635] = 16'b0000000000000000;
	sram_mem[111636] = 16'b0000000000000000;
	sram_mem[111637] = 16'b0000000000000000;
	sram_mem[111638] = 16'b0000000000000000;
	sram_mem[111639] = 16'b0000000000000000;
	sram_mem[111640] = 16'b0000000000000000;
	sram_mem[111641] = 16'b0000000000000000;
	sram_mem[111642] = 16'b0000000000000000;
	sram_mem[111643] = 16'b0000000000000000;
	sram_mem[111644] = 16'b0000000000000000;
	sram_mem[111645] = 16'b0000000000000000;
	sram_mem[111646] = 16'b0000000000000000;
	sram_mem[111647] = 16'b0000000000000000;
	sram_mem[111648] = 16'b0000000000000000;
	sram_mem[111649] = 16'b0000000000000000;
	sram_mem[111650] = 16'b0000000000000000;
	sram_mem[111651] = 16'b0000000000000000;
	sram_mem[111652] = 16'b0000000000000000;
	sram_mem[111653] = 16'b0000000000000000;
	sram_mem[111654] = 16'b0000000000000000;
	sram_mem[111655] = 16'b0000000000000000;
	sram_mem[111656] = 16'b0000000000000000;
	sram_mem[111657] = 16'b0000000000000000;
	sram_mem[111658] = 16'b0000000000000000;
	sram_mem[111659] = 16'b0000000000000000;
	sram_mem[111660] = 16'b0000000000000000;
	sram_mem[111661] = 16'b0000000000000000;
	sram_mem[111662] = 16'b0000000000000000;
	sram_mem[111663] = 16'b0000000000000000;
	sram_mem[111664] = 16'b0000000000000000;
	sram_mem[111665] = 16'b0000000000000000;
	sram_mem[111666] = 16'b0000000000000000;
	sram_mem[111667] = 16'b0000000000000000;
	sram_mem[111668] = 16'b0000000000000000;
	sram_mem[111669] = 16'b0000000000000000;
	sram_mem[111670] = 16'b0000000000000000;
	sram_mem[111671] = 16'b0000000000000000;
	sram_mem[111672] = 16'b0000000000000000;
	sram_mem[111673] = 16'b0000000000000000;
	sram_mem[111674] = 16'b0000000000000000;
	sram_mem[111675] = 16'b0000000000000000;
	sram_mem[111676] = 16'b0000000000000000;
	sram_mem[111677] = 16'b0000000000000000;
	sram_mem[111678] = 16'b0000000000000000;
	sram_mem[111679] = 16'b0000000000000000;
	sram_mem[111680] = 16'b0000000000000000;
	sram_mem[111681] = 16'b0000000000000000;
	sram_mem[111682] = 16'b0000000000000000;
	sram_mem[111683] = 16'b0000000000000000;
	sram_mem[111684] = 16'b0000000000000000;
	sram_mem[111685] = 16'b0000000000000000;
	sram_mem[111686] = 16'b0000000000000000;
	sram_mem[111687] = 16'b0000000000000000;
	sram_mem[111688] = 16'b0000000000000000;
	sram_mem[111689] = 16'b0000000000000000;
	sram_mem[111690] = 16'b0000000000000000;
	sram_mem[111691] = 16'b0000000000000000;
	sram_mem[111692] = 16'b0000000000000000;
	sram_mem[111693] = 16'b0000000000000000;
	sram_mem[111694] = 16'b0000000000000000;
	sram_mem[111695] = 16'b0000000000000000;
	sram_mem[111696] = 16'b0000000000000000;
	sram_mem[111697] = 16'b0000000000000000;
	sram_mem[111698] = 16'b0000000000000000;
	sram_mem[111699] = 16'b0000000000000000;
	sram_mem[111700] = 16'b0000000000000000;
	sram_mem[111701] = 16'b0000000000000000;
	sram_mem[111702] = 16'b0000000000000000;
	sram_mem[111703] = 16'b0000000000000000;
	sram_mem[111704] = 16'b0000000000000000;
	sram_mem[111705] = 16'b0000000000000000;
	sram_mem[111706] = 16'b0000000000000000;
	sram_mem[111707] = 16'b0000000000000000;
	sram_mem[111708] = 16'b0000000000000000;
	sram_mem[111709] = 16'b0000000000000000;
	sram_mem[111710] = 16'b0000000000000000;
	sram_mem[111711] = 16'b0000000000000000;
	sram_mem[111712] = 16'b0000000000000000;
	sram_mem[111713] = 16'b0000000000000000;
	sram_mem[111714] = 16'b0000000000000000;
	sram_mem[111715] = 16'b0000000000000000;
	sram_mem[111716] = 16'b0000000000000000;
	sram_mem[111717] = 16'b0000000000000000;
	sram_mem[111718] = 16'b0000000000000000;
	sram_mem[111719] = 16'b0000000000000000;
	sram_mem[111720] = 16'b0000000000000000;
	sram_mem[111721] = 16'b0000000000000000;
	sram_mem[111722] = 16'b0000000000000000;
	sram_mem[111723] = 16'b0000000000000000;
	sram_mem[111724] = 16'b0000000000000000;
	sram_mem[111725] = 16'b0000000000000000;
	sram_mem[111726] = 16'b0000000000000000;
	sram_mem[111727] = 16'b0000000000000000;
	sram_mem[111728] = 16'b0000000000000000;
	sram_mem[111729] = 16'b0000000000000000;
	sram_mem[111730] = 16'b0000000000000000;
	sram_mem[111731] = 16'b0000000000000000;
	sram_mem[111732] = 16'b0000000000000000;
	sram_mem[111733] = 16'b0000000000000000;
	sram_mem[111734] = 16'b0000000000000000;
	sram_mem[111735] = 16'b0000000000000000;
	sram_mem[111736] = 16'b0000000000000000;
	sram_mem[111737] = 16'b0000000000000000;
	sram_mem[111738] = 16'b0000000000000000;
	sram_mem[111739] = 16'b0000000000000000;
	sram_mem[111740] = 16'b0000000000000000;
	sram_mem[111741] = 16'b0000000000000000;
	sram_mem[111742] = 16'b0000000000000000;
	sram_mem[111743] = 16'b0000000000000000;
	sram_mem[111744] = 16'b0000000000000000;
	sram_mem[111745] = 16'b0000000000000000;
	sram_mem[111746] = 16'b0000000000000000;
	sram_mem[111747] = 16'b0000000000000000;
	sram_mem[111748] = 16'b0000000000000000;
	sram_mem[111749] = 16'b0000000000000000;
	sram_mem[111750] = 16'b0000000000000000;
	sram_mem[111751] = 16'b0000000000000000;
	sram_mem[111752] = 16'b0000000000000000;
	sram_mem[111753] = 16'b0000000000000000;
	sram_mem[111754] = 16'b0000000000000000;
	sram_mem[111755] = 16'b0000000000000000;
	sram_mem[111756] = 16'b0000000000000000;
	sram_mem[111757] = 16'b0000000000000000;
	sram_mem[111758] = 16'b0000000000000000;
	sram_mem[111759] = 16'b0000000000000000;
	sram_mem[111760] = 16'b0000000000000000;
	sram_mem[111761] = 16'b0000000000000000;
	sram_mem[111762] = 16'b0000000000000000;
	sram_mem[111763] = 16'b0000000000000000;
	sram_mem[111764] = 16'b0000000000000000;
	sram_mem[111765] = 16'b0000000000000000;
	sram_mem[111766] = 16'b0000000000000000;
	sram_mem[111767] = 16'b0000000000000000;
	sram_mem[111768] = 16'b0000000000000000;
	sram_mem[111769] = 16'b0000000000000000;
	sram_mem[111770] = 16'b0000000000000000;
	sram_mem[111771] = 16'b0000000000000000;
	sram_mem[111772] = 16'b0000000000000000;
	sram_mem[111773] = 16'b0000000000000000;
	sram_mem[111774] = 16'b0000000000000000;
	sram_mem[111775] = 16'b0000000000000000;
	sram_mem[111776] = 16'b0000000000000000;
	sram_mem[111777] = 16'b0000000000000000;
	sram_mem[111778] = 16'b0000000000000000;
	sram_mem[111779] = 16'b0000000000000000;
	sram_mem[111780] = 16'b0000000000000000;
	sram_mem[111781] = 16'b0000000000000000;
	sram_mem[111782] = 16'b0000000000000000;
	sram_mem[111783] = 16'b0000000000000000;
	sram_mem[111784] = 16'b0000000000000000;
	sram_mem[111785] = 16'b0000000000000000;
	sram_mem[111786] = 16'b0000000000000000;
	sram_mem[111787] = 16'b0000000000000000;
	sram_mem[111788] = 16'b0000000000000000;
	sram_mem[111789] = 16'b0000000000000000;
	sram_mem[111790] = 16'b0000000000000000;
	sram_mem[111791] = 16'b0000000000000000;
	sram_mem[111792] = 16'b0000000000000000;
	sram_mem[111793] = 16'b0000000000000000;
	sram_mem[111794] = 16'b0000000000000000;
	sram_mem[111795] = 16'b0000000000000000;
	sram_mem[111796] = 16'b0000000000000000;
	sram_mem[111797] = 16'b0000000000000000;
	sram_mem[111798] = 16'b0000000000000000;
	sram_mem[111799] = 16'b0000000000000000;
	sram_mem[111800] = 16'b0000000000000000;
	sram_mem[111801] = 16'b0000000000000000;
	sram_mem[111802] = 16'b0000000000000000;
	sram_mem[111803] = 16'b0000000000000000;
	sram_mem[111804] = 16'b0000000000000000;
	sram_mem[111805] = 16'b0000000000000000;
	sram_mem[111806] = 16'b0000000000000000;
	sram_mem[111807] = 16'b0000000000000000;
	sram_mem[111808] = 16'b0000000000000000;
	sram_mem[111809] = 16'b0000000000000000;
	sram_mem[111810] = 16'b0000000000000000;
	sram_mem[111811] = 16'b0000000000000000;
	sram_mem[111812] = 16'b0000000000000000;
	sram_mem[111813] = 16'b0000000000000000;
	sram_mem[111814] = 16'b0000000000000000;
	sram_mem[111815] = 16'b0000000000000000;
	sram_mem[111816] = 16'b0000000000000000;
	sram_mem[111817] = 16'b0000000000000000;
	sram_mem[111818] = 16'b0000000000000000;
	sram_mem[111819] = 16'b0000000000000000;
	sram_mem[111820] = 16'b0000000000000000;
	sram_mem[111821] = 16'b0000000000000000;
	sram_mem[111822] = 16'b0000000000000000;
	sram_mem[111823] = 16'b0000000000000000;
	sram_mem[111824] = 16'b0000000000000000;
	sram_mem[111825] = 16'b0000000000000000;
	sram_mem[111826] = 16'b0000000000000000;
	sram_mem[111827] = 16'b0000000000000000;
	sram_mem[111828] = 16'b0000000000000000;
	sram_mem[111829] = 16'b0000000000000000;
	sram_mem[111830] = 16'b0000000000000000;
	sram_mem[111831] = 16'b0000000000000000;
	sram_mem[111832] = 16'b0000000000000000;
	sram_mem[111833] = 16'b0000000000000000;
	sram_mem[111834] = 16'b0000000000000000;
	sram_mem[111835] = 16'b0000000000000000;
	sram_mem[111836] = 16'b0000000000000000;
	sram_mem[111837] = 16'b0000000000000000;
	sram_mem[111838] = 16'b0000000000000000;
	sram_mem[111839] = 16'b0000000000000000;
	sram_mem[111840] = 16'b0000000000000000;
	sram_mem[111841] = 16'b0000000000000000;
	sram_mem[111842] = 16'b0000000000000000;
	sram_mem[111843] = 16'b0000000000000000;
	sram_mem[111844] = 16'b0000000000000000;
	sram_mem[111845] = 16'b0000000000000000;
	sram_mem[111846] = 16'b0000000000000000;
	sram_mem[111847] = 16'b0000000000000000;
	sram_mem[111848] = 16'b0000000000000000;
	sram_mem[111849] = 16'b0000000000000000;
	sram_mem[111850] = 16'b0000000000000000;
	sram_mem[111851] = 16'b0000000000000000;
	sram_mem[111852] = 16'b0000000000000000;
	sram_mem[111853] = 16'b0000000000000000;
	sram_mem[111854] = 16'b0000000000000000;
	sram_mem[111855] = 16'b0000000000000000;
	sram_mem[111856] = 16'b0000000000000000;
	sram_mem[111857] = 16'b0000000000000000;
	sram_mem[111858] = 16'b0000000000000000;
	sram_mem[111859] = 16'b0000000000000000;
	sram_mem[111860] = 16'b0000000000000000;
	sram_mem[111861] = 16'b0000000000000000;
	sram_mem[111862] = 16'b0000000000000000;
	sram_mem[111863] = 16'b0000000000000000;
	sram_mem[111864] = 16'b0000000000000000;
	sram_mem[111865] = 16'b0000000000000000;
	sram_mem[111866] = 16'b0000000000000000;
	sram_mem[111867] = 16'b0000000000000000;
	sram_mem[111868] = 16'b0000000000000000;
	sram_mem[111869] = 16'b0000000000000000;
	sram_mem[111870] = 16'b0000000000000000;
	sram_mem[111871] = 16'b0000000000000000;
	sram_mem[111872] = 16'b0000000000000000;
	sram_mem[111873] = 16'b0000000000000000;
	sram_mem[111874] = 16'b0000000000000000;
	sram_mem[111875] = 16'b0000000000000000;
	sram_mem[111876] = 16'b0000000000000000;
	sram_mem[111877] = 16'b0000000000000000;
	sram_mem[111878] = 16'b0000000000000000;
	sram_mem[111879] = 16'b0000000000000000;
	sram_mem[111880] = 16'b0000000000000000;
	sram_mem[111881] = 16'b0000000000000000;
	sram_mem[111882] = 16'b0000000000000000;
	sram_mem[111883] = 16'b0000000000000000;
	sram_mem[111884] = 16'b0000000000000000;
	sram_mem[111885] = 16'b0000000000000000;
	sram_mem[111886] = 16'b0000000000000000;
	sram_mem[111887] = 16'b0000000000000000;
	sram_mem[111888] = 16'b0000000000000000;
	sram_mem[111889] = 16'b0000000000000000;
	sram_mem[111890] = 16'b0000000000000000;
	sram_mem[111891] = 16'b0000000000000000;
	sram_mem[111892] = 16'b0000000000000000;
	sram_mem[111893] = 16'b0000000000000000;
	sram_mem[111894] = 16'b0000000000000000;
	sram_mem[111895] = 16'b0000000000000000;
	sram_mem[111896] = 16'b0000000000000000;
	sram_mem[111897] = 16'b0000000000000000;
	sram_mem[111898] = 16'b0000000000000000;
	sram_mem[111899] = 16'b0000000000000000;
	sram_mem[111900] = 16'b0000000000000000;
	sram_mem[111901] = 16'b0000000000000000;
	sram_mem[111902] = 16'b0000000000000000;
	sram_mem[111903] = 16'b0000000000000000;
	sram_mem[111904] = 16'b0000000000000000;
	sram_mem[111905] = 16'b0000000000000000;
	sram_mem[111906] = 16'b0000000000000000;
	sram_mem[111907] = 16'b0000000000000000;
	sram_mem[111908] = 16'b0000000000000000;
	sram_mem[111909] = 16'b0000000000000000;
	sram_mem[111910] = 16'b0000000000000000;
	sram_mem[111911] = 16'b0000000000000000;
	sram_mem[111912] = 16'b0000000000000000;
	sram_mem[111913] = 16'b0000000000000000;
	sram_mem[111914] = 16'b0000000000000000;
	sram_mem[111915] = 16'b0000000000000000;
	sram_mem[111916] = 16'b0000000000000000;
	sram_mem[111917] = 16'b0000000000000000;
	sram_mem[111918] = 16'b0000000000000000;
	sram_mem[111919] = 16'b0000000000000000;
	sram_mem[111920] = 16'b0000000000000000;
	sram_mem[111921] = 16'b0000000000000000;
	sram_mem[111922] = 16'b0000000000000000;
	sram_mem[111923] = 16'b0000000000000000;
	sram_mem[111924] = 16'b0000000000000000;
	sram_mem[111925] = 16'b0000000000000000;
	sram_mem[111926] = 16'b0000000000000000;
	sram_mem[111927] = 16'b0000000000000000;
	sram_mem[111928] = 16'b0000000000000000;
	sram_mem[111929] = 16'b0000000000000000;
	sram_mem[111930] = 16'b0000000000000000;
	sram_mem[111931] = 16'b0000000000000000;
	sram_mem[111932] = 16'b0000000000000000;
	sram_mem[111933] = 16'b0000000000000000;
	sram_mem[111934] = 16'b0000000000000000;
	sram_mem[111935] = 16'b0000000000000000;
	sram_mem[111936] = 16'b0000000000000000;
	sram_mem[111937] = 16'b0000000000000000;
	sram_mem[111938] = 16'b0000000000000000;
	sram_mem[111939] = 16'b0000000000000000;
	sram_mem[111940] = 16'b0000000000000000;
	sram_mem[111941] = 16'b0000000000000000;
	sram_mem[111942] = 16'b0000000000000000;
	sram_mem[111943] = 16'b0000000000000000;
	sram_mem[111944] = 16'b0000000000000000;
	sram_mem[111945] = 16'b0000000000000000;
	sram_mem[111946] = 16'b0000000000000000;
	sram_mem[111947] = 16'b0000000000000000;
	sram_mem[111948] = 16'b0000000000000000;
	sram_mem[111949] = 16'b0000000000000000;
	sram_mem[111950] = 16'b0000000000000000;
	sram_mem[111951] = 16'b0000000000000000;
	sram_mem[111952] = 16'b0000000000000000;
	sram_mem[111953] = 16'b0000000000000000;
	sram_mem[111954] = 16'b0000000000000000;
	sram_mem[111955] = 16'b0000000000000000;
	sram_mem[111956] = 16'b0000000000000000;
	sram_mem[111957] = 16'b0000000000000000;
	sram_mem[111958] = 16'b0000000000000000;
	sram_mem[111959] = 16'b0000000000000000;
	sram_mem[111960] = 16'b0000000000000000;
	sram_mem[111961] = 16'b0000000000000000;
	sram_mem[111962] = 16'b0000000000000000;
	sram_mem[111963] = 16'b0000000000000000;
	sram_mem[111964] = 16'b0000000000000000;
	sram_mem[111965] = 16'b0000000000000000;
	sram_mem[111966] = 16'b0000000000000000;
	sram_mem[111967] = 16'b0000000000000000;
	sram_mem[111968] = 16'b0000000000000000;
	sram_mem[111969] = 16'b0000000000000000;
	sram_mem[111970] = 16'b0000000000000000;
	sram_mem[111971] = 16'b0000000000000000;
	sram_mem[111972] = 16'b0000000000000000;
	sram_mem[111973] = 16'b0000000000000000;
	sram_mem[111974] = 16'b0000000000000000;
	sram_mem[111975] = 16'b0000000000000000;
	sram_mem[111976] = 16'b0000000000000000;
	sram_mem[111977] = 16'b0000000000000000;
	sram_mem[111978] = 16'b0000000000000000;
	sram_mem[111979] = 16'b0000000000000000;
	sram_mem[111980] = 16'b0000000000000000;
	sram_mem[111981] = 16'b0000000000000000;
	sram_mem[111982] = 16'b0000000000000000;
	sram_mem[111983] = 16'b0000000000000000;
	sram_mem[111984] = 16'b0000000000000000;
	sram_mem[111985] = 16'b0000000000000000;
	sram_mem[111986] = 16'b0000000000000000;
	sram_mem[111987] = 16'b0000000000000000;
	sram_mem[111988] = 16'b0000000000000000;
	sram_mem[111989] = 16'b0000000000000000;
	sram_mem[111990] = 16'b0000000000000000;
	sram_mem[111991] = 16'b0000000000000000;
	sram_mem[111992] = 16'b0000000000000000;
	sram_mem[111993] = 16'b0000000000000000;
	sram_mem[111994] = 16'b0000000000000000;
	sram_mem[111995] = 16'b0000000000000000;
	sram_mem[111996] = 16'b0000000000000000;
	sram_mem[111997] = 16'b0000000000000000;
	sram_mem[111998] = 16'b0000000000000000;
	sram_mem[111999] = 16'b0000000000000000;
	sram_mem[112000] = 16'b0000000000000000;
	sram_mem[112001] = 16'b0000000000000000;
	sram_mem[112002] = 16'b0000000000000000;
	sram_mem[112003] = 16'b0000000000000000;
	sram_mem[112004] = 16'b0000000000000000;
	sram_mem[112005] = 16'b0000000000000000;
	sram_mem[112006] = 16'b0000000000000000;
	sram_mem[112007] = 16'b0000000000000000;
	sram_mem[112008] = 16'b0000000000000000;
	sram_mem[112009] = 16'b0000000000000000;
	sram_mem[112010] = 16'b0000000000000000;
	sram_mem[112011] = 16'b0000000000000000;
	sram_mem[112012] = 16'b0000000000000000;
	sram_mem[112013] = 16'b0000000000000000;
	sram_mem[112014] = 16'b0000000000000000;
	sram_mem[112015] = 16'b0000000000000000;
	sram_mem[112016] = 16'b0000000000000000;
	sram_mem[112017] = 16'b0000000000000000;
	sram_mem[112018] = 16'b0000000000000000;
	sram_mem[112019] = 16'b0000000000000000;
	sram_mem[112020] = 16'b0000000000000000;
	sram_mem[112021] = 16'b0000000000000000;
	sram_mem[112022] = 16'b0000000000000000;
	sram_mem[112023] = 16'b0000000000000000;
	sram_mem[112024] = 16'b0000000000000000;
	sram_mem[112025] = 16'b0000000000000000;
	sram_mem[112026] = 16'b0000000000000000;
	sram_mem[112027] = 16'b0000000000000000;
	sram_mem[112028] = 16'b0000000000000000;
	sram_mem[112029] = 16'b0000000000000000;
	sram_mem[112030] = 16'b0000000000000000;
	sram_mem[112031] = 16'b0000000000000000;
	sram_mem[112032] = 16'b0000000000000000;
	sram_mem[112033] = 16'b0000000000000000;
	sram_mem[112034] = 16'b0000000000000000;
	sram_mem[112035] = 16'b0000000000000000;
	sram_mem[112036] = 16'b0000000000000000;
	sram_mem[112037] = 16'b0000000000000000;
	sram_mem[112038] = 16'b0000000000000000;
	sram_mem[112039] = 16'b0000000000000000;
	sram_mem[112040] = 16'b0000000000000000;
	sram_mem[112041] = 16'b0000000000000000;
	sram_mem[112042] = 16'b0000000000000000;
	sram_mem[112043] = 16'b0000000000000000;
	sram_mem[112044] = 16'b0000000000000000;
	sram_mem[112045] = 16'b0000000000000000;
	sram_mem[112046] = 16'b0000000000000000;
	sram_mem[112047] = 16'b0000000000000000;
	sram_mem[112048] = 16'b0000000000000000;
	sram_mem[112049] = 16'b0000000000000000;
	sram_mem[112050] = 16'b0000000000000000;
	sram_mem[112051] = 16'b0000000000000000;
	sram_mem[112052] = 16'b0000000000000000;
	sram_mem[112053] = 16'b0000000000000000;
	sram_mem[112054] = 16'b0000000000000000;
	sram_mem[112055] = 16'b0000000000000000;
	sram_mem[112056] = 16'b0000000000000000;
	sram_mem[112057] = 16'b0000000000000000;
	sram_mem[112058] = 16'b0000000000000000;
	sram_mem[112059] = 16'b0000000000000000;
	sram_mem[112060] = 16'b0000000000000000;
	sram_mem[112061] = 16'b0000000000000000;
	sram_mem[112062] = 16'b0000000000000000;
	sram_mem[112063] = 16'b0000000000000000;
	sram_mem[112064] = 16'b0000000000000000;
	sram_mem[112065] = 16'b0000000000000000;
	sram_mem[112066] = 16'b0000000000000000;
	sram_mem[112067] = 16'b0000000000000000;
	sram_mem[112068] = 16'b0000000000000000;
	sram_mem[112069] = 16'b0000000000000000;
	sram_mem[112070] = 16'b0000000000000000;
	sram_mem[112071] = 16'b0000000000000000;
	sram_mem[112072] = 16'b0000000000000000;
	sram_mem[112073] = 16'b0000000000000000;
	sram_mem[112074] = 16'b0000000000000000;
	sram_mem[112075] = 16'b0000000000000000;
	sram_mem[112076] = 16'b0000000000000000;
	sram_mem[112077] = 16'b0000000000000000;
	sram_mem[112078] = 16'b0000000000000000;
	sram_mem[112079] = 16'b0000000000000000;
	sram_mem[112080] = 16'b0000000000000000;
	sram_mem[112081] = 16'b0000000000000000;
	sram_mem[112082] = 16'b0000000000000000;
	sram_mem[112083] = 16'b0000000000000000;
	sram_mem[112084] = 16'b0000000000000000;
	sram_mem[112085] = 16'b0000000000000000;
	sram_mem[112086] = 16'b0000000000000000;
	sram_mem[112087] = 16'b0000000000000000;
	sram_mem[112088] = 16'b0000000000000000;
	sram_mem[112089] = 16'b0000000000000000;
	sram_mem[112090] = 16'b0000000000000000;
	sram_mem[112091] = 16'b0000000000000000;
	sram_mem[112092] = 16'b0000000000000000;
	sram_mem[112093] = 16'b0000000000000000;
	sram_mem[112094] = 16'b0000000000000000;
	sram_mem[112095] = 16'b0000000000000000;
	sram_mem[112096] = 16'b0000000000000000;
	sram_mem[112097] = 16'b0000000000000000;
	sram_mem[112098] = 16'b0000000000000000;
	sram_mem[112099] = 16'b0000000000000000;
	sram_mem[112100] = 16'b0000000000000000;
	sram_mem[112101] = 16'b0000000000000000;
	sram_mem[112102] = 16'b0000000000000000;
	sram_mem[112103] = 16'b0000000000000000;
	sram_mem[112104] = 16'b0000000000000000;
	sram_mem[112105] = 16'b0000000000000000;
	sram_mem[112106] = 16'b0000000000000000;
	sram_mem[112107] = 16'b0000000000000000;
	sram_mem[112108] = 16'b0000000000000000;
	sram_mem[112109] = 16'b0000000000000000;
	sram_mem[112110] = 16'b0000000000000000;
	sram_mem[112111] = 16'b0000000000000000;
	sram_mem[112112] = 16'b0000000000000000;
	sram_mem[112113] = 16'b0000000000000000;
	sram_mem[112114] = 16'b0000000000000000;
	sram_mem[112115] = 16'b0000000000000000;
	sram_mem[112116] = 16'b0000000000000000;
	sram_mem[112117] = 16'b0000000000000000;
	sram_mem[112118] = 16'b0000000000000000;
	sram_mem[112119] = 16'b0000000000000000;
	sram_mem[112120] = 16'b0000000000000000;
	sram_mem[112121] = 16'b0000000000000000;
	sram_mem[112122] = 16'b0000000000000000;
	sram_mem[112123] = 16'b0000000000000000;
	sram_mem[112124] = 16'b0000000000000000;
	sram_mem[112125] = 16'b0000000000000000;
	sram_mem[112126] = 16'b0000000000000000;
	sram_mem[112127] = 16'b0000000000000000;
	sram_mem[112128] = 16'b0000000000000000;
	sram_mem[112129] = 16'b0000000000000000;
	sram_mem[112130] = 16'b0000000000000000;
	sram_mem[112131] = 16'b0000000000000000;
	sram_mem[112132] = 16'b0000000000000000;
	sram_mem[112133] = 16'b0000000000000000;
	sram_mem[112134] = 16'b0000000000000000;
	sram_mem[112135] = 16'b0000000000000000;
	sram_mem[112136] = 16'b0000000000000000;
	sram_mem[112137] = 16'b0000000000000000;
	sram_mem[112138] = 16'b0000000000000000;
	sram_mem[112139] = 16'b0000000000000000;
	sram_mem[112140] = 16'b0000000000000000;
	sram_mem[112141] = 16'b0000000000000000;
	sram_mem[112142] = 16'b0000000000000000;
	sram_mem[112143] = 16'b0000000000000000;
	sram_mem[112144] = 16'b0000000000000000;
	sram_mem[112145] = 16'b0000000000000000;
	sram_mem[112146] = 16'b0000000000000000;
	sram_mem[112147] = 16'b0000000000000000;
	sram_mem[112148] = 16'b0000000000000000;
	sram_mem[112149] = 16'b0000000000000000;
	sram_mem[112150] = 16'b0000000000000000;
	sram_mem[112151] = 16'b0000000000000000;
	sram_mem[112152] = 16'b0000000000000000;
	sram_mem[112153] = 16'b0000000000000000;
	sram_mem[112154] = 16'b0000000000000000;
	sram_mem[112155] = 16'b0000000000000000;
	sram_mem[112156] = 16'b0000000000000000;
	sram_mem[112157] = 16'b0000000000000000;
	sram_mem[112158] = 16'b0000000000000000;
	sram_mem[112159] = 16'b0000000000000000;
	sram_mem[112160] = 16'b0000000000000000;
	sram_mem[112161] = 16'b0000000000000000;
	sram_mem[112162] = 16'b0000000000000000;
	sram_mem[112163] = 16'b0000000000000000;
	sram_mem[112164] = 16'b0000000000000000;
	sram_mem[112165] = 16'b0000000000000000;
	sram_mem[112166] = 16'b0000000000000000;
	sram_mem[112167] = 16'b0000000000000000;
	sram_mem[112168] = 16'b0000000000000000;
	sram_mem[112169] = 16'b0000000000000000;
	sram_mem[112170] = 16'b0000000000000000;
	sram_mem[112171] = 16'b0000000000000000;
	sram_mem[112172] = 16'b0000000000000000;
	sram_mem[112173] = 16'b0000000000000000;
	sram_mem[112174] = 16'b0000000000000000;
	sram_mem[112175] = 16'b0000000000000000;
	sram_mem[112176] = 16'b0000000000000000;
	sram_mem[112177] = 16'b0000000000000000;
	sram_mem[112178] = 16'b0000000000000000;
	sram_mem[112179] = 16'b0000000000000000;
	sram_mem[112180] = 16'b0000000000000000;
	sram_mem[112181] = 16'b0000000000000000;
	sram_mem[112182] = 16'b0000000000000000;
	sram_mem[112183] = 16'b0000000000000000;
	sram_mem[112184] = 16'b0000000000000000;
	sram_mem[112185] = 16'b0000000000000000;
	sram_mem[112186] = 16'b0000000000000000;
	sram_mem[112187] = 16'b0000000000000000;
	sram_mem[112188] = 16'b0000000000000000;
	sram_mem[112189] = 16'b0000000000000000;
	sram_mem[112190] = 16'b0000000000000000;
	sram_mem[112191] = 16'b0000000000000000;
	sram_mem[112192] = 16'b0000000000000000;
	sram_mem[112193] = 16'b0000000000000000;
	sram_mem[112194] = 16'b0000000000000000;
	sram_mem[112195] = 16'b0000000000000000;
	sram_mem[112196] = 16'b0000000000000000;
	sram_mem[112197] = 16'b0000000000000000;
	sram_mem[112198] = 16'b0000000000000000;
	sram_mem[112199] = 16'b0000000000000000;
	sram_mem[112200] = 16'b0000000000000000;
	sram_mem[112201] = 16'b0000000000000000;
	sram_mem[112202] = 16'b0000000000000000;
	sram_mem[112203] = 16'b0000000000000000;
	sram_mem[112204] = 16'b0000000000000000;
	sram_mem[112205] = 16'b0000000000000000;
	sram_mem[112206] = 16'b0000000000000000;
	sram_mem[112207] = 16'b0000000000000000;
	sram_mem[112208] = 16'b0000000000000000;
	sram_mem[112209] = 16'b0000000000000000;
	sram_mem[112210] = 16'b0000000000000000;
	sram_mem[112211] = 16'b0000000000000000;
	sram_mem[112212] = 16'b0000000000000000;
	sram_mem[112213] = 16'b0000000000000000;
	sram_mem[112214] = 16'b0000000000000000;
	sram_mem[112215] = 16'b0000000000000000;
	sram_mem[112216] = 16'b0000000000000000;
	sram_mem[112217] = 16'b0000000000000000;
	sram_mem[112218] = 16'b0000000000000000;
	sram_mem[112219] = 16'b0000000000000000;
	sram_mem[112220] = 16'b0000000000000000;
	sram_mem[112221] = 16'b0000000000000000;
	sram_mem[112222] = 16'b0000000000000000;
	sram_mem[112223] = 16'b0000000000000000;
	sram_mem[112224] = 16'b0000000000000000;
	sram_mem[112225] = 16'b0000000000000000;
	sram_mem[112226] = 16'b0000000000000000;
	sram_mem[112227] = 16'b0000000000000000;
	sram_mem[112228] = 16'b0000000000000000;
	sram_mem[112229] = 16'b0000000000000000;
	sram_mem[112230] = 16'b0000000000000000;
	sram_mem[112231] = 16'b0000000000000000;
	sram_mem[112232] = 16'b0000000000000000;
	sram_mem[112233] = 16'b0000000000000000;
	sram_mem[112234] = 16'b0000000000000000;
	sram_mem[112235] = 16'b0000000000000000;
	sram_mem[112236] = 16'b0000000000000000;
	sram_mem[112237] = 16'b0000000000000000;
	sram_mem[112238] = 16'b0000000000000000;
	sram_mem[112239] = 16'b0000000000000000;
	sram_mem[112240] = 16'b0000000000000000;
	sram_mem[112241] = 16'b0000000000000000;
	sram_mem[112242] = 16'b0000000000000000;
	sram_mem[112243] = 16'b0000000000000000;
	sram_mem[112244] = 16'b0000000000000000;
	sram_mem[112245] = 16'b0000000000000000;
	sram_mem[112246] = 16'b0000000000000000;
	sram_mem[112247] = 16'b0000000000000000;
	sram_mem[112248] = 16'b0000000000000000;
	sram_mem[112249] = 16'b0000000000000000;
	sram_mem[112250] = 16'b0000000000000000;
	sram_mem[112251] = 16'b0000000000000000;
	sram_mem[112252] = 16'b0000000000000000;
	sram_mem[112253] = 16'b0000000000000000;
	sram_mem[112254] = 16'b0000000000000000;
	sram_mem[112255] = 16'b0000000000000000;
	sram_mem[112256] = 16'b0000000000000000;
	sram_mem[112257] = 16'b0000000000000000;
	sram_mem[112258] = 16'b0000000000000000;
	sram_mem[112259] = 16'b0000000000000000;
	sram_mem[112260] = 16'b0000000000000000;
	sram_mem[112261] = 16'b0000000000000000;
	sram_mem[112262] = 16'b0000000000000000;
	sram_mem[112263] = 16'b0000000000000000;
	sram_mem[112264] = 16'b0000000000000000;
	sram_mem[112265] = 16'b0000000000000000;
	sram_mem[112266] = 16'b0000000000000000;
	sram_mem[112267] = 16'b0000000000000000;
	sram_mem[112268] = 16'b0000000000000000;
	sram_mem[112269] = 16'b0000000000000000;
	sram_mem[112270] = 16'b0000000000000000;
	sram_mem[112271] = 16'b0000000000000000;
	sram_mem[112272] = 16'b0000000000000000;
	sram_mem[112273] = 16'b0000000000000000;
	sram_mem[112274] = 16'b0000000000000000;
	sram_mem[112275] = 16'b0000000000000000;
	sram_mem[112276] = 16'b0000000000000000;
	sram_mem[112277] = 16'b0000000000000000;
	sram_mem[112278] = 16'b0000000000000000;
	sram_mem[112279] = 16'b0000000000000000;
	sram_mem[112280] = 16'b0000000000000000;
	sram_mem[112281] = 16'b0000000000000000;
	sram_mem[112282] = 16'b0000000000000000;
	sram_mem[112283] = 16'b0000000000000000;
	sram_mem[112284] = 16'b0000000000000000;
	sram_mem[112285] = 16'b0000000000000000;
	sram_mem[112286] = 16'b0000000000000000;
	sram_mem[112287] = 16'b0000000000000000;
	sram_mem[112288] = 16'b0000000000000000;
	sram_mem[112289] = 16'b0000000000000000;
	sram_mem[112290] = 16'b0000000000000000;
	sram_mem[112291] = 16'b0000000000000000;
	sram_mem[112292] = 16'b0000000000000000;
	sram_mem[112293] = 16'b0000000000000000;
	sram_mem[112294] = 16'b0000000000000000;
	sram_mem[112295] = 16'b0000000000000000;
	sram_mem[112296] = 16'b0000000000000000;
	sram_mem[112297] = 16'b0000000000000000;
	sram_mem[112298] = 16'b0000000000000000;
	sram_mem[112299] = 16'b0000000000000000;
	sram_mem[112300] = 16'b0000000000000000;
	sram_mem[112301] = 16'b0000000000000000;
	sram_mem[112302] = 16'b0000000000000000;
	sram_mem[112303] = 16'b0000000000000000;
	sram_mem[112304] = 16'b0000000000000000;
	sram_mem[112305] = 16'b0000000000000000;
	sram_mem[112306] = 16'b0000000000000000;
	sram_mem[112307] = 16'b0000000000000000;
	sram_mem[112308] = 16'b0000000000000000;
	sram_mem[112309] = 16'b0000000000000000;
	sram_mem[112310] = 16'b0000000000000000;
	sram_mem[112311] = 16'b0000000000000000;
	sram_mem[112312] = 16'b0000000000000000;
	sram_mem[112313] = 16'b0000000000000000;
	sram_mem[112314] = 16'b0000000000000000;
	sram_mem[112315] = 16'b0000000000000000;
	sram_mem[112316] = 16'b0000000000000000;
	sram_mem[112317] = 16'b0000000000000000;
	sram_mem[112318] = 16'b0000000000000000;
	sram_mem[112319] = 16'b0000000000000000;
	sram_mem[112320] = 16'b0000000000000000;
	sram_mem[112321] = 16'b0000000000000000;
	sram_mem[112322] = 16'b0000000000000000;
	sram_mem[112323] = 16'b0000000000000000;
	sram_mem[112324] = 16'b0000000000000000;
	sram_mem[112325] = 16'b0000000000000000;
	sram_mem[112326] = 16'b0000000000000000;
	sram_mem[112327] = 16'b0000000000000000;
	sram_mem[112328] = 16'b0000000000000000;
	sram_mem[112329] = 16'b0000000000000000;
	sram_mem[112330] = 16'b0000000000000000;
	sram_mem[112331] = 16'b0000000000000000;
	sram_mem[112332] = 16'b0000000000000000;
	sram_mem[112333] = 16'b0000000000000000;
	sram_mem[112334] = 16'b0000000000000000;
	sram_mem[112335] = 16'b0000000000000000;
	sram_mem[112336] = 16'b0000000000000000;
	sram_mem[112337] = 16'b0000000000000000;
	sram_mem[112338] = 16'b0000000000000000;
	sram_mem[112339] = 16'b0000000000000000;
	sram_mem[112340] = 16'b0000000000000000;
	sram_mem[112341] = 16'b0000000000000000;
	sram_mem[112342] = 16'b0000000000000000;
	sram_mem[112343] = 16'b0000000000000000;
	sram_mem[112344] = 16'b0000000000000000;
	sram_mem[112345] = 16'b0000000000000000;
	sram_mem[112346] = 16'b0000000000000000;
	sram_mem[112347] = 16'b0000000000000000;
	sram_mem[112348] = 16'b0000000000000000;
	sram_mem[112349] = 16'b0000000000000000;
	sram_mem[112350] = 16'b0000000000000000;
	sram_mem[112351] = 16'b0000000000000000;
	sram_mem[112352] = 16'b0000000000000000;
	sram_mem[112353] = 16'b0000000000000000;
	sram_mem[112354] = 16'b0000000000000000;
	sram_mem[112355] = 16'b0000000000000000;
	sram_mem[112356] = 16'b0000000000000000;
	sram_mem[112357] = 16'b0000000000000000;
	sram_mem[112358] = 16'b0000000000000000;
	sram_mem[112359] = 16'b0000000000000000;
	sram_mem[112360] = 16'b0000000000000000;
	sram_mem[112361] = 16'b0000000000000000;
	sram_mem[112362] = 16'b0000000000000000;
	sram_mem[112363] = 16'b0000000000000000;
	sram_mem[112364] = 16'b0000000000000000;
	sram_mem[112365] = 16'b0000000000000000;
	sram_mem[112366] = 16'b0000000000000000;
	sram_mem[112367] = 16'b0000000000000000;
	sram_mem[112368] = 16'b0000000000000000;
	sram_mem[112369] = 16'b0000000000000000;
	sram_mem[112370] = 16'b0000000000000000;
	sram_mem[112371] = 16'b0000000000000000;
	sram_mem[112372] = 16'b0000000000000000;
	sram_mem[112373] = 16'b0000000000000000;
	sram_mem[112374] = 16'b0000000000000000;
	sram_mem[112375] = 16'b0000000000000000;
	sram_mem[112376] = 16'b0000000000000000;
	sram_mem[112377] = 16'b0000000000000000;
	sram_mem[112378] = 16'b0000000000000000;
	sram_mem[112379] = 16'b0000000000000000;
	sram_mem[112380] = 16'b0000000000000000;
	sram_mem[112381] = 16'b0000000000000000;
	sram_mem[112382] = 16'b0000000000000000;
	sram_mem[112383] = 16'b0000000000000000;
	sram_mem[112384] = 16'b0000000000000000;
	sram_mem[112385] = 16'b0000000000000000;
	sram_mem[112386] = 16'b0000000000000000;
	sram_mem[112387] = 16'b0000000000000000;
	sram_mem[112388] = 16'b0000000000000000;
	sram_mem[112389] = 16'b0000000000000000;
	sram_mem[112390] = 16'b0000000000000000;
	sram_mem[112391] = 16'b0000000000000000;
	sram_mem[112392] = 16'b0000000000000000;
	sram_mem[112393] = 16'b0000000000000000;
	sram_mem[112394] = 16'b0000000000000000;
	sram_mem[112395] = 16'b0000000000000000;
	sram_mem[112396] = 16'b0000000000000000;
	sram_mem[112397] = 16'b0000000000000000;
	sram_mem[112398] = 16'b0000000000000000;
	sram_mem[112399] = 16'b0000000000000000;
	sram_mem[112400] = 16'b0000000000000000;
	sram_mem[112401] = 16'b0000000000000000;
	sram_mem[112402] = 16'b0000000000000000;
	sram_mem[112403] = 16'b0000000000000000;
	sram_mem[112404] = 16'b0000000000000000;
	sram_mem[112405] = 16'b0000000000000000;
	sram_mem[112406] = 16'b0000000000000000;
	sram_mem[112407] = 16'b0000000000000000;
	sram_mem[112408] = 16'b0000000000000000;
	sram_mem[112409] = 16'b0000000000000000;
	sram_mem[112410] = 16'b0000000000000000;
	sram_mem[112411] = 16'b0000000000000000;
	sram_mem[112412] = 16'b0000000000000000;
	sram_mem[112413] = 16'b0000000000000000;
	sram_mem[112414] = 16'b0000000000000000;
	sram_mem[112415] = 16'b0000000000000000;
	sram_mem[112416] = 16'b0000000000000000;
	sram_mem[112417] = 16'b0000000000000000;
	sram_mem[112418] = 16'b0000000000000000;
	sram_mem[112419] = 16'b0000000000000000;
	sram_mem[112420] = 16'b0000000000000000;
	sram_mem[112421] = 16'b0000000000000000;
	sram_mem[112422] = 16'b0000000000000000;
	sram_mem[112423] = 16'b0000000000000000;
	sram_mem[112424] = 16'b0000000000000000;
	sram_mem[112425] = 16'b0000000000000000;
	sram_mem[112426] = 16'b0000000000000000;
	sram_mem[112427] = 16'b0000000000000000;
	sram_mem[112428] = 16'b0000000000000000;
	sram_mem[112429] = 16'b0000000000000000;
	sram_mem[112430] = 16'b0000000000000000;
	sram_mem[112431] = 16'b0000000000000000;
	sram_mem[112432] = 16'b0000000000000000;
	sram_mem[112433] = 16'b0000000000000000;
	sram_mem[112434] = 16'b0000000000000000;
	sram_mem[112435] = 16'b0000000000000000;
	sram_mem[112436] = 16'b0000000000000000;
	sram_mem[112437] = 16'b0000000000000000;
	sram_mem[112438] = 16'b0000000000000000;
	sram_mem[112439] = 16'b0000000000000000;
	sram_mem[112440] = 16'b0000000000000000;
	sram_mem[112441] = 16'b0000000000000000;
	sram_mem[112442] = 16'b0000000000000000;
	sram_mem[112443] = 16'b0000000000000000;
	sram_mem[112444] = 16'b0000000000000000;
	sram_mem[112445] = 16'b0000000000000000;
	sram_mem[112446] = 16'b0000000000000000;
	sram_mem[112447] = 16'b0000000000000000;
	sram_mem[112448] = 16'b0000000000000000;
	sram_mem[112449] = 16'b0000000000000000;
	sram_mem[112450] = 16'b0000000000000000;
	sram_mem[112451] = 16'b0000000000000000;
	sram_mem[112452] = 16'b0000000000000000;
	sram_mem[112453] = 16'b0000000000000000;
	sram_mem[112454] = 16'b0000000000000000;
	sram_mem[112455] = 16'b0000000000000000;
	sram_mem[112456] = 16'b0000000000000000;
	sram_mem[112457] = 16'b0000000000000000;
	sram_mem[112458] = 16'b0000000000000000;
	sram_mem[112459] = 16'b0000000000000000;
	sram_mem[112460] = 16'b0000000000000000;
	sram_mem[112461] = 16'b0000000000000000;
	sram_mem[112462] = 16'b0000000000000000;
	sram_mem[112463] = 16'b0000000000000000;
	sram_mem[112464] = 16'b0000000000000000;
	sram_mem[112465] = 16'b0000000000000000;
	sram_mem[112466] = 16'b0000000000000000;
	sram_mem[112467] = 16'b0000000000000000;
	sram_mem[112468] = 16'b0000000000000000;
	sram_mem[112469] = 16'b0000000000000000;
	sram_mem[112470] = 16'b0000000000000000;
	sram_mem[112471] = 16'b0000000000000000;
	sram_mem[112472] = 16'b0000000000000000;
	sram_mem[112473] = 16'b0000000000000000;
	sram_mem[112474] = 16'b0000000000000000;
	sram_mem[112475] = 16'b0000000000000000;
	sram_mem[112476] = 16'b0000000000000000;
	sram_mem[112477] = 16'b0000000000000000;
	sram_mem[112478] = 16'b0000000000000000;
	sram_mem[112479] = 16'b0000000000000000;
	sram_mem[112480] = 16'b0000000000000000;
	sram_mem[112481] = 16'b0000000000000000;
	sram_mem[112482] = 16'b0000000000000000;
	sram_mem[112483] = 16'b0000000000000000;
	sram_mem[112484] = 16'b0000000000000000;
	sram_mem[112485] = 16'b0000000000000000;
	sram_mem[112486] = 16'b0000000000000000;
	sram_mem[112487] = 16'b0000000000000000;
	sram_mem[112488] = 16'b0000000000000000;
	sram_mem[112489] = 16'b0000000000000000;
	sram_mem[112490] = 16'b0000000000000000;
	sram_mem[112491] = 16'b0000000000000000;
	sram_mem[112492] = 16'b0000000000000000;
	sram_mem[112493] = 16'b0000000000000000;
	sram_mem[112494] = 16'b0000000000000000;
	sram_mem[112495] = 16'b0000000000000000;
	sram_mem[112496] = 16'b0000000000000000;
	sram_mem[112497] = 16'b0000000000000000;
	sram_mem[112498] = 16'b0000000000000000;
	sram_mem[112499] = 16'b0000000000000000;
	sram_mem[112500] = 16'b0000000000000000;
	sram_mem[112501] = 16'b0000000000000000;
	sram_mem[112502] = 16'b0000000000000000;
	sram_mem[112503] = 16'b0000000000000000;
	sram_mem[112504] = 16'b0000000000000000;
	sram_mem[112505] = 16'b0000000000000000;
	sram_mem[112506] = 16'b0000000000000000;
	sram_mem[112507] = 16'b0000000000000000;
	sram_mem[112508] = 16'b0000000000000000;
	sram_mem[112509] = 16'b0000000000000000;
	sram_mem[112510] = 16'b0000000000000000;
	sram_mem[112511] = 16'b0000000000000000;
	sram_mem[112512] = 16'b0000000000000000;
	sram_mem[112513] = 16'b0000000000000000;
	sram_mem[112514] = 16'b0000000000000000;
	sram_mem[112515] = 16'b0000000000000000;
	sram_mem[112516] = 16'b0000000000000000;
	sram_mem[112517] = 16'b0000000000000000;
	sram_mem[112518] = 16'b0000000000000000;
	sram_mem[112519] = 16'b0000000000000000;
	sram_mem[112520] = 16'b0000000000000000;
	sram_mem[112521] = 16'b0000000000000000;
	sram_mem[112522] = 16'b0000000000000000;
	sram_mem[112523] = 16'b0000000000000000;
	sram_mem[112524] = 16'b0000000000000000;
	sram_mem[112525] = 16'b0000000000000000;
	sram_mem[112526] = 16'b0000000000000000;
	sram_mem[112527] = 16'b0000000000000000;
	sram_mem[112528] = 16'b0000000000000000;
	sram_mem[112529] = 16'b0000000000000000;
	sram_mem[112530] = 16'b0000000000000000;
	sram_mem[112531] = 16'b0000000000000000;
	sram_mem[112532] = 16'b0000000000000000;
	sram_mem[112533] = 16'b0000000000000000;
	sram_mem[112534] = 16'b0000000000000000;
	sram_mem[112535] = 16'b0000000000000000;
	sram_mem[112536] = 16'b0000000000000000;
	sram_mem[112537] = 16'b0000000000000000;
	sram_mem[112538] = 16'b0000000000000000;
	sram_mem[112539] = 16'b0000000000000000;
	sram_mem[112540] = 16'b0000000000000000;
	sram_mem[112541] = 16'b0000000000000000;
	sram_mem[112542] = 16'b0000000000000000;
	sram_mem[112543] = 16'b0000000000000000;
	sram_mem[112544] = 16'b0000000000000000;
	sram_mem[112545] = 16'b0000000000000000;
	sram_mem[112546] = 16'b0000000000000000;
	sram_mem[112547] = 16'b0000000000000000;
	sram_mem[112548] = 16'b0000000000000000;
	sram_mem[112549] = 16'b0000000000000000;
	sram_mem[112550] = 16'b0000000000000000;
	sram_mem[112551] = 16'b0000000000000000;
	sram_mem[112552] = 16'b0000000000000000;
	sram_mem[112553] = 16'b0000000000000000;
	sram_mem[112554] = 16'b0000000000000000;
	sram_mem[112555] = 16'b0000000000000000;
	sram_mem[112556] = 16'b0000000000000000;
	sram_mem[112557] = 16'b0000000000000000;
	sram_mem[112558] = 16'b0000000000000000;
	sram_mem[112559] = 16'b0000000000000000;
	sram_mem[112560] = 16'b0000000000000000;
	sram_mem[112561] = 16'b0000000000000000;
	sram_mem[112562] = 16'b0000000000000000;
	sram_mem[112563] = 16'b0000000000000000;
	sram_mem[112564] = 16'b0000000000000000;
	sram_mem[112565] = 16'b0000000000000000;
	sram_mem[112566] = 16'b0000000000000000;
	sram_mem[112567] = 16'b0000000000000000;
	sram_mem[112568] = 16'b0000000000000000;
	sram_mem[112569] = 16'b0000000000000000;
	sram_mem[112570] = 16'b0000000000000000;
	sram_mem[112571] = 16'b0000000000000000;
	sram_mem[112572] = 16'b0000000000000000;
	sram_mem[112573] = 16'b0000000000000000;
	sram_mem[112574] = 16'b0000000000000000;
	sram_mem[112575] = 16'b0000000000000000;
	sram_mem[112576] = 16'b0000000000000000;
	sram_mem[112577] = 16'b0000000000000000;
	sram_mem[112578] = 16'b0000000000000000;
	sram_mem[112579] = 16'b0000000000000000;
	sram_mem[112580] = 16'b0000000000000000;
	sram_mem[112581] = 16'b0000000000000000;
	sram_mem[112582] = 16'b0000000000000000;
	sram_mem[112583] = 16'b0000000000000000;
	sram_mem[112584] = 16'b0000000000000000;
	sram_mem[112585] = 16'b0000000000000000;
	sram_mem[112586] = 16'b0000000000000000;
	sram_mem[112587] = 16'b0000000000000000;
	sram_mem[112588] = 16'b0000000000000000;
	sram_mem[112589] = 16'b0000000000000000;
	sram_mem[112590] = 16'b0000000000000000;
	sram_mem[112591] = 16'b0000000000000000;
	sram_mem[112592] = 16'b0000000000000000;
	sram_mem[112593] = 16'b0000000000000000;
	sram_mem[112594] = 16'b0000000000000000;
	sram_mem[112595] = 16'b0000000000000000;
	sram_mem[112596] = 16'b0000000000000000;
	sram_mem[112597] = 16'b0000000000000000;
	sram_mem[112598] = 16'b0000000000000000;
	sram_mem[112599] = 16'b0000000000000000;
	sram_mem[112600] = 16'b0000000000000000;
	sram_mem[112601] = 16'b0000000000000000;
	sram_mem[112602] = 16'b0000000000000000;
	sram_mem[112603] = 16'b0000000000000000;
	sram_mem[112604] = 16'b0000000000000000;
	sram_mem[112605] = 16'b0000000000000000;
	sram_mem[112606] = 16'b0000000000000000;
	sram_mem[112607] = 16'b0000000000000000;
	sram_mem[112608] = 16'b0000000000000000;
	sram_mem[112609] = 16'b0000000000000000;
	sram_mem[112610] = 16'b0000000000000000;
	sram_mem[112611] = 16'b0000000000000000;
	sram_mem[112612] = 16'b0000000000000000;
	sram_mem[112613] = 16'b0000000000000000;
	sram_mem[112614] = 16'b0000000000000000;
	sram_mem[112615] = 16'b0000000000000000;
	sram_mem[112616] = 16'b0000000000000000;
	sram_mem[112617] = 16'b0000000000000000;
	sram_mem[112618] = 16'b0000000000000000;
	sram_mem[112619] = 16'b0000000000000000;
	sram_mem[112620] = 16'b0000000000000000;
	sram_mem[112621] = 16'b0000000000000000;
	sram_mem[112622] = 16'b0000000000000000;
	sram_mem[112623] = 16'b0000000000000000;
	sram_mem[112624] = 16'b0000000000000000;
	sram_mem[112625] = 16'b0000000000000000;
	sram_mem[112626] = 16'b0000000000000000;
	sram_mem[112627] = 16'b0000000000000000;
	sram_mem[112628] = 16'b0000000000000000;
	sram_mem[112629] = 16'b0000000000000000;
	sram_mem[112630] = 16'b0000000000000000;
	sram_mem[112631] = 16'b0000000000000000;
	sram_mem[112632] = 16'b0000000000000000;
	sram_mem[112633] = 16'b0000000000000000;
	sram_mem[112634] = 16'b0000000000000000;
	sram_mem[112635] = 16'b0000000000000000;
	sram_mem[112636] = 16'b0000000000000000;
	sram_mem[112637] = 16'b0000000000000000;
	sram_mem[112638] = 16'b0000000000000000;
	sram_mem[112639] = 16'b0000000000000000;
	sram_mem[112640] = 16'b0000000000000000;
	sram_mem[112641] = 16'b0000000000000000;
	sram_mem[112642] = 16'b0000000000000000;
	sram_mem[112643] = 16'b0000000000000000;
	sram_mem[112644] = 16'b0000000000000000;
	sram_mem[112645] = 16'b0000000000000000;
	sram_mem[112646] = 16'b0000000000000000;
	sram_mem[112647] = 16'b0000000000000000;
	sram_mem[112648] = 16'b0000000000000000;
	sram_mem[112649] = 16'b0000000000000000;
	sram_mem[112650] = 16'b0000000000000000;
	sram_mem[112651] = 16'b0000000000000000;
	sram_mem[112652] = 16'b0000000000000000;
	sram_mem[112653] = 16'b0000000000000000;
	sram_mem[112654] = 16'b0000000000000000;
	sram_mem[112655] = 16'b0000000000000000;
	sram_mem[112656] = 16'b0000000000000000;
	sram_mem[112657] = 16'b0000000000000000;
	sram_mem[112658] = 16'b0000000000000000;
	sram_mem[112659] = 16'b0000000000000000;
	sram_mem[112660] = 16'b0000000000000000;
	sram_mem[112661] = 16'b0000000000000000;
	sram_mem[112662] = 16'b0000000000000000;
	sram_mem[112663] = 16'b0000000000000000;
	sram_mem[112664] = 16'b0000000000000000;
	sram_mem[112665] = 16'b0000000000000000;
	sram_mem[112666] = 16'b0000000000000000;
	sram_mem[112667] = 16'b0000000000000000;
	sram_mem[112668] = 16'b0000000000000000;
	sram_mem[112669] = 16'b0000000000000000;
	sram_mem[112670] = 16'b0000000000000000;
	sram_mem[112671] = 16'b0000000000000000;
	sram_mem[112672] = 16'b0000000000000000;
	sram_mem[112673] = 16'b0000000000000000;
	sram_mem[112674] = 16'b0000000000000000;
	sram_mem[112675] = 16'b0000000000000000;
	sram_mem[112676] = 16'b0000000000000000;
	sram_mem[112677] = 16'b0000000000000000;
	sram_mem[112678] = 16'b0000000000000000;
	sram_mem[112679] = 16'b0000000000000000;
	sram_mem[112680] = 16'b0000000000000000;
	sram_mem[112681] = 16'b0000000000000000;
	sram_mem[112682] = 16'b0000000000000000;
	sram_mem[112683] = 16'b0000000000000000;
	sram_mem[112684] = 16'b0000000000000000;
	sram_mem[112685] = 16'b0000000000000000;
	sram_mem[112686] = 16'b0000000000000000;
	sram_mem[112687] = 16'b0000000000000000;
	sram_mem[112688] = 16'b0000000000000000;
	sram_mem[112689] = 16'b0000000000000000;
	sram_mem[112690] = 16'b0000000000000000;
	sram_mem[112691] = 16'b0000000000000000;
	sram_mem[112692] = 16'b0000000000000000;
	sram_mem[112693] = 16'b0000000000000000;
	sram_mem[112694] = 16'b0000000000000000;
	sram_mem[112695] = 16'b0000000000000000;
	sram_mem[112696] = 16'b0000000000000000;
	sram_mem[112697] = 16'b0000000000000000;
	sram_mem[112698] = 16'b0000000000000000;
	sram_mem[112699] = 16'b0000000000000000;
	sram_mem[112700] = 16'b0000000000000000;
	sram_mem[112701] = 16'b0000000000000000;
	sram_mem[112702] = 16'b0000000000000000;
	sram_mem[112703] = 16'b0000000000000000;
	sram_mem[112704] = 16'b0000000000000000;
	sram_mem[112705] = 16'b0000000000000000;
	sram_mem[112706] = 16'b0000000000000000;
	sram_mem[112707] = 16'b0000000000000000;
	sram_mem[112708] = 16'b0000000000000000;
	sram_mem[112709] = 16'b0000000000000000;
	sram_mem[112710] = 16'b0000000000000000;
	sram_mem[112711] = 16'b0000000000000000;
	sram_mem[112712] = 16'b0000000000000000;
	sram_mem[112713] = 16'b0000000000000000;
	sram_mem[112714] = 16'b0000000000000000;
	sram_mem[112715] = 16'b0000000000000000;
	sram_mem[112716] = 16'b0000000000000000;
	sram_mem[112717] = 16'b0000000000000000;
	sram_mem[112718] = 16'b0000000000000000;
	sram_mem[112719] = 16'b0000000000000000;
	sram_mem[112720] = 16'b0000000000000000;
	sram_mem[112721] = 16'b0000000000000000;
	sram_mem[112722] = 16'b0000000000000000;
	sram_mem[112723] = 16'b0000000000000000;
	sram_mem[112724] = 16'b0000000000000000;
	sram_mem[112725] = 16'b0000000000000000;
	sram_mem[112726] = 16'b0000000000000000;
	sram_mem[112727] = 16'b0000000000000000;
	sram_mem[112728] = 16'b0000000000000000;
	sram_mem[112729] = 16'b0000000000000000;
	sram_mem[112730] = 16'b0000000000000000;
	sram_mem[112731] = 16'b0000000000000000;
	sram_mem[112732] = 16'b0000000000000000;
	sram_mem[112733] = 16'b0000000000000000;
	sram_mem[112734] = 16'b0000000000000000;
	sram_mem[112735] = 16'b0000000000000000;
	sram_mem[112736] = 16'b0000000000000000;
	sram_mem[112737] = 16'b0000000000000000;
	sram_mem[112738] = 16'b0000000000000000;
	sram_mem[112739] = 16'b0000000000000000;
	sram_mem[112740] = 16'b0000000000000000;
	sram_mem[112741] = 16'b0000000000000000;
	sram_mem[112742] = 16'b0000000000000000;
	sram_mem[112743] = 16'b0000000000000000;
	sram_mem[112744] = 16'b0000000000000000;
	sram_mem[112745] = 16'b0000000000000000;
	sram_mem[112746] = 16'b0000000000000000;
	sram_mem[112747] = 16'b0000000000000000;
	sram_mem[112748] = 16'b0000000000000000;
	sram_mem[112749] = 16'b0000000000000000;
	sram_mem[112750] = 16'b0000000000000000;
	sram_mem[112751] = 16'b0000000000000000;
	sram_mem[112752] = 16'b0000000000000000;
	sram_mem[112753] = 16'b0000000000000000;
	sram_mem[112754] = 16'b0000000000000000;
	sram_mem[112755] = 16'b0000000000000000;
	sram_mem[112756] = 16'b0000000000000000;
	sram_mem[112757] = 16'b0000000000000000;
	sram_mem[112758] = 16'b0000000000000000;
	sram_mem[112759] = 16'b0000000000000000;
	sram_mem[112760] = 16'b0000000000000000;
	sram_mem[112761] = 16'b0000000000000000;
	sram_mem[112762] = 16'b0000000000000000;
	sram_mem[112763] = 16'b0000000000000000;
	sram_mem[112764] = 16'b0000000000000000;
	sram_mem[112765] = 16'b0000000000000000;
	sram_mem[112766] = 16'b0000000000000000;
	sram_mem[112767] = 16'b0000000000000000;
	sram_mem[112768] = 16'b0000000000000000;
	sram_mem[112769] = 16'b0000000000000000;
	sram_mem[112770] = 16'b0000000000000000;
	sram_mem[112771] = 16'b0000000000000000;
	sram_mem[112772] = 16'b0000000000000000;
	sram_mem[112773] = 16'b0000000000000000;
	sram_mem[112774] = 16'b0000000000000000;
	sram_mem[112775] = 16'b0000000000000000;
	sram_mem[112776] = 16'b0000000000000000;
	sram_mem[112777] = 16'b0000000000000000;
	sram_mem[112778] = 16'b0000000000000000;
	sram_mem[112779] = 16'b0000000000000000;
	sram_mem[112780] = 16'b0000000000000000;
	sram_mem[112781] = 16'b0000000000000000;
	sram_mem[112782] = 16'b0000000000000000;
	sram_mem[112783] = 16'b0000000000000000;
	sram_mem[112784] = 16'b0000000000000000;
	sram_mem[112785] = 16'b0000000000000000;
	sram_mem[112786] = 16'b0000000000000000;
	sram_mem[112787] = 16'b0000000000000000;
	sram_mem[112788] = 16'b0000000000000000;
	sram_mem[112789] = 16'b0000000000000000;
	sram_mem[112790] = 16'b0000000000000000;
	sram_mem[112791] = 16'b0000000000000000;
	sram_mem[112792] = 16'b0000000000000000;
	sram_mem[112793] = 16'b0000000000000000;
	sram_mem[112794] = 16'b0000000000000000;
	sram_mem[112795] = 16'b0000000000000000;
	sram_mem[112796] = 16'b0000000000000000;
	sram_mem[112797] = 16'b0000000000000000;
	sram_mem[112798] = 16'b0000000000000000;
	sram_mem[112799] = 16'b0000000000000000;
	sram_mem[112800] = 16'b0000000000000000;
	sram_mem[112801] = 16'b0000000000000000;
	sram_mem[112802] = 16'b0000000000000000;
	sram_mem[112803] = 16'b0000000000000000;
	sram_mem[112804] = 16'b0000000000000000;
	sram_mem[112805] = 16'b0000000000000000;
	sram_mem[112806] = 16'b0000000000000000;
	sram_mem[112807] = 16'b0000000000000000;
	sram_mem[112808] = 16'b0000000000000000;
	sram_mem[112809] = 16'b0000000000000000;
	sram_mem[112810] = 16'b0000000000000000;
	sram_mem[112811] = 16'b0000000000000000;
	sram_mem[112812] = 16'b0000000000000000;
	sram_mem[112813] = 16'b0000000000000000;
	sram_mem[112814] = 16'b0000000000000000;
	sram_mem[112815] = 16'b0000000000000000;
	sram_mem[112816] = 16'b0000000000000000;
	sram_mem[112817] = 16'b0000000000000000;
	sram_mem[112818] = 16'b0000000000000000;
	sram_mem[112819] = 16'b0000000000000000;
	sram_mem[112820] = 16'b0000000000000000;
	sram_mem[112821] = 16'b0000000000000000;
	sram_mem[112822] = 16'b0000000000000000;
	sram_mem[112823] = 16'b0000000000000000;
	sram_mem[112824] = 16'b0000000000000000;
	sram_mem[112825] = 16'b0000000000000000;
	sram_mem[112826] = 16'b0000000000000000;
	sram_mem[112827] = 16'b0000000000000000;
	sram_mem[112828] = 16'b0000000000000000;
	sram_mem[112829] = 16'b0000000000000000;
	sram_mem[112830] = 16'b0000000000000000;
	sram_mem[112831] = 16'b0000000000000000;
	sram_mem[112832] = 16'b0000000000000000;
	sram_mem[112833] = 16'b0000000000000000;
	sram_mem[112834] = 16'b0000000000000000;
	sram_mem[112835] = 16'b0000000000000000;
	sram_mem[112836] = 16'b0000000000000000;
	sram_mem[112837] = 16'b0000000000000000;
	sram_mem[112838] = 16'b0000000000000000;
	sram_mem[112839] = 16'b0000000000000000;
	sram_mem[112840] = 16'b0000000000000000;
	sram_mem[112841] = 16'b0000000000000000;
	sram_mem[112842] = 16'b0000000000000000;
	sram_mem[112843] = 16'b0000000000000000;
	sram_mem[112844] = 16'b0000000000000000;
	sram_mem[112845] = 16'b0000000000000000;
	sram_mem[112846] = 16'b0000000000000000;
	sram_mem[112847] = 16'b0000000000000000;
	sram_mem[112848] = 16'b0000000000000000;
	sram_mem[112849] = 16'b0000000000000000;
	sram_mem[112850] = 16'b0000000000000000;
	sram_mem[112851] = 16'b0000000000000000;
	sram_mem[112852] = 16'b0000000000000000;
	sram_mem[112853] = 16'b0000000000000000;
	sram_mem[112854] = 16'b0000000000000000;
	sram_mem[112855] = 16'b0000000000000000;
	sram_mem[112856] = 16'b0000000000000000;
	sram_mem[112857] = 16'b0000000000000000;
	sram_mem[112858] = 16'b0000000000000000;
	sram_mem[112859] = 16'b0000000000000000;
	sram_mem[112860] = 16'b0000000000000000;
	sram_mem[112861] = 16'b0000000000000000;
	sram_mem[112862] = 16'b0000000000000000;
	sram_mem[112863] = 16'b0000000000000000;
	sram_mem[112864] = 16'b0000000000000000;
	sram_mem[112865] = 16'b0000000000000000;
	sram_mem[112866] = 16'b0000000000000000;
	sram_mem[112867] = 16'b0000000000000000;
	sram_mem[112868] = 16'b0000000000000000;
	sram_mem[112869] = 16'b0000000000000000;
	sram_mem[112870] = 16'b0000000000000000;
	sram_mem[112871] = 16'b0000000000000000;
	sram_mem[112872] = 16'b0000000000000000;
	sram_mem[112873] = 16'b0000000000000000;
	sram_mem[112874] = 16'b0000000000000000;
	sram_mem[112875] = 16'b0000000000000000;
	sram_mem[112876] = 16'b0000000000000000;
	sram_mem[112877] = 16'b0000000000000000;
	sram_mem[112878] = 16'b0000000000000000;
	sram_mem[112879] = 16'b0000000000000000;
	sram_mem[112880] = 16'b0000000000000000;
	sram_mem[112881] = 16'b0000000000000000;
	sram_mem[112882] = 16'b0000000000000000;
	sram_mem[112883] = 16'b0000000000000000;
	sram_mem[112884] = 16'b0000000000000000;
	sram_mem[112885] = 16'b0000000000000000;
	sram_mem[112886] = 16'b0000000000000000;
	sram_mem[112887] = 16'b0000000000000000;
	sram_mem[112888] = 16'b0000000000000000;
	sram_mem[112889] = 16'b0000000000000000;
	sram_mem[112890] = 16'b0000000000000000;
	sram_mem[112891] = 16'b0000000000000000;
	sram_mem[112892] = 16'b0000000000000000;
	sram_mem[112893] = 16'b0000000000000000;
	sram_mem[112894] = 16'b0000000000000000;
	sram_mem[112895] = 16'b0000000000000000;
	sram_mem[112896] = 16'b0000000000000000;
	sram_mem[112897] = 16'b0000000000000000;
	sram_mem[112898] = 16'b0000000000000000;
	sram_mem[112899] = 16'b0000000000000000;
	sram_mem[112900] = 16'b0000000000000000;
	sram_mem[112901] = 16'b0000000000000000;
	sram_mem[112902] = 16'b0000000000000000;
	sram_mem[112903] = 16'b0000000000000000;
	sram_mem[112904] = 16'b0000000000000000;
	sram_mem[112905] = 16'b0000000000000000;
	sram_mem[112906] = 16'b0000000000000000;
	sram_mem[112907] = 16'b0000000000000000;
	sram_mem[112908] = 16'b0000000000000000;
	sram_mem[112909] = 16'b0000000000000000;
	sram_mem[112910] = 16'b0000000000000000;
	sram_mem[112911] = 16'b0000000000000000;
	sram_mem[112912] = 16'b0000000000000000;
	sram_mem[112913] = 16'b0000000000000000;
	sram_mem[112914] = 16'b0000000000000000;
	sram_mem[112915] = 16'b0000000000000000;
	sram_mem[112916] = 16'b0000000000000000;
	sram_mem[112917] = 16'b0000000000000000;
	sram_mem[112918] = 16'b0000000000000000;
	sram_mem[112919] = 16'b0000000000000000;
	sram_mem[112920] = 16'b0000000000000000;
	sram_mem[112921] = 16'b0000000000000000;
	sram_mem[112922] = 16'b0000000000000000;
	sram_mem[112923] = 16'b0000000000000000;
	sram_mem[112924] = 16'b0000000000000000;
	sram_mem[112925] = 16'b0000000000000000;
	sram_mem[112926] = 16'b0000000000000000;
	sram_mem[112927] = 16'b0000000000000000;
	sram_mem[112928] = 16'b0000000000000000;
	sram_mem[112929] = 16'b0000000000000000;
	sram_mem[112930] = 16'b0000000000000000;
	sram_mem[112931] = 16'b0000000000000000;
	sram_mem[112932] = 16'b0000000000000000;
	sram_mem[112933] = 16'b0000000000000000;
	sram_mem[112934] = 16'b0000000000000000;
	sram_mem[112935] = 16'b0000000000000000;
	sram_mem[112936] = 16'b0000000000000000;
	sram_mem[112937] = 16'b0000000000000000;
	sram_mem[112938] = 16'b0000000000000000;
	sram_mem[112939] = 16'b0000000000000000;
	sram_mem[112940] = 16'b0000000000000000;
	sram_mem[112941] = 16'b0000000000000000;
	sram_mem[112942] = 16'b0000000000000000;
	sram_mem[112943] = 16'b0000000000000000;
	sram_mem[112944] = 16'b0000000000000000;
	sram_mem[112945] = 16'b0000000000000000;
	sram_mem[112946] = 16'b0000000000000000;
	sram_mem[112947] = 16'b0000000000000000;
	sram_mem[112948] = 16'b0000000000000000;
	sram_mem[112949] = 16'b0000000000000000;
	sram_mem[112950] = 16'b0000000000000000;
	sram_mem[112951] = 16'b0000000000000000;
	sram_mem[112952] = 16'b0000000000000000;
	sram_mem[112953] = 16'b0000000000000000;
	sram_mem[112954] = 16'b0000000000000000;
	sram_mem[112955] = 16'b0000000000000000;
	sram_mem[112956] = 16'b0000000000000000;
	sram_mem[112957] = 16'b0000000000000000;
	sram_mem[112958] = 16'b0000000000000000;
	sram_mem[112959] = 16'b0000000000000000;
	sram_mem[112960] = 16'b0000000000000000;
	sram_mem[112961] = 16'b0000000000000000;
	sram_mem[112962] = 16'b0000000000000000;
	sram_mem[112963] = 16'b0000000000000000;
	sram_mem[112964] = 16'b0000000000000000;
	sram_mem[112965] = 16'b0000000000000000;
	sram_mem[112966] = 16'b0000000000000000;
	sram_mem[112967] = 16'b0000000000000000;
	sram_mem[112968] = 16'b0000000000000000;
	sram_mem[112969] = 16'b0000000000000000;
	sram_mem[112970] = 16'b0000000000000000;
	sram_mem[112971] = 16'b0000000000000000;
	sram_mem[112972] = 16'b0000000000000000;
	sram_mem[112973] = 16'b0000000000000000;
	sram_mem[112974] = 16'b0000000000000000;
	sram_mem[112975] = 16'b0000000000000000;
	sram_mem[112976] = 16'b0000000000000000;
	sram_mem[112977] = 16'b0000000000000000;
	sram_mem[112978] = 16'b0000000000000000;
	sram_mem[112979] = 16'b0000000000000000;
	sram_mem[112980] = 16'b0000000000000000;
	sram_mem[112981] = 16'b0000000000000000;
	sram_mem[112982] = 16'b0000000000000000;
	sram_mem[112983] = 16'b0000000000000000;
	sram_mem[112984] = 16'b0000000000000000;
	sram_mem[112985] = 16'b0000000000000000;
	sram_mem[112986] = 16'b0000000000000000;
	sram_mem[112987] = 16'b0000000000000000;
	sram_mem[112988] = 16'b0000000000000000;
	sram_mem[112989] = 16'b0000000000000000;
	sram_mem[112990] = 16'b0000000000000000;
	sram_mem[112991] = 16'b0000000000000000;
	sram_mem[112992] = 16'b0000000000000000;
	sram_mem[112993] = 16'b0000000000000000;
	sram_mem[112994] = 16'b0000000000000000;
	sram_mem[112995] = 16'b0000000000000000;
	sram_mem[112996] = 16'b0000000000000000;
	sram_mem[112997] = 16'b0000000000000000;
	sram_mem[112998] = 16'b0000000000000000;
	sram_mem[112999] = 16'b0000000000000000;
	sram_mem[113000] = 16'b0000000000000000;
	sram_mem[113001] = 16'b0000000000000000;
	sram_mem[113002] = 16'b0000000000000000;
	sram_mem[113003] = 16'b0000000000000000;
	sram_mem[113004] = 16'b0000000000000000;
	sram_mem[113005] = 16'b0000000000000000;
	sram_mem[113006] = 16'b0000000000000000;
	sram_mem[113007] = 16'b0000000000000000;
	sram_mem[113008] = 16'b0000000000000000;
	sram_mem[113009] = 16'b0000000000000000;
	sram_mem[113010] = 16'b0000000000000000;
	sram_mem[113011] = 16'b0000000000000000;
	sram_mem[113012] = 16'b0000000000000000;
	sram_mem[113013] = 16'b0000000000000000;
	sram_mem[113014] = 16'b0000000000000000;
	sram_mem[113015] = 16'b0000000000000000;
	sram_mem[113016] = 16'b0000000000000000;
	sram_mem[113017] = 16'b0000000000000000;
	sram_mem[113018] = 16'b0000000000000000;
	sram_mem[113019] = 16'b0000000000000000;
	sram_mem[113020] = 16'b0000000000000000;
	sram_mem[113021] = 16'b0000000000000000;
	sram_mem[113022] = 16'b0000000000000000;
	sram_mem[113023] = 16'b0000000000000000;
	sram_mem[113024] = 16'b0000000000000000;
	sram_mem[113025] = 16'b0000000000000000;
	sram_mem[113026] = 16'b0000000000000000;
	sram_mem[113027] = 16'b0000000000000000;
	sram_mem[113028] = 16'b0000000000000000;
	sram_mem[113029] = 16'b0000000000000000;
	sram_mem[113030] = 16'b0000000000000000;
	sram_mem[113031] = 16'b0000000000000000;
	sram_mem[113032] = 16'b0000000000000000;
	sram_mem[113033] = 16'b0000000000000000;
	sram_mem[113034] = 16'b0000000000000000;
	sram_mem[113035] = 16'b0000000000000000;
	sram_mem[113036] = 16'b0000000000000000;
	sram_mem[113037] = 16'b0000000000000000;
	sram_mem[113038] = 16'b0000000000000000;
	sram_mem[113039] = 16'b0000000000000000;
	sram_mem[113040] = 16'b0000000000000000;
	sram_mem[113041] = 16'b0000000000000000;
	sram_mem[113042] = 16'b0000000000000000;
	sram_mem[113043] = 16'b0000000000000000;
	sram_mem[113044] = 16'b0000000000000000;
	sram_mem[113045] = 16'b0000000000000000;
	sram_mem[113046] = 16'b0000000000000000;
	sram_mem[113047] = 16'b0000000000000000;
	sram_mem[113048] = 16'b0000000000000000;
	sram_mem[113049] = 16'b0000000000000000;
	sram_mem[113050] = 16'b0000000000000000;
	sram_mem[113051] = 16'b0000000000000000;
	sram_mem[113052] = 16'b0000000000000000;
	sram_mem[113053] = 16'b0000000000000000;
	sram_mem[113054] = 16'b0000000000000000;
	sram_mem[113055] = 16'b0000000000000000;
	sram_mem[113056] = 16'b0000000000000000;
	sram_mem[113057] = 16'b0000000000000000;
	sram_mem[113058] = 16'b0000000000000000;
	sram_mem[113059] = 16'b0000000000000000;
	sram_mem[113060] = 16'b0000000000000000;
	sram_mem[113061] = 16'b0000000000000000;
	sram_mem[113062] = 16'b0000000000000000;
	sram_mem[113063] = 16'b0000000000000000;
	sram_mem[113064] = 16'b0000000000000000;
	sram_mem[113065] = 16'b0000000000000000;
	sram_mem[113066] = 16'b0000000000000000;
	sram_mem[113067] = 16'b0000000000000000;
	sram_mem[113068] = 16'b0000000000000000;
	sram_mem[113069] = 16'b0000000000000000;
	sram_mem[113070] = 16'b0000000000000000;
	sram_mem[113071] = 16'b0000000000000000;
	sram_mem[113072] = 16'b0000000000000000;
	sram_mem[113073] = 16'b0000000000000000;
	sram_mem[113074] = 16'b0000000000000000;
	sram_mem[113075] = 16'b0000000000000000;
	sram_mem[113076] = 16'b0000000000000000;
	sram_mem[113077] = 16'b0000000000000000;
	sram_mem[113078] = 16'b0000000000000000;
	sram_mem[113079] = 16'b0000000000000000;
	sram_mem[113080] = 16'b0000000000000000;
	sram_mem[113081] = 16'b0000000000000000;
	sram_mem[113082] = 16'b0000000000000000;
	sram_mem[113083] = 16'b0000000000000000;
	sram_mem[113084] = 16'b0000000000000000;
	sram_mem[113085] = 16'b0000000000000000;
	sram_mem[113086] = 16'b0000000000000000;
	sram_mem[113087] = 16'b0000000000000000;
	sram_mem[113088] = 16'b0000000000000000;
	sram_mem[113089] = 16'b0000000000000000;
	sram_mem[113090] = 16'b0000000000000000;
	sram_mem[113091] = 16'b0000000000000000;
	sram_mem[113092] = 16'b0000000000000000;
	sram_mem[113093] = 16'b0000000000000000;
	sram_mem[113094] = 16'b0000000000000000;
	sram_mem[113095] = 16'b0000000000000000;
	sram_mem[113096] = 16'b0000000000000000;
	sram_mem[113097] = 16'b0000000000000000;
	sram_mem[113098] = 16'b0000000000000000;
	sram_mem[113099] = 16'b0000000000000000;
	sram_mem[113100] = 16'b0000000000000000;
	sram_mem[113101] = 16'b0000000000000000;
	sram_mem[113102] = 16'b0000000000000000;
	sram_mem[113103] = 16'b0000000000000000;
	sram_mem[113104] = 16'b0000000000000000;
	sram_mem[113105] = 16'b0000000000000000;
	sram_mem[113106] = 16'b0000000000000000;
	sram_mem[113107] = 16'b0000000000000000;
	sram_mem[113108] = 16'b0000000000000000;
	sram_mem[113109] = 16'b0000000000000000;
	sram_mem[113110] = 16'b0000000000000000;
	sram_mem[113111] = 16'b0000000000000000;
	sram_mem[113112] = 16'b0000000000000000;
	sram_mem[113113] = 16'b0000000000000000;
	sram_mem[113114] = 16'b0000000000000000;
	sram_mem[113115] = 16'b0000000000000000;
	sram_mem[113116] = 16'b0000000000000000;
	sram_mem[113117] = 16'b0000000000000000;
	sram_mem[113118] = 16'b0000000000000000;
	sram_mem[113119] = 16'b0000000000000000;
	sram_mem[113120] = 16'b0000000000000000;
	sram_mem[113121] = 16'b0000000000000000;
	sram_mem[113122] = 16'b0000000000000000;
	sram_mem[113123] = 16'b0000000000000000;
	sram_mem[113124] = 16'b0000000000000000;
	sram_mem[113125] = 16'b0000000000000000;
	sram_mem[113126] = 16'b0000000000000000;
	sram_mem[113127] = 16'b0000000000000000;
	sram_mem[113128] = 16'b0000000000000000;
	sram_mem[113129] = 16'b0000000000000000;
	sram_mem[113130] = 16'b0000000000000000;
	sram_mem[113131] = 16'b0000000000000000;
	sram_mem[113132] = 16'b0000000000000000;
	sram_mem[113133] = 16'b0000000000000000;
	sram_mem[113134] = 16'b0000000000000000;
	sram_mem[113135] = 16'b0000000000000000;
	sram_mem[113136] = 16'b0000000000000000;
	sram_mem[113137] = 16'b0000000000000000;
	sram_mem[113138] = 16'b0000000000000000;
	sram_mem[113139] = 16'b0000000000000000;
	sram_mem[113140] = 16'b0000000000000000;
	sram_mem[113141] = 16'b0000000000000000;
	sram_mem[113142] = 16'b0000000000000000;
	sram_mem[113143] = 16'b0000000000000000;
	sram_mem[113144] = 16'b0000000000000000;
	sram_mem[113145] = 16'b0000000000000000;
	sram_mem[113146] = 16'b0000000000000000;
	sram_mem[113147] = 16'b0000000000000000;
	sram_mem[113148] = 16'b0000000000000000;
	sram_mem[113149] = 16'b0000000000000000;
	sram_mem[113150] = 16'b0000000000000000;
	sram_mem[113151] = 16'b0000000000000000;
	sram_mem[113152] = 16'b0000000000000000;
	sram_mem[113153] = 16'b0000000000000000;
	sram_mem[113154] = 16'b0000000000000000;
	sram_mem[113155] = 16'b0000000000000000;
	sram_mem[113156] = 16'b0000000000000000;
	sram_mem[113157] = 16'b0000000000000000;
	sram_mem[113158] = 16'b0000000000000000;
	sram_mem[113159] = 16'b0000000000000000;
	sram_mem[113160] = 16'b0000000000000000;
	sram_mem[113161] = 16'b0000000000000000;
	sram_mem[113162] = 16'b0000000000000000;
	sram_mem[113163] = 16'b0000000000000000;
	sram_mem[113164] = 16'b0000000000000000;
	sram_mem[113165] = 16'b0000000000000000;
	sram_mem[113166] = 16'b0000000000000000;
	sram_mem[113167] = 16'b0000000000000000;
	sram_mem[113168] = 16'b0000000000000000;
	sram_mem[113169] = 16'b0000000000000000;
	sram_mem[113170] = 16'b0000000000000000;
	sram_mem[113171] = 16'b0000000000000000;
	sram_mem[113172] = 16'b0000000000000000;
	sram_mem[113173] = 16'b0000000000000000;
	sram_mem[113174] = 16'b0000000000000000;
	sram_mem[113175] = 16'b0000000000000000;
	sram_mem[113176] = 16'b0000000000000000;
	sram_mem[113177] = 16'b0000000000000000;
	sram_mem[113178] = 16'b0000000000000000;
	sram_mem[113179] = 16'b0000000000000000;
	sram_mem[113180] = 16'b0000000000000000;
	sram_mem[113181] = 16'b0000000000000000;
	sram_mem[113182] = 16'b0000000000000000;
	sram_mem[113183] = 16'b0000000000000000;
	sram_mem[113184] = 16'b0000000000000000;
	sram_mem[113185] = 16'b0000000000000000;
	sram_mem[113186] = 16'b0000000000000000;
	sram_mem[113187] = 16'b0000000000000000;
	sram_mem[113188] = 16'b0000000000000000;
	sram_mem[113189] = 16'b0000000000000000;
	sram_mem[113190] = 16'b0000000000000000;
	sram_mem[113191] = 16'b0000000000000000;
	sram_mem[113192] = 16'b0000000000000000;
	sram_mem[113193] = 16'b0000000000000000;
	sram_mem[113194] = 16'b0000000000000000;
	sram_mem[113195] = 16'b0000000000000000;
	sram_mem[113196] = 16'b0000000000000000;
	sram_mem[113197] = 16'b0000000000000000;
	sram_mem[113198] = 16'b0000000000000000;
	sram_mem[113199] = 16'b0000000000000000;
	sram_mem[113200] = 16'b0000000000000000;
	sram_mem[113201] = 16'b0000000000000000;
	sram_mem[113202] = 16'b0000000000000000;
	sram_mem[113203] = 16'b0000000000000000;
	sram_mem[113204] = 16'b0000000000000000;
	sram_mem[113205] = 16'b0000000000000000;
	sram_mem[113206] = 16'b0000000000000000;
	sram_mem[113207] = 16'b0000000000000000;
	sram_mem[113208] = 16'b0000000000000000;
	sram_mem[113209] = 16'b0000000000000000;
	sram_mem[113210] = 16'b0000000000000000;
	sram_mem[113211] = 16'b0000000000000000;
	sram_mem[113212] = 16'b0000000000000000;
	sram_mem[113213] = 16'b0000000000000000;
	sram_mem[113214] = 16'b0000000000000000;
	sram_mem[113215] = 16'b0000000000000000;
	sram_mem[113216] = 16'b0000000000000000;
	sram_mem[113217] = 16'b0000000000000000;
	sram_mem[113218] = 16'b0000000000000000;
	sram_mem[113219] = 16'b0000000000000000;
	sram_mem[113220] = 16'b0000000000000000;
	sram_mem[113221] = 16'b0000000000000000;
	sram_mem[113222] = 16'b0000000000000000;
	sram_mem[113223] = 16'b0000000000000000;
	sram_mem[113224] = 16'b0000000000000000;
	sram_mem[113225] = 16'b0000000000000000;
	sram_mem[113226] = 16'b0000000000000000;
	sram_mem[113227] = 16'b0000000000000000;
	sram_mem[113228] = 16'b0000000000000000;
	sram_mem[113229] = 16'b0000000000000000;
	sram_mem[113230] = 16'b0000000000000000;
	sram_mem[113231] = 16'b0000000000000000;
	sram_mem[113232] = 16'b0000000000000000;
	sram_mem[113233] = 16'b0000000000000000;
	sram_mem[113234] = 16'b0000000000000000;
	sram_mem[113235] = 16'b0000000000000000;
	sram_mem[113236] = 16'b0000000000000000;
	sram_mem[113237] = 16'b0000000000000000;
	sram_mem[113238] = 16'b0000000000000000;
	sram_mem[113239] = 16'b0000000000000000;
	sram_mem[113240] = 16'b0000000000000000;
	sram_mem[113241] = 16'b0000000000000000;
	sram_mem[113242] = 16'b0000000000000000;
	sram_mem[113243] = 16'b0000000000000000;
	sram_mem[113244] = 16'b0000000000000000;
	sram_mem[113245] = 16'b0000000000000000;
	sram_mem[113246] = 16'b0000000000000000;
	sram_mem[113247] = 16'b0000000000000000;
	sram_mem[113248] = 16'b0000000000000000;
	sram_mem[113249] = 16'b0000000000000000;
	sram_mem[113250] = 16'b0000000000000000;
	sram_mem[113251] = 16'b0000000000000000;
	sram_mem[113252] = 16'b0000000000000000;
	sram_mem[113253] = 16'b0000000000000000;
	sram_mem[113254] = 16'b0000000000000000;
	sram_mem[113255] = 16'b0000000000000000;
	sram_mem[113256] = 16'b0000000000000000;
	sram_mem[113257] = 16'b0000000000000000;
	sram_mem[113258] = 16'b0000000000000000;
	sram_mem[113259] = 16'b0000000000000000;
	sram_mem[113260] = 16'b0000000000000000;
	sram_mem[113261] = 16'b0000000000000000;
	sram_mem[113262] = 16'b0000000000000000;
	sram_mem[113263] = 16'b0000000000000000;
	sram_mem[113264] = 16'b0000000000000000;
	sram_mem[113265] = 16'b0000000000000000;
	sram_mem[113266] = 16'b0000000000000000;
	sram_mem[113267] = 16'b0000000000000000;
	sram_mem[113268] = 16'b0000000000000000;
	sram_mem[113269] = 16'b0000000000000000;
	sram_mem[113270] = 16'b0000000000000000;
	sram_mem[113271] = 16'b0000000000000000;
	sram_mem[113272] = 16'b0000000000000000;
	sram_mem[113273] = 16'b0000000000000000;
	sram_mem[113274] = 16'b0000000000000000;
	sram_mem[113275] = 16'b0000000000000000;
	sram_mem[113276] = 16'b0000000000000000;
	sram_mem[113277] = 16'b0000000000000000;
	sram_mem[113278] = 16'b0000000000000000;
	sram_mem[113279] = 16'b0000000000000000;
	sram_mem[113280] = 16'b0000000000000000;
	sram_mem[113281] = 16'b0000000000000000;
	sram_mem[113282] = 16'b0000000000000000;
	sram_mem[113283] = 16'b0000000000000000;
	sram_mem[113284] = 16'b0000000000000000;
	sram_mem[113285] = 16'b0000000000000000;
	sram_mem[113286] = 16'b0000000000000000;
	sram_mem[113287] = 16'b0000000000000000;
	sram_mem[113288] = 16'b0000000000000000;
	sram_mem[113289] = 16'b0000000000000000;
	sram_mem[113290] = 16'b0000000000000000;
	sram_mem[113291] = 16'b0000000000000000;
	sram_mem[113292] = 16'b0000000000000000;
	sram_mem[113293] = 16'b0000000000000000;
	sram_mem[113294] = 16'b0000000000000000;
	sram_mem[113295] = 16'b0000000000000000;
	sram_mem[113296] = 16'b0000000000000000;
	sram_mem[113297] = 16'b0000000000000000;
	sram_mem[113298] = 16'b0000000000000000;
	sram_mem[113299] = 16'b0000000000000000;
	sram_mem[113300] = 16'b0000000000000000;
	sram_mem[113301] = 16'b0000000000000000;
	sram_mem[113302] = 16'b0000000000000000;
	sram_mem[113303] = 16'b0000000000000000;
	sram_mem[113304] = 16'b0000000000000000;
	sram_mem[113305] = 16'b0000000000000000;
	sram_mem[113306] = 16'b0000000000000000;
	sram_mem[113307] = 16'b0000000000000000;
	sram_mem[113308] = 16'b0000000000000000;
	sram_mem[113309] = 16'b0000000000000000;
	sram_mem[113310] = 16'b0000000000000000;
	sram_mem[113311] = 16'b0000000000000000;
	sram_mem[113312] = 16'b0000000000000000;
	sram_mem[113313] = 16'b0000000000000000;
	sram_mem[113314] = 16'b0000000000000000;
	sram_mem[113315] = 16'b0000000000000000;
	sram_mem[113316] = 16'b0000000000000000;
	sram_mem[113317] = 16'b0000000000000000;
	sram_mem[113318] = 16'b0000000000000000;
	sram_mem[113319] = 16'b0000000000000000;
	sram_mem[113320] = 16'b0000000000000000;
	sram_mem[113321] = 16'b0000000000000000;
	sram_mem[113322] = 16'b0000000000000000;
	sram_mem[113323] = 16'b0000000000000000;
	sram_mem[113324] = 16'b0000000000000000;
	sram_mem[113325] = 16'b0000000000000000;
	sram_mem[113326] = 16'b0000000000000000;
	sram_mem[113327] = 16'b0000000000000000;
	sram_mem[113328] = 16'b0000000000000000;
	sram_mem[113329] = 16'b0000000000000000;
	sram_mem[113330] = 16'b0000000000000000;
	sram_mem[113331] = 16'b0000000000000000;
	sram_mem[113332] = 16'b0000000000000000;
	sram_mem[113333] = 16'b0000000000000000;
	sram_mem[113334] = 16'b0000000000000000;
	sram_mem[113335] = 16'b0000000000000000;
	sram_mem[113336] = 16'b0000000000000000;
	sram_mem[113337] = 16'b0000000000000000;
	sram_mem[113338] = 16'b0000000000000000;
	sram_mem[113339] = 16'b0000000000000000;
	sram_mem[113340] = 16'b0000000000000000;
	sram_mem[113341] = 16'b0000000000000000;
	sram_mem[113342] = 16'b0000000000000000;
	sram_mem[113343] = 16'b0000000000000000;
	sram_mem[113344] = 16'b0000000000000000;
	sram_mem[113345] = 16'b0000000000000000;
	sram_mem[113346] = 16'b0000000000000000;
	sram_mem[113347] = 16'b0000000000000000;
	sram_mem[113348] = 16'b0000000000000000;
	sram_mem[113349] = 16'b0000000000000000;
	sram_mem[113350] = 16'b0000000000000000;
	sram_mem[113351] = 16'b0000000000000000;
	sram_mem[113352] = 16'b0000000000000000;
	sram_mem[113353] = 16'b0000000000000000;
	sram_mem[113354] = 16'b0000000000000000;
	sram_mem[113355] = 16'b0000000000000000;
	sram_mem[113356] = 16'b0000000000000000;
	sram_mem[113357] = 16'b0000000000000000;
	sram_mem[113358] = 16'b0000000000000000;
	sram_mem[113359] = 16'b0000000000000000;
	sram_mem[113360] = 16'b0000000000000000;
	sram_mem[113361] = 16'b0000000000000000;
	sram_mem[113362] = 16'b0000000000000000;
	sram_mem[113363] = 16'b0000000000000000;
	sram_mem[113364] = 16'b0000000000000000;
	sram_mem[113365] = 16'b0000000000000000;
	sram_mem[113366] = 16'b0000000000000000;
	sram_mem[113367] = 16'b0000000000000000;
	sram_mem[113368] = 16'b0000000000000000;
	sram_mem[113369] = 16'b0000000000000000;
	sram_mem[113370] = 16'b0000000000000000;
	sram_mem[113371] = 16'b0000000000000000;
	sram_mem[113372] = 16'b0000000000000000;
	sram_mem[113373] = 16'b0000000000000000;
	sram_mem[113374] = 16'b0000000000000000;
	sram_mem[113375] = 16'b0000000000000000;
	sram_mem[113376] = 16'b0000000000000000;
	sram_mem[113377] = 16'b0000000000000000;
	sram_mem[113378] = 16'b0000000000000000;
	sram_mem[113379] = 16'b0000000000000000;
	sram_mem[113380] = 16'b0000000000000000;
	sram_mem[113381] = 16'b0000000000000000;
	sram_mem[113382] = 16'b0000000000000000;
	sram_mem[113383] = 16'b0000000000000000;
	sram_mem[113384] = 16'b0000000000000000;
	sram_mem[113385] = 16'b0000000000000000;
	sram_mem[113386] = 16'b0000000000000000;
	sram_mem[113387] = 16'b0000000000000000;
	sram_mem[113388] = 16'b0000000000000000;
	sram_mem[113389] = 16'b0000000000000000;
	sram_mem[113390] = 16'b0000000000000000;
	sram_mem[113391] = 16'b0000000000000000;
	sram_mem[113392] = 16'b0000000000000000;
	sram_mem[113393] = 16'b0000000000000000;
	sram_mem[113394] = 16'b0000000000000000;
	sram_mem[113395] = 16'b0000000000000000;
	sram_mem[113396] = 16'b0000000000000000;
	sram_mem[113397] = 16'b0000000000000000;
	sram_mem[113398] = 16'b0000000000000000;
	sram_mem[113399] = 16'b0000000000000000;
	sram_mem[113400] = 16'b0000000000000000;
	sram_mem[113401] = 16'b0000000000000000;
	sram_mem[113402] = 16'b0000000000000000;
	sram_mem[113403] = 16'b0000000000000000;
	sram_mem[113404] = 16'b0000000000000000;
	sram_mem[113405] = 16'b0000000000000000;
	sram_mem[113406] = 16'b0000000000000000;
	sram_mem[113407] = 16'b0000000000000000;
	sram_mem[113408] = 16'b0000000000000000;
	sram_mem[113409] = 16'b0000000000000000;
	sram_mem[113410] = 16'b0000000000000000;
	sram_mem[113411] = 16'b0000000000000000;
	sram_mem[113412] = 16'b0000000000000000;
	sram_mem[113413] = 16'b0000000000000000;
	sram_mem[113414] = 16'b0000000000000000;
	sram_mem[113415] = 16'b0000000000000000;
	sram_mem[113416] = 16'b0000000000000000;
	sram_mem[113417] = 16'b0000000000000000;
	sram_mem[113418] = 16'b0000000000000000;
	sram_mem[113419] = 16'b0000000000000000;
	sram_mem[113420] = 16'b0000000000000000;
	sram_mem[113421] = 16'b0000000000000000;
	sram_mem[113422] = 16'b0000000000000000;
	sram_mem[113423] = 16'b0000000000000000;
	sram_mem[113424] = 16'b0000000000000000;
	sram_mem[113425] = 16'b0000000000000000;
	sram_mem[113426] = 16'b0000000000000000;
	sram_mem[113427] = 16'b0000000000000000;
	sram_mem[113428] = 16'b0000000000000000;
	sram_mem[113429] = 16'b0000000000000000;
	sram_mem[113430] = 16'b0000000000000000;
	sram_mem[113431] = 16'b0000000000000000;
	sram_mem[113432] = 16'b0000000000000000;
	sram_mem[113433] = 16'b0000000000000000;
	sram_mem[113434] = 16'b0000000000000000;
	sram_mem[113435] = 16'b0000000000000000;
	sram_mem[113436] = 16'b0000000000000000;
	sram_mem[113437] = 16'b0000000000000000;
	sram_mem[113438] = 16'b0000000000000000;
	sram_mem[113439] = 16'b0000000000000000;
	sram_mem[113440] = 16'b0000000000000000;
	sram_mem[113441] = 16'b0000000000000000;
	sram_mem[113442] = 16'b0000000000000000;
	sram_mem[113443] = 16'b0000000000000000;
	sram_mem[113444] = 16'b0000000000000000;
	sram_mem[113445] = 16'b0000000000000000;
	sram_mem[113446] = 16'b0000000000000000;
	sram_mem[113447] = 16'b0000000000000000;
	sram_mem[113448] = 16'b0000000000000000;
	sram_mem[113449] = 16'b0000000000000000;
	sram_mem[113450] = 16'b0000000000000000;
	sram_mem[113451] = 16'b0000000000000000;
	sram_mem[113452] = 16'b0000000000000000;
	sram_mem[113453] = 16'b0000000000000000;
	sram_mem[113454] = 16'b0000000000000000;
	sram_mem[113455] = 16'b0000000000000000;
	sram_mem[113456] = 16'b0000000000000000;
	sram_mem[113457] = 16'b0000000000000000;
	sram_mem[113458] = 16'b0000000000000000;
	sram_mem[113459] = 16'b0000000000000000;
	sram_mem[113460] = 16'b0000000000000000;
	sram_mem[113461] = 16'b0000000000000000;
	sram_mem[113462] = 16'b0000000000000000;
	sram_mem[113463] = 16'b0000000000000000;
	sram_mem[113464] = 16'b0000000000000000;
	sram_mem[113465] = 16'b0000000000000000;
	sram_mem[113466] = 16'b0000000000000000;
	sram_mem[113467] = 16'b0000000000000000;
	sram_mem[113468] = 16'b0000000000000000;
	sram_mem[113469] = 16'b0000000000000000;
	sram_mem[113470] = 16'b0000000000000000;
	sram_mem[113471] = 16'b0000000000000000;
	sram_mem[113472] = 16'b0000000000000000;
	sram_mem[113473] = 16'b0000000000000000;
	sram_mem[113474] = 16'b0000000000000000;
	sram_mem[113475] = 16'b0000000000000000;
	sram_mem[113476] = 16'b0000000000000000;
	sram_mem[113477] = 16'b0000000000000000;
	sram_mem[113478] = 16'b0000000000000000;
	sram_mem[113479] = 16'b0000000000000000;
	sram_mem[113480] = 16'b0000000000000000;
	sram_mem[113481] = 16'b0000000000000000;
	sram_mem[113482] = 16'b0000000000000000;
	sram_mem[113483] = 16'b0000000000000000;
	sram_mem[113484] = 16'b0000000000000000;
	sram_mem[113485] = 16'b0000000000000000;
	sram_mem[113486] = 16'b0000000000000000;
	sram_mem[113487] = 16'b0000000000000000;
	sram_mem[113488] = 16'b0000000000000000;
	sram_mem[113489] = 16'b0000000000000000;
	sram_mem[113490] = 16'b0000000000000000;
	sram_mem[113491] = 16'b0000000000000000;
	sram_mem[113492] = 16'b0000000000000000;
	sram_mem[113493] = 16'b0000000000000000;
	sram_mem[113494] = 16'b0000000000000000;
	sram_mem[113495] = 16'b0000000000000000;
	sram_mem[113496] = 16'b0000000000000000;
	sram_mem[113497] = 16'b0000000000000000;
	sram_mem[113498] = 16'b0000000000000000;
	sram_mem[113499] = 16'b0000000000000000;
	sram_mem[113500] = 16'b0000000000000000;
	sram_mem[113501] = 16'b0000000000000000;
	sram_mem[113502] = 16'b0000000000000000;
	sram_mem[113503] = 16'b0000000000000000;
	sram_mem[113504] = 16'b0000000000000000;
	sram_mem[113505] = 16'b0000000000000000;
	sram_mem[113506] = 16'b0000000000000000;
	sram_mem[113507] = 16'b0000000000000000;
	sram_mem[113508] = 16'b0000000000000000;
	sram_mem[113509] = 16'b0000000000000000;
	sram_mem[113510] = 16'b0000000000000000;
	sram_mem[113511] = 16'b0000000000000000;
	sram_mem[113512] = 16'b0000000000000000;
	sram_mem[113513] = 16'b0000000000000000;
	sram_mem[113514] = 16'b0000000000000000;
	sram_mem[113515] = 16'b0000000000000000;
	sram_mem[113516] = 16'b0000000000000000;
	sram_mem[113517] = 16'b0000000000000000;
	sram_mem[113518] = 16'b0000000000000000;
	sram_mem[113519] = 16'b0000000000000000;
	sram_mem[113520] = 16'b0000000000000000;
	sram_mem[113521] = 16'b0000000000000000;
	sram_mem[113522] = 16'b0000000000000000;
	sram_mem[113523] = 16'b0000000000000000;
	sram_mem[113524] = 16'b0000000000000000;
	sram_mem[113525] = 16'b0000000000000000;
	sram_mem[113526] = 16'b0000000000000000;
	sram_mem[113527] = 16'b0000000000000000;
	sram_mem[113528] = 16'b0000000000000000;
	sram_mem[113529] = 16'b0000000000000000;
	sram_mem[113530] = 16'b0000000000000000;
	sram_mem[113531] = 16'b0000000000000000;
	sram_mem[113532] = 16'b0000000000000000;
	sram_mem[113533] = 16'b0000000000000000;
	sram_mem[113534] = 16'b0000000000000000;
	sram_mem[113535] = 16'b0000000000000000;
	sram_mem[113536] = 16'b0000000000000000;
	sram_mem[113537] = 16'b0000000000000000;
	sram_mem[113538] = 16'b0000000000000000;
	sram_mem[113539] = 16'b0000000000000000;
	sram_mem[113540] = 16'b0000000000000000;
	sram_mem[113541] = 16'b0000000000000000;
	sram_mem[113542] = 16'b0000000000000000;
	sram_mem[113543] = 16'b0000000000000000;
	sram_mem[113544] = 16'b0000000000000000;
	sram_mem[113545] = 16'b0000000000000000;
	sram_mem[113546] = 16'b0000000000000000;
	sram_mem[113547] = 16'b0000000000000000;
	sram_mem[113548] = 16'b0000000000000000;
	sram_mem[113549] = 16'b0000000000000000;
	sram_mem[113550] = 16'b0000000000000000;
	sram_mem[113551] = 16'b0000000000000000;
	sram_mem[113552] = 16'b0000000000000000;
	sram_mem[113553] = 16'b0000000000000000;
	sram_mem[113554] = 16'b0000000000000000;
	sram_mem[113555] = 16'b0000000000000000;
	sram_mem[113556] = 16'b0000000000000000;
	sram_mem[113557] = 16'b0000000000000000;
	sram_mem[113558] = 16'b0000000000000000;
	sram_mem[113559] = 16'b0000000000000000;
	sram_mem[113560] = 16'b0000000000000000;
	sram_mem[113561] = 16'b0000000000000000;
	sram_mem[113562] = 16'b0000000000000000;
	sram_mem[113563] = 16'b0000000000000000;
	sram_mem[113564] = 16'b0000000000000000;
	sram_mem[113565] = 16'b0000000000000000;
	sram_mem[113566] = 16'b0000000000000000;
	sram_mem[113567] = 16'b0000000000000000;
	sram_mem[113568] = 16'b0000000000000000;
	sram_mem[113569] = 16'b0000000000000000;
	sram_mem[113570] = 16'b0000000000000000;
	sram_mem[113571] = 16'b0000000000000000;
	sram_mem[113572] = 16'b0000000000000000;
	sram_mem[113573] = 16'b0000000000000000;
	sram_mem[113574] = 16'b0000000000000000;
	sram_mem[113575] = 16'b0000000000000000;
	sram_mem[113576] = 16'b0000000000000000;
	sram_mem[113577] = 16'b0000000000000000;
	sram_mem[113578] = 16'b0000000000000000;
	sram_mem[113579] = 16'b0000000000000000;
	sram_mem[113580] = 16'b0000000000000000;
	sram_mem[113581] = 16'b0000000000000000;
	sram_mem[113582] = 16'b0000000000000000;
	sram_mem[113583] = 16'b0000000000000000;
	sram_mem[113584] = 16'b0000000000000000;
	sram_mem[113585] = 16'b0000000000000000;
	sram_mem[113586] = 16'b0000000000000000;
	sram_mem[113587] = 16'b0000000000000000;
	sram_mem[113588] = 16'b0000000000000000;
	sram_mem[113589] = 16'b0000000000000000;
	sram_mem[113590] = 16'b0000000000000000;
	sram_mem[113591] = 16'b0000000000000000;
	sram_mem[113592] = 16'b0000000000000000;
	sram_mem[113593] = 16'b0000000000000000;
	sram_mem[113594] = 16'b0000000000000000;
	sram_mem[113595] = 16'b0000000000000000;
	sram_mem[113596] = 16'b0000000000000000;
	sram_mem[113597] = 16'b0000000000000000;
	sram_mem[113598] = 16'b0000000000000000;
	sram_mem[113599] = 16'b0000000000000000;
	sram_mem[113600] = 16'b0000000000000000;
	sram_mem[113601] = 16'b0000000000000000;
	sram_mem[113602] = 16'b0000000000000000;
	sram_mem[113603] = 16'b0000000000000000;
	sram_mem[113604] = 16'b0000000000000000;
	sram_mem[113605] = 16'b0000000000000000;
	sram_mem[113606] = 16'b0000000000000000;
	sram_mem[113607] = 16'b0000000000000000;
	sram_mem[113608] = 16'b0000000000000000;
	sram_mem[113609] = 16'b0000000000000000;
	sram_mem[113610] = 16'b0000000000000000;
	sram_mem[113611] = 16'b0000000000000000;
	sram_mem[113612] = 16'b0000000000000000;
	sram_mem[113613] = 16'b0000000000000000;
	sram_mem[113614] = 16'b0000000000000000;
	sram_mem[113615] = 16'b0000000000000000;
	sram_mem[113616] = 16'b0000000000000000;
	sram_mem[113617] = 16'b0000000000000000;
	sram_mem[113618] = 16'b0000000000000000;
	sram_mem[113619] = 16'b0000000000000000;
	sram_mem[113620] = 16'b0000000000000000;
	sram_mem[113621] = 16'b0000000000000000;
	sram_mem[113622] = 16'b0000000000000000;
	sram_mem[113623] = 16'b0000000000000000;
	sram_mem[113624] = 16'b0000000000000000;
	sram_mem[113625] = 16'b0000000000000000;
	sram_mem[113626] = 16'b0000000000000000;
	sram_mem[113627] = 16'b0000000000000000;
	sram_mem[113628] = 16'b0000000000000000;
	sram_mem[113629] = 16'b0000000000000000;
	sram_mem[113630] = 16'b0000000000000000;
	sram_mem[113631] = 16'b0000000000000000;
	sram_mem[113632] = 16'b0000000000000000;
	sram_mem[113633] = 16'b0000000000000000;
	sram_mem[113634] = 16'b0000000000000000;
	sram_mem[113635] = 16'b0000000000000000;
	sram_mem[113636] = 16'b0000000000000000;
	sram_mem[113637] = 16'b0000000000000000;
	sram_mem[113638] = 16'b0000000000000000;
	sram_mem[113639] = 16'b0000000000000000;
	sram_mem[113640] = 16'b0000000000000000;
	sram_mem[113641] = 16'b0000000000000000;
	sram_mem[113642] = 16'b0000000000000000;
	sram_mem[113643] = 16'b0000000000000000;
	sram_mem[113644] = 16'b0000000000000000;
	sram_mem[113645] = 16'b0000000000000000;
	sram_mem[113646] = 16'b0000000000000000;
	sram_mem[113647] = 16'b0000000000000000;
	sram_mem[113648] = 16'b0000000000000000;
	sram_mem[113649] = 16'b0000000000000000;
	sram_mem[113650] = 16'b0000000000000000;
	sram_mem[113651] = 16'b0000000000000000;
	sram_mem[113652] = 16'b0000000000000000;
	sram_mem[113653] = 16'b0000000000000000;
	sram_mem[113654] = 16'b0000000000000000;
	sram_mem[113655] = 16'b0000000000000000;
	sram_mem[113656] = 16'b0000000000000000;
	sram_mem[113657] = 16'b0000000000000000;
	sram_mem[113658] = 16'b0000000000000000;
	sram_mem[113659] = 16'b0000000000000000;
	sram_mem[113660] = 16'b0000000000000000;
	sram_mem[113661] = 16'b0000000000000000;
	sram_mem[113662] = 16'b0000000000000000;
	sram_mem[113663] = 16'b0000000000000000;
	sram_mem[113664] = 16'b0000000000000000;
	sram_mem[113665] = 16'b0000000000000000;
	sram_mem[113666] = 16'b0000000000000000;
	sram_mem[113667] = 16'b0000000000000000;
	sram_mem[113668] = 16'b0000000000000000;
	sram_mem[113669] = 16'b0000000000000000;
	sram_mem[113670] = 16'b0000000000000000;
	sram_mem[113671] = 16'b0000000000000000;
	sram_mem[113672] = 16'b0000000000000000;
	sram_mem[113673] = 16'b0000000000000000;
	sram_mem[113674] = 16'b0000000000000000;
	sram_mem[113675] = 16'b0000000000000000;
	sram_mem[113676] = 16'b0000000000000000;
	sram_mem[113677] = 16'b0000000000000000;
	sram_mem[113678] = 16'b0000000000000000;
	sram_mem[113679] = 16'b0000000000000000;
	sram_mem[113680] = 16'b0000000000000000;
	sram_mem[113681] = 16'b0000000000000000;
	sram_mem[113682] = 16'b0000000000000000;
	sram_mem[113683] = 16'b0000000000000000;
	sram_mem[113684] = 16'b0000000000000000;
	sram_mem[113685] = 16'b0000000000000000;
	sram_mem[113686] = 16'b0000000000000000;
	sram_mem[113687] = 16'b0000000000000000;
	sram_mem[113688] = 16'b0000000000000000;
	sram_mem[113689] = 16'b0000000000000000;
	sram_mem[113690] = 16'b0000000000000000;
	sram_mem[113691] = 16'b0000000000000000;
	sram_mem[113692] = 16'b0000000000000000;
	sram_mem[113693] = 16'b0000000000000000;
	sram_mem[113694] = 16'b0000000000000000;
	sram_mem[113695] = 16'b0000000000000000;
	sram_mem[113696] = 16'b0000000000000000;
	sram_mem[113697] = 16'b0000000000000000;
	sram_mem[113698] = 16'b0000000000000000;
	sram_mem[113699] = 16'b0000000000000000;
	sram_mem[113700] = 16'b0000000000000000;
	sram_mem[113701] = 16'b0000000000000000;
	sram_mem[113702] = 16'b0000000000000000;
	sram_mem[113703] = 16'b0000000000000000;
	sram_mem[113704] = 16'b0000000000000000;
	sram_mem[113705] = 16'b0000000000000000;
	sram_mem[113706] = 16'b0000000000000000;
	sram_mem[113707] = 16'b0000000000000000;
	sram_mem[113708] = 16'b0000000000000000;
	sram_mem[113709] = 16'b0000000000000000;
	sram_mem[113710] = 16'b0000000000000000;
	sram_mem[113711] = 16'b0000000000000000;
	sram_mem[113712] = 16'b0000000000000000;
	sram_mem[113713] = 16'b0000000000000000;
	sram_mem[113714] = 16'b0000000000000000;
	sram_mem[113715] = 16'b0000000000000000;
	sram_mem[113716] = 16'b0000000000000000;
	sram_mem[113717] = 16'b0000000000000000;
	sram_mem[113718] = 16'b0000000000000000;
	sram_mem[113719] = 16'b0000000000000000;
	sram_mem[113720] = 16'b0000000000000000;
	sram_mem[113721] = 16'b0000000000000000;
	sram_mem[113722] = 16'b0000000000000000;
	sram_mem[113723] = 16'b0000000000000000;
	sram_mem[113724] = 16'b0000000000000000;
	sram_mem[113725] = 16'b0000000000000000;
	sram_mem[113726] = 16'b0000000000000000;
	sram_mem[113727] = 16'b0000000000000000;
	sram_mem[113728] = 16'b0000000000000000;
	sram_mem[113729] = 16'b0000000000000000;
	sram_mem[113730] = 16'b0000000000000000;
	sram_mem[113731] = 16'b0000000000000000;
	sram_mem[113732] = 16'b0000000000000000;
	sram_mem[113733] = 16'b0000000000000000;
	sram_mem[113734] = 16'b0000000000000000;
	sram_mem[113735] = 16'b0000000000000000;
	sram_mem[113736] = 16'b0000000000000000;
	sram_mem[113737] = 16'b0000000000000000;
	sram_mem[113738] = 16'b0000000000000000;
	sram_mem[113739] = 16'b0000000000000000;
	sram_mem[113740] = 16'b0000000000000000;
	sram_mem[113741] = 16'b0000000000000000;
	sram_mem[113742] = 16'b0000000000000000;
	sram_mem[113743] = 16'b0000000000000000;
	sram_mem[113744] = 16'b0000000000000000;
	sram_mem[113745] = 16'b0000000000000000;
	sram_mem[113746] = 16'b0000000000000000;
	sram_mem[113747] = 16'b0000000000000000;
	sram_mem[113748] = 16'b0000000000000000;
	sram_mem[113749] = 16'b0000000000000000;
	sram_mem[113750] = 16'b0000000000000000;
	sram_mem[113751] = 16'b0000000000000000;
	sram_mem[113752] = 16'b0000000000000000;
	sram_mem[113753] = 16'b0000000000000000;
	sram_mem[113754] = 16'b0000000000000000;
	sram_mem[113755] = 16'b0000000000000000;
	sram_mem[113756] = 16'b0000000000000000;
	sram_mem[113757] = 16'b0000000000000000;
	sram_mem[113758] = 16'b0000000000000000;
	sram_mem[113759] = 16'b0000000000000000;
	sram_mem[113760] = 16'b0000000000000000;
	sram_mem[113761] = 16'b0000000000000000;
	sram_mem[113762] = 16'b0000000000000000;
	sram_mem[113763] = 16'b0000000000000000;
	sram_mem[113764] = 16'b0000000000000000;
	sram_mem[113765] = 16'b0000000000000000;
	sram_mem[113766] = 16'b0000000000000000;
	sram_mem[113767] = 16'b0000000000000000;
	sram_mem[113768] = 16'b0000000000000000;
	sram_mem[113769] = 16'b0000000000000000;
	sram_mem[113770] = 16'b0000000000000000;
	sram_mem[113771] = 16'b0000000000000000;
	sram_mem[113772] = 16'b0000000000000000;
	sram_mem[113773] = 16'b0000000000000000;
	sram_mem[113774] = 16'b0000000000000000;
	sram_mem[113775] = 16'b0000000000000000;
	sram_mem[113776] = 16'b0000000000000000;
	sram_mem[113777] = 16'b0000000000000000;
	sram_mem[113778] = 16'b0000000000000000;
	sram_mem[113779] = 16'b0000000000000000;
	sram_mem[113780] = 16'b0000000000000000;
	sram_mem[113781] = 16'b0000000000000000;
	sram_mem[113782] = 16'b0000000000000000;
	sram_mem[113783] = 16'b0000000000000000;
	sram_mem[113784] = 16'b0000000000000000;
	sram_mem[113785] = 16'b0000000000000000;
	sram_mem[113786] = 16'b0000000000000000;
	sram_mem[113787] = 16'b0000000000000000;
	sram_mem[113788] = 16'b0000000000000000;
	sram_mem[113789] = 16'b0000000000000000;
	sram_mem[113790] = 16'b0000000000000000;
	sram_mem[113791] = 16'b0000000000000000;
	sram_mem[113792] = 16'b0000000000000000;
	sram_mem[113793] = 16'b0000000000000000;
	sram_mem[113794] = 16'b0000000000000000;
	sram_mem[113795] = 16'b0000000000000000;
	sram_mem[113796] = 16'b0000000000000000;
	sram_mem[113797] = 16'b0000000000000000;
	sram_mem[113798] = 16'b0000000000000000;
	sram_mem[113799] = 16'b0000000000000000;
	sram_mem[113800] = 16'b0000000000000000;
	sram_mem[113801] = 16'b0000000000000000;
	sram_mem[113802] = 16'b0000000000000000;
	sram_mem[113803] = 16'b0000000000000000;
	sram_mem[113804] = 16'b0000000000000000;
	sram_mem[113805] = 16'b0000000000000000;
	sram_mem[113806] = 16'b0000000000000000;
	sram_mem[113807] = 16'b0000000000000000;
	sram_mem[113808] = 16'b0000000000000000;
	sram_mem[113809] = 16'b0000000000000000;
	sram_mem[113810] = 16'b0000000000000000;
	sram_mem[113811] = 16'b0000000000000000;
	sram_mem[113812] = 16'b0000000000000000;
	sram_mem[113813] = 16'b0000000000000000;
	sram_mem[113814] = 16'b0000000000000000;
	sram_mem[113815] = 16'b0000000000000000;
	sram_mem[113816] = 16'b0000000000000000;
	sram_mem[113817] = 16'b0000000000000000;
	sram_mem[113818] = 16'b0000000000000000;
	sram_mem[113819] = 16'b0000000000000000;
	sram_mem[113820] = 16'b0000000000000000;
	sram_mem[113821] = 16'b0000000000000000;
	sram_mem[113822] = 16'b0000000000000000;
	sram_mem[113823] = 16'b0000000000000000;
	sram_mem[113824] = 16'b0000000000000000;
	sram_mem[113825] = 16'b0000000000000000;
	sram_mem[113826] = 16'b0000000000000000;
	sram_mem[113827] = 16'b0000000000000000;
	sram_mem[113828] = 16'b0000000000000000;
	sram_mem[113829] = 16'b0000000000000000;
	sram_mem[113830] = 16'b0000000000000000;
	sram_mem[113831] = 16'b0000000000000000;
	sram_mem[113832] = 16'b0000000000000000;
	sram_mem[113833] = 16'b0000000000000000;
	sram_mem[113834] = 16'b0000000000000000;
	sram_mem[113835] = 16'b0000000000000000;
	sram_mem[113836] = 16'b0000000000000000;
	sram_mem[113837] = 16'b0000000000000000;
	sram_mem[113838] = 16'b0000000000000000;
	sram_mem[113839] = 16'b0000000000000000;
	sram_mem[113840] = 16'b0000000000000000;
	sram_mem[113841] = 16'b0000000000000000;
	sram_mem[113842] = 16'b0000000000000000;
	sram_mem[113843] = 16'b0000000000000000;
	sram_mem[113844] = 16'b0000000000000000;
	sram_mem[113845] = 16'b0000000000000000;
	sram_mem[113846] = 16'b0000000000000000;
	sram_mem[113847] = 16'b0000000000000000;
	sram_mem[113848] = 16'b0000000000000000;
	sram_mem[113849] = 16'b0000000000000000;
	sram_mem[113850] = 16'b0000000000000000;
	sram_mem[113851] = 16'b0000000000000000;
	sram_mem[113852] = 16'b0000000000000000;
	sram_mem[113853] = 16'b0000000000000000;
	sram_mem[113854] = 16'b0000000000000000;
	sram_mem[113855] = 16'b0000000000000000;
	sram_mem[113856] = 16'b0000000000000000;
	sram_mem[113857] = 16'b0000000000000000;
	sram_mem[113858] = 16'b0000000000000000;
	sram_mem[113859] = 16'b0000000000000000;
	sram_mem[113860] = 16'b0000000000000000;
	sram_mem[113861] = 16'b0000000000000000;
	sram_mem[113862] = 16'b0000000000000000;
	sram_mem[113863] = 16'b0000000000000000;
	sram_mem[113864] = 16'b0000000000000000;
	sram_mem[113865] = 16'b0000000000000000;
	sram_mem[113866] = 16'b0000000000000000;
	sram_mem[113867] = 16'b0000000000000000;
	sram_mem[113868] = 16'b0000000000000000;
	sram_mem[113869] = 16'b0000000000000000;
	sram_mem[113870] = 16'b0000000000000000;
	sram_mem[113871] = 16'b0000000000000000;
	sram_mem[113872] = 16'b0000000000000000;
	sram_mem[113873] = 16'b0000000000000000;
	sram_mem[113874] = 16'b0000000000000000;
	sram_mem[113875] = 16'b0000000000000000;
	sram_mem[113876] = 16'b0000000000000000;
	sram_mem[113877] = 16'b0000000000000000;
	sram_mem[113878] = 16'b0000000000000000;
	sram_mem[113879] = 16'b0000000000000000;
	sram_mem[113880] = 16'b0000000000000000;
	sram_mem[113881] = 16'b0000000000000000;
	sram_mem[113882] = 16'b0000000000000000;
	sram_mem[113883] = 16'b0000000000000000;
	sram_mem[113884] = 16'b0000000000000000;
	sram_mem[113885] = 16'b0000000000000000;
	sram_mem[113886] = 16'b0000000000000000;
	sram_mem[113887] = 16'b0000000000000000;
	sram_mem[113888] = 16'b0000000000000000;
	sram_mem[113889] = 16'b0000000000000000;
	sram_mem[113890] = 16'b0000000000000000;
	sram_mem[113891] = 16'b0000000000000000;
	sram_mem[113892] = 16'b0000000000000000;
	sram_mem[113893] = 16'b0000000000000000;
	sram_mem[113894] = 16'b0000000000000000;
	sram_mem[113895] = 16'b0000000000000000;
	sram_mem[113896] = 16'b0000000000000000;
	sram_mem[113897] = 16'b0000000000000000;
	sram_mem[113898] = 16'b0000000000000000;
	sram_mem[113899] = 16'b0000000000000000;
	sram_mem[113900] = 16'b0000000000000000;
	sram_mem[113901] = 16'b0000000000000000;
	sram_mem[113902] = 16'b0000000000000000;
	sram_mem[113903] = 16'b0000000000000000;
	sram_mem[113904] = 16'b0000000000000000;
	sram_mem[113905] = 16'b0000000000000000;
	sram_mem[113906] = 16'b0000000000000000;
	sram_mem[113907] = 16'b0000000000000000;
	sram_mem[113908] = 16'b0000000000000000;
	sram_mem[113909] = 16'b0000000000000000;
	sram_mem[113910] = 16'b0000000000000000;
	sram_mem[113911] = 16'b0000000000000000;
	sram_mem[113912] = 16'b0000000000000000;
	sram_mem[113913] = 16'b0000000000000000;
	sram_mem[113914] = 16'b0000000000000000;
	sram_mem[113915] = 16'b0000000000000000;
	sram_mem[113916] = 16'b0000000000000000;
	sram_mem[113917] = 16'b0000000000000000;
	sram_mem[113918] = 16'b0000000000000000;
	sram_mem[113919] = 16'b0000000000000000;
	sram_mem[113920] = 16'b0000000000000000;
	sram_mem[113921] = 16'b0000000000000000;
	sram_mem[113922] = 16'b0000000000000000;
	sram_mem[113923] = 16'b0000000000000000;
	sram_mem[113924] = 16'b0000000000000000;
	sram_mem[113925] = 16'b0000000000000000;
	sram_mem[113926] = 16'b0000000000000000;
	sram_mem[113927] = 16'b0000000000000000;
	sram_mem[113928] = 16'b0000000000000000;
	sram_mem[113929] = 16'b0000000000000000;
	sram_mem[113930] = 16'b0000000000000000;
	sram_mem[113931] = 16'b0000000000000000;
	sram_mem[113932] = 16'b0000000000000000;
	sram_mem[113933] = 16'b0000000000000000;
	sram_mem[113934] = 16'b0000000000000000;
	sram_mem[113935] = 16'b0000000000000000;
	sram_mem[113936] = 16'b0000000000000000;
	sram_mem[113937] = 16'b0000000000000000;
	sram_mem[113938] = 16'b0000000000000000;
	sram_mem[113939] = 16'b0000000000000000;
	sram_mem[113940] = 16'b0000000000000000;
	sram_mem[113941] = 16'b0000000000000000;
	sram_mem[113942] = 16'b0000000000000000;
	sram_mem[113943] = 16'b0000000000000000;
	sram_mem[113944] = 16'b0000000000000000;
	sram_mem[113945] = 16'b0000000000000000;
	sram_mem[113946] = 16'b0000000000000000;
	sram_mem[113947] = 16'b0000000000000000;
	sram_mem[113948] = 16'b0000000000000000;
	sram_mem[113949] = 16'b0000000000000000;
	sram_mem[113950] = 16'b0000000000000000;
	sram_mem[113951] = 16'b0000000000000000;
	sram_mem[113952] = 16'b0000000000000000;
	sram_mem[113953] = 16'b0000000000000000;
	sram_mem[113954] = 16'b0000000000000000;
	sram_mem[113955] = 16'b0000000000000000;
	sram_mem[113956] = 16'b0000000000000000;
	sram_mem[113957] = 16'b0000000000000000;
	sram_mem[113958] = 16'b0000000000000000;
	sram_mem[113959] = 16'b0000000000000000;
	sram_mem[113960] = 16'b0000000000000000;
	sram_mem[113961] = 16'b0000000000000000;
	sram_mem[113962] = 16'b0000000000000000;
	sram_mem[113963] = 16'b0000000000000000;
	sram_mem[113964] = 16'b0000000000000000;
	sram_mem[113965] = 16'b0000000000000000;
	sram_mem[113966] = 16'b0000000000000000;
	sram_mem[113967] = 16'b0000000000000000;
	sram_mem[113968] = 16'b0000000000000000;
	sram_mem[113969] = 16'b0000000000000000;
	sram_mem[113970] = 16'b0000000000000000;
	sram_mem[113971] = 16'b0000000000000000;
	sram_mem[113972] = 16'b0000000000000000;
	sram_mem[113973] = 16'b0000000000000000;
	sram_mem[113974] = 16'b0000000000000000;
	sram_mem[113975] = 16'b0000000000000000;
	sram_mem[113976] = 16'b0000000000000000;
	sram_mem[113977] = 16'b0000000000000000;
	sram_mem[113978] = 16'b0000000000000000;
	sram_mem[113979] = 16'b0000000000000000;
	sram_mem[113980] = 16'b0000000000000000;
	sram_mem[113981] = 16'b0000000000000000;
	sram_mem[113982] = 16'b0000000000000000;
	sram_mem[113983] = 16'b0000000000000000;
	sram_mem[113984] = 16'b0000000000000000;
	sram_mem[113985] = 16'b0000000000000000;
	sram_mem[113986] = 16'b0000000000000000;
	sram_mem[113987] = 16'b0000000000000000;
	sram_mem[113988] = 16'b0000000000000000;
	sram_mem[113989] = 16'b0000000000000000;
	sram_mem[113990] = 16'b0000000000000000;
	sram_mem[113991] = 16'b0000000000000000;
	sram_mem[113992] = 16'b0000000000000000;
	sram_mem[113993] = 16'b0000000000000000;
	sram_mem[113994] = 16'b0000000000000000;
	sram_mem[113995] = 16'b0000000000000000;
	sram_mem[113996] = 16'b0000000000000000;
	sram_mem[113997] = 16'b0000000000000000;
	sram_mem[113998] = 16'b0000000000000000;
	sram_mem[113999] = 16'b0000000000000000;
	sram_mem[114000] = 16'b0000000000000000;
	sram_mem[114001] = 16'b0000000000000000;
	sram_mem[114002] = 16'b0000000000000000;
	sram_mem[114003] = 16'b0000000000000000;
	sram_mem[114004] = 16'b0000000000000000;
	sram_mem[114005] = 16'b0000000000000000;
	sram_mem[114006] = 16'b0000000000000000;
	sram_mem[114007] = 16'b0000000000000000;
	sram_mem[114008] = 16'b0000000000000000;
	sram_mem[114009] = 16'b0000000000000000;
	sram_mem[114010] = 16'b0000000000000000;
	sram_mem[114011] = 16'b0000000000000000;
	sram_mem[114012] = 16'b0000000000000000;
	sram_mem[114013] = 16'b0000000000000000;
	sram_mem[114014] = 16'b0000000000000000;
	sram_mem[114015] = 16'b0000000000000000;
	sram_mem[114016] = 16'b0000000000000000;
	sram_mem[114017] = 16'b0000000000000000;
	sram_mem[114018] = 16'b0000000000000000;
	sram_mem[114019] = 16'b0000000000000000;
	sram_mem[114020] = 16'b0000000000000000;
	sram_mem[114021] = 16'b0000000000000000;
	sram_mem[114022] = 16'b0000000000000000;
	sram_mem[114023] = 16'b0000000000000000;
	sram_mem[114024] = 16'b0000000000000000;
	sram_mem[114025] = 16'b0000000000000000;
	sram_mem[114026] = 16'b0000000000000000;
	sram_mem[114027] = 16'b0000000000000000;
	sram_mem[114028] = 16'b0000000000000000;
	sram_mem[114029] = 16'b0000000000000000;
	sram_mem[114030] = 16'b0000000000000000;
	sram_mem[114031] = 16'b0000000000000000;
	sram_mem[114032] = 16'b0000000000000000;
	sram_mem[114033] = 16'b0000000000000000;
	sram_mem[114034] = 16'b0000000000000000;
	sram_mem[114035] = 16'b0000000000000000;
	sram_mem[114036] = 16'b0000000000000000;
	sram_mem[114037] = 16'b0000000000000000;
	sram_mem[114038] = 16'b0000000000000000;
	sram_mem[114039] = 16'b0000000000000000;
	sram_mem[114040] = 16'b0000000000000000;
	sram_mem[114041] = 16'b0000000000000000;
	sram_mem[114042] = 16'b0000000000000000;
	sram_mem[114043] = 16'b0000000000000000;
	sram_mem[114044] = 16'b0000000000000000;
	sram_mem[114045] = 16'b0000000000000000;
	sram_mem[114046] = 16'b0000000000000000;
	sram_mem[114047] = 16'b0000000000000000;
	sram_mem[114048] = 16'b0000000000000000;
	sram_mem[114049] = 16'b0000000000000000;
	sram_mem[114050] = 16'b0000000000000000;
	sram_mem[114051] = 16'b0000000000000000;
	sram_mem[114052] = 16'b0000000000000000;
	sram_mem[114053] = 16'b0000000000000000;
	sram_mem[114054] = 16'b0000000000000000;
	sram_mem[114055] = 16'b0000000000000000;
	sram_mem[114056] = 16'b0000000000000000;
	sram_mem[114057] = 16'b0000000000000000;
	sram_mem[114058] = 16'b0000000000000000;
	sram_mem[114059] = 16'b0000000000000000;
	sram_mem[114060] = 16'b0000000000000000;
	sram_mem[114061] = 16'b0000000000000000;
	sram_mem[114062] = 16'b0000000000000000;
	sram_mem[114063] = 16'b0000000000000000;
	sram_mem[114064] = 16'b0000000000000000;
	sram_mem[114065] = 16'b0000000000000000;
	sram_mem[114066] = 16'b0000000000000000;
	sram_mem[114067] = 16'b0000000000000000;
	sram_mem[114068] = 16'b0000000000000000;
	sram_mem[114069] = 16'b0000000000000000;
	sram_mem[114070] = 16'b0000000000000000;
	sram_mem[114071] = 16'b0000000000000000;
	sram_mem[114072] = 16'b0000000000000000;
	sram_mem[114073] = 16'b0000000000000000;
	sram_mem[114074] = 16'b0000000000000000;
	sram_mem[114075] = 16'b0000000000000000;
	sram_mem[114076] = 16'b0000000000000000;
	sram_mem[114077] = 16'b0000000000000000;
	sram_mem[114078] = 16'b0000000000000000;
	sram_mem[114079] = 16'b0000000000000000;
	sram_mem[114080] = 16'b0000000000000000;
	sram_mem[114081] = 16'b0000000000000000;
	sram_mem[114082] = 16'b0000000000000000;
	sram_mem[114083] = 16'b0000000000000000;
	sram_mem[114084] = 16'b0000000000000000;
	sram_mem[114085] = 16'b0000000000000000;
	sram_mem[114086] = 16'b0000000000000000;
	sram_mem[114087] = 16'b0000000000000000;
	sram_mem[114088] = 16'b0000000000000000;
	sram_mem[114089] = 16'b0000000000000000;
	sram_mem[114090] = 16'b0000000000000000;
	sram_mem[114091] = 16'b0000000000000000;
	sram_mem[114092] = 16'b0000000000000000;
	sram_mem[114093] = 16'b0000000000000000;
	sram_mem[114094] = 16'b0000000000000000;
	sram_mem[114095] = 16'b0000000000000000;
	sram_mem[114096] = 16'b0000000000000000;
	sram_mem[114097] = 16'b0000000000000000;
	sram_mem[114098] = 16'b0000000000000000;
	sram_mem[114099] = 16'b0000000000000000;
	sram_mem[114100] = 16'b0000000000000000;
	sram_mem[114101] = 16'b0000000000000000;
	sram_mem[114102] = 16'b0000000000000000;
	sram_mem[114103] = 16'b0000000000000000;
	sram_mem[114104] = 16'b0000000000000000;
	sram_mem[114105] = 16'b0000000000000000;
	sram_mem[114106] = 16'b0000000000000000;
	sram_mem[114107] = 16'b0000000000000000;
	sram_mem[114108] = 16'b0000000000000000;
	sram_mem[114109] = 16'b0000000000000000;
	sram_mem[114110] = 16'b0000000000000000;
	sram_mem[114111] = 16'b0000000000000000;
	sram_mem[114112] = 16'b0000000000000000;
	sram_mem[114113] = 16'b0000000000000000;
	sram_mem[114114] = 16'b0000000000000000;
	sram_mem[114115] = 16'b0000000000000000;
	sram_mem[114116] = 16'b0000000000000000;
	sram_mem[114117] = 16'b0000000000000000;
	sram_mem[114118] = 16'b0000000000000000;
	sram_mem[114119] = 16'b0000000000000000;
	sram_mem[114120] = 16'b0000000000000000;
	sram_mem[114121] = 16'b0000000000000000;
	sram_mem[114122] = 16'b0000000000000000;
	sram_mem[114123] = 16'b0000000000000000;
	sram_mem[114124] = 16'b0000000000000000;
	sram_mem[114125] = 16'b0000000000000000;
	sram_mem[114126] = 16'b0000000000000000;
	sram_mem[114127] = 16'b0000000000000000;
	sram_mem[114128] = 16'b0000000000000000;
	sram_mem[114129] = 16'b0000000000000000;
	sram_mem[114130] = 16'b0000000000000000;
	sram_mem[114131] = 16'b0000000000000000;
	sram_mem[114132] = 16'b0000000000000000;
	sram_mem[114133] = 16'b0000000000000000;
	sram_mem[114134] = 16'b0000000000000000;
	sram_mem[114135] = 16'b0000000000000000;
	sram_mem[114136] = 16'b0000000000000000;
	sram_mem[114137] = 16'b0000000000000000;
	sram_mem[114138] = 16'b0000000000000000;
	sram_mem[114139] = 16'b0000000000000000;
	sram_mem[114140] = 16'b0000000000000000;
	sram_mem[114141] = 16'b0000000000000000;
	sram_mem[114142] = 16'b0000000000000000;
	sram_mem[114143] = 16'b0000000000000000;
	sram_mem[114144] = 16'b0000000000000000;
	sram_mem[114145] = 16'b0000000000000000;
	sram_mem[114146] = 16'b0000000000000000;
	sram_mem[114147] = 16'b0000000000000000;
	sram_mem[114148] = 16'b0000000000000000;
	sram_mem[114149] = 16'b0000000000000000;
	sram_mem[114150] = 16'b0000000000000000;
	sram_mem[114151] = 16'b0000000000000000;
	sram_mem[114152] = 16'b0000000000000000;
	sram_mem[114153] = 16'b0000000000000000;
	sram_mem[114154] = 16'b0000000000000000;
	sram_mem[114155] = 16'b0000000000000000;
	sram_mem[114156] = 16'b0000000000000000;
	sram_mem[114157] = 16'b0000000000000000;
	sram_mem[114158] = 16'b0000000000000000;
	sram_mem[114159] = 16'b0000000000000000;
	sram_mem[114160] = 16'b0000000000000000;
	sram_mem[114161] = 16'b0000000000000000;
	sram_mem[114162] = 16'b0000000000000000;
	sram_mem[114163] = 16'b0000000000000000;
	sram_mem[114164] = 16'b0000000000000000;
	sram_mem[114165] = 16'b0000000000000000;
	sram_mem[114166] = 16'b0000000000000000;
	sram_mem[114167] = 16'b0000000000000000;
	sram_mem[114168] = 16'b0000000000000000;
	sram_mem[114169] = 16'b0000000000000000;
	sram_mem[114170] = 16'b0000000000000000;
	sram_mem[114171] = 16'b0000000000000000;
	sram_mem[114172] = 16'b0000000000000000;
	sram_mem[114173] = 16'b0000000000000000;
	sram_mem[114174] = 16'b0000000000000000;
	sram_mem[114175] = 16'b0000000000000000;
	sram_mem[114176] = 16'b0000000000000000;
	sram_mem[114177] = 16'b0000000000000000;
	sram_mem[114178] = 16'b0000000000000000;
	sram_mem[114179] = 16'b0000000000000000;
	sram_mem[114180] = 16'b0000000000000000;
	sram_mem[114181] = 16'b0000000000000000;
	sram_mem[114182] = 16'b0000000000000000;
	sram_mem[114183] = 16'b0000000000000000;
	sram_mem[114184] = 16'b0000000000000000;
	sram_mem[114185] = 16'b0000000000000000;
	sram_mem[114186] = 16'b0000000000000000;
	sram_mem[114187] = 16'b0000000000000000;
	sram_mem[114188] = 16'b0000000000000000;
	sram_mem[114189] = 16'b0000000000000000;
	sram_mem[114190] = 16'b0000000000000000;
	sram_mem[114191] = 16'b0000000000000000;
	sram_mem[114192] = 16'b0000000000000000;
	sram_mem[114193] = 16'b0000000000000000;
	sram_mem[114194] = 16'b0000000000000000;
	sram_mem[114195] = 16'b0000000000000000;
	sram_mem[114196] = 16'b0000000000000000;
	sram_mem[114197] = 16'b0000000000000000;
	sram_mem[114198] = 16'b0000000000000000;
	sram_mem[114199] = 16'b0000000000000000;
	sram_mem[114200] = 16'b0000000000000000;
	sram_mem[114201] = 16'b0000000000000000;
	sram_mem[114202] = 16'b0000000000000000;
	sram_mem[114203] = 16'b0000000000000000;
	sram_mem[114204] = 16'b0000000000000000;
	sram_mem[114205] = 16'b0000000000000000;
	sram_mem[114206] = 16'b0000000000000000;
	sram_mem[114207] = 16'b0000000000000000;
	sram_mem[114208] = 16'b0000000000000000;
	sram_mem[114209] = 16'b0000000000000000;
	sram_mem[114210] = 16'b0000000000000000;
	sram_mem[114211] = 16'b0000000000000000;
	sram_mem[114212] = 16'b0000000000000000;
	sram_mem[114213] = 16'b0000000000000000;
	sram_mem[114214] = 16'b0000000000000000;
	sram_mem[114215] = 16'b0000000000000000;
	sram_mem[114216] = 16'b0000000000000000;
	sram_mem[114217] = 16'b0000000000000000;
	sram_mem[114218] = 16'b0000000000000000;
	sram_mem[114219] = 16'b0000000000000000;
	sram_mem[114220] = 16'b0000000000000000;
	sram_mem[114221] = 16'b0000000000000000;
	sram_mem[114222] = 16'b0000000000000000;
	sram_mem[114223] = 16'b0000000000000000;
	sram_mem[114224] = 16'b0000000000000000;
	sram_mem[114225] = 16'b0000000000000000;
	sram_mem[114226] = 16'b0000000000000000;
	sram_mem[114227] = 16'b0000000000000000;
	sram_mem[114228] = 16'b0000000000000000;
	sram_mem[114229] = 16'b0000000000000000;
	sram_mem[114230] = 16'b0000000000000000;
	sram_mem[114231] = 16'b0000000000000000;
	sram_mem[114232] = 16'b0000000000000000;
	sram_mem[114233] = 16'b0000000000000000;
	sram_mem[114234] = 16'b0000000000000000;
	sram_mem[114235] = 16'b0000000000000000;
	sram_mem[114236] = 16'b0000000000000000;
	sram_mem[114237] = 16'b0000000000000000;
	sram_mem[114238] = 16'b0000000000000000;
	sram_mem[114239] = 16'b0000000000000000;
	sram_mem[114240] = 16'b0000000000000000;
	sram_mem[114241] = 16'b0000000000000000;
	sram_mem[114242] = 16'b0000000000000000;
	sram_mem[114243] = 16'b0000000000000000;
	sram_mem[114244] = 16'b0000000000000000;
	sram_mem[114245] = 16'b0000000000000000;
	sram_mem[114246] = 16'b0000000000000000;
	sram_mem[114247] = 16'b0000000000000000;
	sram_mem[114248] = 16'b0000000000000000;
	sram_mem[114249] = 16'b0000000000000000;
	sram_mem[114250] = 16'b0000000000000000;
	sram_mem[114251] = 16'b0000000000000000;
	sram_mem[114252] = 16'b0000000000000000;
	sram_mem[114253] = 16'b0000000000000000;
	sram_mem[114254] = 16'b0000000000000000;
	sram_mem[114255] = 16'b0000000000000000;
	sram_mem[114256] = 16'b0000000000000000;
	sram_mem[114257] = 16'b0000000000000000;
	sram_mem[114258] = 16'b0000000000000000;
	sram_mem[114259] = 16'b0000000000000000;
	sram_mem[114260] = 16'b0000000000000000;
	sram_mem[114261] = 16'b0000000000000000;
	sram_mem[114262] = 16'b0000000000000000;
	sram_mem[114263] = 16'b0000000000000000;
	sram_mem[114264] = 16'b0000000000000000;
	sram_mem[114265] = 16'b0000000000000000;
	sram_mem[114266] = 16'b0000000000000000;
	sram_mem[114267] = 16'b0000000000000000;
	sram_mem[114268] = 16'b0000000000000000;
	sram_mem[114269] = 16'b0000000000000000;
	sram_mem[114270] = 16'b0000000000000000;
	sram_mem[114271] = 16'b0000000000000000;
	sram_mem[114272] = 16'b0000000000000000;
	sram_mem[114273] = 16'b0000000000000000;
	sram_mem[114274] = 16'b0000000000000000;
	sram_mem[114275] = 16'b0000000000000000;
	sram_mem[114276] = 16'b0000000000000000;
	sram_mem[114277] = 16'b0000000000000000;
	sram_mem[114278] = 16'b0000000000000000;
	sram_mem[114279] = 16'b0000000000000000;
	sram_mem[114280] = 16'b0000000000000000;
	sram_mem[114281] = 16'b0000000000000000;
	sram_mem[114282] = 16'b0000000000000000;
	sram_mem[114283] = 16'b0000000000000000;
	sram_mem[114284] = 16'b0000000000000000;
	sram_mem[114285] = 16'b0000000000000000;
	sram_mem[114286] = 16'b0000000000000000;
	sram_mem[114287] = 16'b0000000000000000;
	sram_mem[114288] = 16'b0000000000000000;
	sram_mem[114289] = 16'b0000000000000000;
	sram_mem[114290] = 16'b0000000000000000;
	sram_mem[114291] = 16'b0000000000000000;
	sram_mem[114292] = 16'b0000000000000000;
	sram_mem[114293] = 16'b0000000000000000;
	sram_mem[114294] = 16'b0000000000000000;
	sram_mem[114295] = 16'b0000000000000000;
	sram_mem[114296] = 16'b0000000000000000;
	sram_mem[114297] = 16'b0000000000000000;
	sram_mem[114298] = 16'b0000000000000000;
	sram_mem[114299] = 16'b0000000000000000;
	sram_mem[114300] = 16'b0000000000000000;
	sram_mem[114301] = 16'b0000000000000000;
	sram_mem[114302] = 16'b0000000000000000;
	sram_mem[114303] = 16'b0000000000000000;
	sram_mem[114304] = 16'b0000000000000000;
	sram_mem[114305] = 16'b0000000000000000;
	sram_mem[114306] = 16'b0000000000000000;
	sram_mem[114307] = 16'b0000000000000000;
	sram_mem[114308] = 16'b0000000000000000;
	sram_mem[114309] = 16'b0000000000000000;
	sram_mem[114310] = 16'b0000000000000000;
	sram_mem[114311] = 16'b0000000000000000;
	sram_mem[114312] = 16'b0000000000000000;
	sram_mem[114313] = 16'b0000000000000000;
	sram_mem[114314] = 16'b0000000000000000;
	sram_mem[114315] = 16'b0000000000000000;
	sram_mem[114316] = 16'b0000000000000000;
	sram_mem[114317] = 16'b0000000000000000;
	sram_mem[114318] = 16'b0000000000000000;
	sram_mem[114319] = 16'b0000000000000000;
	sram_mem[114320] = 16'b0000000000000000;
	sram_mem[114321] = 16'b0000000000000000;
	sram_mem[114322] = 16'b0000000000000000;
	sram_mem[114323] = 16'b0000000000000000;
	sram_mem[114324] = 16'b0000000000000000;
	sram_mem[114325] = 16'b0000000000000000;
	sram_mem[114326] = 16'b0000000000000000;
	sram_mem[114327] = 16'b0000000000000000;
	sram_mem[114328] = 16'b0000000000000000;
	sram_mem[114329] = 16'b0000000000000000;
	sram_mem[114330] = 16'b0000000000000000;
	sram_mem[114331] = 16'b0000000000000000;
	sram_mem[114332] = 16'b0000000000000000;
	sram_mem[114333] = 16'b0000000000000000;
	sram_mem[114334] = 16'b0000000000000000;
	sram_mem[114335] = 16'b0000000000000000;
	sram_mem[114336] = 16'b0000000000000000;
	sram_mem[114337] = 16'b0000000000000000;
	sram_mem[114338] = 16'b0000000000000000;
	sram_mem[114339] = 16'b0000000000000000;
	sram_mem[114340] = 16'b0000000000000000;
	sram_mem[114341] = 16'b0000000000000000;
	sram_mem[114342] = 16'b0000000000000000;
	sram_mem[114343] = 16'b0000000000000000;
	sram_mem[114344] = 16'b0000000000000000;
	sram_mem[114345] = 16'b0000000000000000;
	sram_mem[114346] = 16'b0000000000000000;
	sram_mem[114347] = 16'b0000000000000000;
	sram_mem[114348] = 16'b0000000000000000;
	sram_mem[114349] = 16'b0000000000000000;
	sram_mem[114350] = 16'b0000000000000000;
	sram_mem[114351] = 16'b0000000000000000;
	sram_mem[114352] = 16'b0000000000000000;
	sram_mem[114353] = 16'b0000000000000000;
	sram_mem[114354] = 16'b0000000000000000;
	sram_mem[114355] = 16'b0000000000000000;
	sram_mem[114356] = 16'b0000000000000000;
	sram_mem[114357] = 16'b0000000000000000;
	sram_mem[114358] = 16'b0000000000000000;
	sram_mem[114359] = 16'b0000000000000000;
	sram_mem[114360] = 16'b0000000000000000;
	sram_mem[114361] = 16'b0000000000000000;
	sram_mem[114362] = 16'b0000000000000000;
	sram_mem[114363] = 16'b0000000000000000;
	sram_mem[114364] = 16'b0000000000000000;
	sram_mem[114365] = 16'b0000000000000000;
	sram_mem[114366] = 16'b0000000000000000;
	sram_mem[114367] = 16'b0000000000000000;
	sram_mem[114368] = 16'b0000000000000000;
	sram_mem[114369] = 16'b0000000000000000;
	sram_mem[114370] = 16'b0000000000000000;
	sram_mem[114371] = 16'b0000000000000000;
	sram_mem[114372] = 16'b0000000000000000;
	sram_mem[114373] = 16'b0000000000000000;
	sram_mem[114374] = 16'b0000000000000000;
	sram_mem[114375] = 16'b0000000000000000;
	sram_mem[114376] = 16'b0000000000000000;
	sram_mem[114377] = 16'b0000000000000000;
	sram_mem[114378] = 16'b0000000000000000;
	sram_mem[114379] = 16'b0000000000000000;
	sram_mem[114380] = 16'b0000000000000000;
	sram_mem[114381] = 16'b0000000000000000;
	sram_mem[114382] = 16'b0000000000000000;
	sram_mem[114383] = 16'b0000000000000000;
	sram_mem[114384] = 16'b0000000000000000;
	sram_mem[114385] = 16'b0000000000000000;
	sram_mem[114386] = 16'b0000000000000000;
	sram_mem[114387] = 16'b0000000000000000;
	sram_mem[114388] = 16'b0000000000000000;
	sram_mem[114389] = 16'b0000000000000000;
	sram_mem[114390] = 16'b0000000000000000;
	sram_mem[114391] = 16'b0000000000000000;
	sram_mem[114392] = 16'b0000000000000000;
	sram_mem[114393] = 16'b0000000000000000;
	sram_mem[114394] = 16'b0000000000000000;
	sram_mem[114395] = 16'b0000000000000000;
	sram_mem[114396] = 16'b0000000000000000;
	sram_mem[114397] = 16'b0000000000000000;
	sram_mem[114398] = 16'b0000000000000000;
	sram_mem[114399] = 16'b0000000000000000;
	sram_mem[114400] = 16'b0000000000000000;
	sram_mem[114401] = 16'b0000000000000000;
	sram_mem[114402] = 16'b0000000000000000;
	sram_mem[114403] = 16'b0000000000000000;
	sram_mem[114404] = 16'b0000000000000000;
	sram_mem[114405] = 16'b0000000000000000;
	sram_mem[114406] = 16'b0000000000000000;
	sram_mem[114407] = 16'b0000000000000000;
	sram_mem[114408] = 16'b0000000000000000;
	sram_mem[114409] = 16'b0000000000000000;
	sram_mem[114410] = 16'b0000000000000000;
	sram_mem[114411] = 16'b0000000000000000;
	sram_mem[114412] = 16'b0000000000000000;
	sram_mem[114413] = 16'b0000000000000000;
	sram_mem[114414] = 16'b0000000000000000;
	sram_mem[114415] = 16'b0000000000000000;
	sram_mem[114416] = 16'b0000000000000000;
	sram_mem[114417] = 16'b0000000000000000;
	sram_mem[114418] = 16'b0000000000000000;
	sram_mem[114419] = 16'b0000000000000000;
	sram_mem[114420] = 16'b0000000000000000;
	sram_mem[114421] = 16'b0000000000000000;
	sram_mem[114422] = 16'b0000000000000000;
	sram_mem[114423] = 16'b0000000000000000;
	sram_mem[114424] = 16'b0000000000000000;
	sram_mem[114425] = 16'b0000000000000000;
	sram_mem[114426] = 16'b0000000000000000;
	sram_mem[114427] = 16'b0000000000000000;
	sram_mem[114428] = 16'b0000000000000000;
	sram_mem[114429] = 16'b0000000000000000;
	sram_mem[114430] = 16'b0000000000000000;
	sram_mem[114431] = 16'b0000000000000000;
	sram_mem[114432] = 16'b0000000000000000;
	sram_mem[114433] = 16'b0000000000000000;
	sram_mem[114434] = 16'b0000000000000000;
	sram_mem[114435] = 16'b0000000000000000;
	sram_mem[114436] = 16'b0000000000000000;
	sram_mem[114437] = 16'b0000000000000000;
	sram_mem[114438] = 16'b0000000000000000;
	sram_mem[114439] = 16'b0000000000000000;
	sram_mem[114440] = 16'b0000000000000000;
	sram_mem[114441] = 16'b0000000000000000;
	sram_mem[114442] = 16'b0000000000000000;
	sram_mem[114443] = 16'b0000000000000000;
	sram_mem[114444] = 16'b0000000000000000;
	sram_mem[114445] = 16'b0000000000000000;
	sram_mem[114446] = 16'b0000000000000000;
	sram_mem[114447] = 16'b0000000000000000;
	sram_mem[114448] = 16'b0000000000000000;
	sram_mem[114449] = 16'b0000000000000000;
	sram_mem[114450] = 16'b0000000000000000;
	sram_mem[114451] = 16'b0000000000000000;
	sram_mem[114452] = 16'b0000000000000000;
	sram_mem[114453] = 16'b0000000000000000;
	sram_mem[114454] = 16'b0000000000000000;
	sram_mem[114455] = 16'b0000000000000000;
	sram_mem[114456] = 16'b0000000000000000;
	sram_mem[114457] = 16'b0000000000000000;
	sram_mem[114458] = 16'b0000000000000000;
	sram_mem[114459] = 16'b0000000000000000;
	sram_mem[114460] = 16'b0000000000000000;
	sram_mem[114461] = 16'b0000000000000000;
	sram_mem[114462] = 16'b0000000000000000;
	sram_mem[114463] = 16'b0000000000000000;
	sram_mem[114464] = 16'b0000000000000000;
	sram_mem[114465] = 16'b0000000000000000;
	sram_mem[114466] = 16'b0000000000000000;
	sram_mem[114467] = 16'b0000000000000000;
	sram_mem[114468] = 16'b0000000000000000;
	sram_mem[114469] = 16'b0000000000000000;
	sram_mem[114470] = 16'b0000000000000000;
	sram_mem[114471] = 16'b0000000000000000;
	sram_mem[114472] = 16'b0000000000000000;
	sram_mem[114473] = 16'b0000000000000000;
	sram_mem[114474] = 16'b0000000000000000;
	sram_mem[114475] = 16'b0000000000000000;
	sram_mem[114476] = 16'b0000000000000000;
	sram_mem[114477] = 16'b0000000000000000;
	sram_mem[114478] = 16'b0000000000000000;
	sram_mem[114479] = 16'b0000000000000000;
	sram_mem[114480] = 16'b0000000000000000;
	sram_mem[114481] = 16'b0000000000000000;
	sram_mem[114482] = 16'b0000000000000000;
	sram_mem[114483] = 16'b0000000000000000;
	sram_mem[114484] = 16'b0000000000000000;
	sram_mem[114485] = 16'b0000000000000000;
	sram_mem[114486] = 16'b0000000000000000;
	sram_mem[114487] = 16'b0000000000000000;
	sram_mem[114488] = 16'b0000000000000000;
	sram_mem[114489] = 16'b0000000000000000;
	sram_mem[114490] = 16'b0000000000000000;
	sram_mem[114491] = 16'b0000000000000000;
	sram_mem[114492] = 16'b0000000000000000;
	sram_mem[114493] = 16'b0000000000000000;
	sram_mem[114494] = 16'b0000000000000000;
	sram_mem[114495] = 16'b0000000000000000;
	sram_mem[114496] = 16'b0000000000000000;
	sram_mem[114497] = 16'b0000000000000000;
	sram_mem[114498] = 16'b0000000000000000;
	sram_mem[114499] = 16'b0000000000000000;
	sram_mem[114500] = 16'b0000000000000000;
	sram_mem[114501] = 16'b0000000000000000;
	sram_mem[114502] = 16'b0000000000000000;
	sram_mem[114503] = 16'b0000000000000000;
	sram_mem[114504] = 16'b0000000000000000;
	sram_mem[114505] = 16'b0000000000000000;
	sram_mem[114506] = 16'b0000000000000000;
	sram_mem[114507] = 16'b0000000000000000;
	sram_mem[114508] = 16'b0000000000000000;
	sram_mem[114509] = 16'b0000000000000000;
	sram_mem[114510] = 16'b0000000000000000;
	sram_mem[114511] = 16'b0000000000000000;
	sram_mem[114512] = 16'b0000000000000000;
	sram_mem[114513] = 16'b0000000000000000;
	sram_mem[114514] = 16'b0000000000000000;
	sram_mem[114515] = 16'b0000000000000000;
	sram_mem[114516] = 16'b0000000000000000;
	sram_mem[114517] = 16'b0000000000000000;
	sram_mem[114518] = 16'b0000000000000000;
	sram_mem[114519] = 16'b0000000000000000;
	sram_mem[114520] = 16'b0000000000000000;
	sram_mem[114521] = 16'b0000000000000000;
	sram_mem[114522] = 16'b0000000000000000;
	sram_mem[114523] = 16'b0000000000000000;
	sram_mem[114524] = 16'b0000000000000000;
	sram_mem[114525] = 16'b0000000000000000;
	sram_mem[114526] = 16'b0000000000000000;
	sram_mem[114527] = 16'b0000000000000000;
	sram_mem[114528] = 16'b0000000000000000;
	sram_mem[114529] = 16'b0000000000000000;
	sram_mem[114530] = 16'b0000000000000000;
	sram_mem[114531] = 16'b0000000000000000;
	sram_mem[114532] = 16'b0000000000000000;
	sram_mem[114533] = 16'b0000000000000000;
	sram_mem[114534] = 16'b0000000000000000;
	sram_mem[114535] = 16'b0000000000000000;
	sram_mem[114536] = 16'b0000000000000000;
	sram_mem[114537] = 16'b0000000000000000;
	sram_mem[114538] = 16'b0000000000000000;
	sram_mem[114539] = 16'b0000000000000000;
	sram_mem[114540] = 16'b0000000000000000;
	sram_mem[114541] = 16'b0000000000000000;
	sram_mem[114542] = 16'b0000000000000000;
	sram_mem[114543] = 16'b0000000000000000;
	sram_mem[114544] = 16'b0000000000000000;
	sram_mem[114545] = 16'b0000000000000000;
	sram_mem[114546] = 16'b0000000000000000;
	sram_mem[114547] = 16'b0000000000000000;
	sram_mem[114548] = 16'b0000000000000000;
	sram_mem[114549] = 16'b0000000000000000;
	sram_mem[114550] = 16'b0000000000000000;
	sram_mem[114551] = 16'b0000000000000000;
	sram_mem[114552] = 16'b0000000000000000;
	sram_mem[114553] = 16'b0000000000000000;
	sram_mem[114554] = 16'b0000000000000000;
	sram_mem[114555] = 16'b0000000000000000;
	sram_mem[114556] = 16'b0000000000000000;
	sram_mem[114557] = 16'b0000000000000000;
	sram_mem[114558] = 16'b0000000000000000;
	sram_mem[114559] = 16'b0000000000000000;
	sram_mem[114560] = 16'b0000000000000000;
	sram_mem[114561] = 16'b0000000000000000;
	sram_mem[114562] = 16'b0000000000000000;
	sram_mem[114563] = 16'b0000000000000000;
	sram_mem[114564] = 16'b0000000000000000;
	sram_mem[114565] = 16'b0000000000000000;
	sram_mem[114566] = 16'b0000000000000000;
	sram_mem[114567] = 16'b0000000000000000;
	sram_mem[114568] = 16'b0000000000000000;
	sram_mem[114569] = 16'b0000000000000000;
	sram_mem[114570] = 16'b0000000000000000;
	sram_mem[114571] = 16'b0000000000000000;
	sram_mem[114572] = 16'b0000000000000000;
	sram_mem[114573] = 16'b0000000000000000;
	sram_mem[114574] = 16'b0000000000000000;
	sram_mem[114575] = 16'b0000000000000000;
	sram_mem[114576] = 16'b0000000000000000;
	sram_mem[114577] = 16'b0000000000000000;
	sram_mem[114578] = 16'b0000000000000000;
	sram_mem[114579] = 16'b0000000000000000;
	sram_mem[114580] = 16'b0000000000000000;
	sram_mem[114581] = 16'b0000000000000000;
	sram_mem[114582] = 16'b0000000000000000;
	sram_mem[114583] = 16'b0000000000000000;
	sram_mem[114584] = 16'b0000000000000000;
	sram_mem[114585] = 16'b0000000000000000;
	sram_mem[114586] = 16'b0000000000000000;
	sram_mem[114587] = 16'b0000000000000000;
	sram_mem[114588] = 16'b0000000000000000;
	sram_mem[114589] = 16'b0000000000000000;
	sram_mem[114590] = 16'b0000000000000000;
	sram_mem[114591] = 16'b0000000000000000;
	sram_mem[114592] = 16'b0000000000000000;
	sram_mem[114593] = 16'b0000000000000000;
	sram_mem[114594] = 16'b0000000000000000;
	sram_mem[114595] = 16'b0000000000000000;
	sram_mem[114596] = 16'b0000000000000000;
	sram_mem[114597] = 16'b0000000000000000;
	sram_mem[114598] = 16'b0000000000000000;
	sram_mem[114599] = 16'b0000000000000000;
	sram_mem[114600] = 16'b0000000000000000;
	sram_mem[114601] = 16'b0000000000000000;
	sram_mem[114602] = 16'b0000000000000000;
	sram_mem[114603] = 16'b0000000000000000;
	sram_mem[114604] = 16'b0000000000000000;
	sram_mem[114605] = 16'b0000000000000000;
	sram_mem[114606] = 16'b0000000000000000;
	sram_mem[114607] = 16'b0000000000000000;
	sram_mem[114608] = 16'b0000000000000000;
	sram_mem[114609] = 16'b0000000000000000;
	sram_mem[114610] = 16'b0000000000000000;
	sram_mem[114611] = 16'b0000000000000000;
	sram_mem[114612] = 16'b0000000000000000;
	sram_mem[114613] = 16'b0000000000000000;
	sram_mem[114614] = 16'b0000000000000000;
	sram_mem[114615] = 16'b0000000000000000;
	sram_mem[114616] = 16'b0000000000000000;
	sram_mem[114617] = 16'b0000000000000000;
	sram_mem[114618] = 16'b0000000000000000;
	sram_mem[114619] = 16'b0000000000000000;
	sram_mem[114620] = 16'b0000000000000000;
	sram_mem[114621] = 16'b0000000000000000;
	sram_mem[114622] = 16'b0000000000000000;
	sram_mem[114623] = 16'b0000000000000000;
	sram_mem[114624] = 16'b0000000000000000;
	sram_mem[114625] = 16'b0000000000000000;
	sram_mem[114626] = 16'b0000000000000000;
	sram_mem[114627] = 16'b0000000000000000;
	sram_mem[114628] = 16'b0000000000000000;
	sram_mem[114629] = 16'b0000000000000000;
	sram_mem[114630] = 16'b0000000000000000;
	sram_mem[114631] = 16'b0000000000000000;
	sram_mem[114632] = 16'b0000000000000000;
	sram_mem[114633] = 16'b0000000000000000;
	sram_mem[114634] = 16'b0000000000000000;
	sram_mem[114635] = 16'b0000000000000000;
	sram_mem[114636] = 16'b0000000000000000;
	sram_mem[114637] = 16'b0000000000000000;
	sram_mem[114638] = 16'b0000000000000000;
	sram_mem[114639] = 16'b0000000000000000;
	sram_mem[114640] = 16'b0000000000000000;
	sram_mem[114641] = 16'b0000000000000000;
	sram_mem[114642] = 16'b0000000000000000;
	sram_mem[114643] = 16'b0000000000000000;
	sram_mem[114644] = 16'b0000000000000000;
	sram_mem[114645] = 16'b0000000000000000;
	sram_mem[114646] = 16'b0000000000000000;
	sram_mem[114647] = 16'b0000000000000000;
	sram_mem[114648] = 16'b0000000000000000;
	sram_mem[114649] = 16'b0000000000000000;
	sram_mem[114650] = 16'b0000000000000000;
	sram_mem[114651] = 16'b0000000000000000;
	sram_mem[114652] = 16'b0000000000000000;
	sram_mem[114653] = 16'b0000000000000000;
	sram_mem[114654] = 16'b0000000000000000;
	sram_mem[114655] = 16'b0000000000000000;
	sram_mem[114656] = 16'b0000000000000000;
	sram_mem[114657] = 16'b0000000000000000;
	sram_mem[114658] = 16'b0000000000000000;
	sram_mem[114659] = 16'b0000000000000000;
	sram_mem[114660] = 16'b0000000000000000;
	sram_mem[114661] = 16'b0000000000000000;
	sram_mem[114662] = 16'b0000000000000000;
	sram_mem[114663] = 16'b0000000000000000;
	sram_mem[114664] = 16'b0000000000000000;
	sram_mem[114665] = 16'b0000000000000000;
	sram_mem[114666] = 16'b0000000000000000;
	sram_mem[114667] = 16'b0000000000000000;
	sram_mem[114668] = 16'b0000000000000000;
	sram_mem[114669] = 16'b0000000000000000;
	sram_mem[114670] = 16'b0000000000000000;
	sram_mem[114671] = 16'b0000000000000000;
	sram_mem[114672] = 16'b0000000000000000;
	sram_mem[114673] = 16'b0000000000000000;
	sram_mem[114674] = 16'b0000000000000000;
	sram_mem[114675] = 16'b0000000000000000;
	sram_mem[114676] = 16'b0000000000000000;
	sram_mem[114677] = 16'b0000000000000000;
	sram_mem[114678] = 16'b0000000000000000;
	sram_mem[114679] = 16'b0000000000000000;
	sram_mem[114680] = 16'b0000000000000000;
	sram_mem[114681] = 16'b0000000000000000;
	sram_mem[114682] = 16'b0000000000000000;
	sram_mem[114683] = 16'b0000000000000000;
	sram_mem[114684] = 16'b0000000000000000;
	sram_mem[114685] = 16'b0000000000000000;
	sram_mem[114686] = 16'b0000000000000000;
	sram_mem[114687] = 16'b0000000000000000;
	sram_mem[114688] = 16'b0000000000000000;
	sram_mem[114689] = 16'b0000000000000000;
	sram_mem[114690] = 16'b0000000000000000;
	sram_mem[114691] = 16'b0000000000000000;
	sram_mem[114692] = 16'b0000000000000000;
	sram_mem[114693] = 16'b0000000000000000;
	sram_mem[114694] = 16'b0000000000000000;
	sram_mem[114695] = 16'b0000000000000000;
	sram_mem[114696] = 16'b0000000000000000;
	sram_mem[114697] = 16'b0000000000000000;
	sram_mem[114698] = 16'b0000000000000000;
	sram_mem[114699] = 16'b0000000000000000;
	sram_mem[114700] = 16'b0000000000000000;
	sram_mem[114701] = 16'b0000000000000000;
	sram_mem[114702] = 16'b0000000000000000;
	sram_mem[114703] = 16'b0000000000000000;
	sram_mem[114704] = 16'b0000000000000000;
	sram_mem[114705] = 16'b0000000000000000;
	sram_mem[114706] = 16'b0000000000000000;
	sram_mem[114707] = 16'b0000000000000000;
	sram_mem[114708] = 16'b0000000000000000;
	sram_mem[114709] = 16'b0000000000000000;
	sram_mem[114710] = 16'b0000000000000000;
	sram_mem[114711] = 16'b0000000000000000;
	sram_mem[114712] = 16'b0000000000000000;
	sram_mem[114713] = 16'b0000000000000000;
	sram_mem[114714] = 16'b0000000000000000;
	sram_mem[114715] = 16'b0000000000000000;
	sram_mem[114716] = 16'b0000000000000000;
	sram_mem[114717] = 16'b0000000000000000;
	sram_mem[114718] = 16'b0000000000000000;
	sram_mem[114719] = 16'b0000000000000000;
	sram_mem[114720] = 16'b0000000000000000;
	sram_mem[114721] = 16'b0000000000000000;
	sram_mem[114722] = 16'b0000000000000000;
	sram_mem[114723] = 16'b0000000000000000;
	sram_mem[114724] = 16'b0000000000000000;
	sram_mem[114725] = 16'b0000000000000000;
	sram_mem[114726] = 16'b0000000000000000;
	sram_mem[114727] = 16'b0000000000000000;
	sram_mem[114728] = 16'b0000000000000000;
	sram_mem[114729] = 16'b0000000000000000;
	sram_mem[114730] = 16'b0000000000000000;
	sram_mem[114731] = 16'b0000000000000000;
	sram_mem[114732] = 16'b0000000000000000;
	sram_mem[114733] = 16'b0000000000000000;
	sram_mem[114734] = 16'b0000000000000000;
	sram_mem[114735] = 16'b0000000000000000;
	sram_mem[114736] = 16'b0000000000000000;
	sram_mem[114737] = 16'b0000000000000000;
	sram_mem[114738] = 16'b0000000000000000;
	sram_mem[114739] = 16'b0000000000000000;
	sram_mem[114740] = 16'b0000000000000000;
	sram_mem[114741] = 16'b0000000000000000;
	sram_mem[114742] = 16'b0000000000000000;
	sram_mem[114743] = 16'b0000000000000000;
	sram_mem[114744] = 16'b0000000000000000;
	sram_mem[114745] = 16'b0000000000000000;
	sram_mem[114746] = 16'b0000000000000000;
	sram_mem[114747] = 16'b0000000000000000;
	sram_mem[114748] = 16'b0000000000000000;
	sram_mem[114749] = 16'b0000000000000000;
	sram_mem[114750] = 16'b0000000000000000;
	sram_mem[114751] = 16'b0000000000000000;
	sram_mem[114752] = 16'b0000000000000000;
	sram_mem[114753] = 16'b0000000000000000;
	sram_mem[114754] = 16'b0000000000000000;
	sram_mem[114755] = 16'b0000000000000000;
	sram_mem[114756] = 16'b0000000000000000;
	sram_mem[114757] = 16'b0000000000000000;
	sram_mem[114758] = 16'b0000000000000000;
	sram_mem[114759] = 16'b0000000000000000;
	sram_mem[114760] = 16'b0000000000000000;
	sram_mem[114761] = 16'b0000000000000000;
	sram_mem[114762] = 16'b0000000000000000;
	sram_mem[114763] = 16'b0000000000000000;
	sram_mem[114764] = 16'b0000000000000000;
	sram_mem[114765] = 16'b0000000000000000;
	sram_mem[114766] = 16'b0000000000000000;
	sram_mem[114767] = 16'b0000000000000000;
	sram_mem[114768] = 16'b0000000000000000;
	sram_mem[114769] = 16'b0000000000000000;
	sram_mem[114770] = 16'b0000000000000000;
	sram_mem[114771] = 16'b0000000000000000;
	sram_mem[114772] = 16'b0000000000000000;
	sram_mem[114773] = 16'b0000000000000000;
	sram_mem[114774] = 16'b0000000000000000;
	sram_mem[114775] = 16'b0000000000000000;
	sram_mem[114776] = 16'b0000000000000000;
	sram_mem[114777] = 16'b0000000000000000;
	sram_mem[114778] = 16'b0000000000000000;
	sram_mem[114779] = 16'b0000000000000000;
	sram_mem[114780] = 16'b0000000000000000;
	sram_mem[114781] = 16'b0000000000000000;
	sram_mem[114782] = 16'b0000000000000000;
	sram_mem[114783] = 16'b0000000000000000;
	sram_mem[114784] = 16'b0000000000000000;
	sram_mem[114785] = 16'b0000000000000000;
	sram_mem[114786] = 16'b0000000000000000;
	sram_mem[114787] = 16'b0000000000000000;
	sram_mem[114788] = 16'b0000000000000000;
	sram_mem[114789] = 16'b0000000000000000;
	sram_mem[114790] = 16'b0000000000000000;
	sram_mem[114791] = 16'b0000000000000000;
	sram_mem[114792] = 16'b0000000000000000;
	sram_mem[114793] = 16'b0000000000000000;
	sram_mem[114794] = 16'b0000000000000000;
	sram_mem[114795] = 16'b0000000000000000;
	sram_mem[114796] = 16'b0000000000000000;
	sram_mem[114797] = 16'b0000000000000000;
	sram_mem[114798] = 16'b0000000000000000;
	sram_mem[114799] = 16'b0000000000000000;
	sram_mem[114800] = 16'b0000000000000000;
	sram_mem[114801] = 16'b0000000000000000;
	sram_mem[114802] = 16'b0000000000000000;
	sram_mem[114803] = 16'b0000000000000000;
	sram_mem[114804] = 16'b0000000000000000;
	sram_mem[114805] = 16'b0000000000000000;
	sram_mem[114806] = 16'b0000000000000000;
	sram_mem[114807] = 16'b0000000000000000;
	sram_mem[114808] = 16'b0000000000000000;
	sram_mem[114809] = 16'b0000000000000000;
	sram_mem[114810] = 16'b0000000000000000;
	sram_mem[114811] = 16'b0000000000000000;
	sram_mem[114812] = 16'b0000000000000000;
	sram_mem[114813] = 16'b0000000000000000;
	sram_mem[114814] = 16'b0000000000000000;
	sram_mem[114815] = 16'b0000000000000000;
	sram_mem[114816] = 16'b0000000000000000;
	sram_mem[114817] = 16'b0000000000000000;
	sram_mem[114818] = 16'b0000000000000000;
	sram_mem[114819] = 16'b0000000000000000;
	sram_mem[114820] = 16'b0000000000000000;
	sram_mem[114821] = 16'b0000000000000000;
	sram_mem[114822] = 16'b0000000000000000;
	sram_mem[114823] = 16'b0000000000000000;
	sram_mem[114824] = 16'b0000000000000000;
	sram_mem[114825] = 16'b0000000000000000;
	sram_mem[114826] = 16'b0000000000000000;
	sram_mem[114827] = 16'b0000000000000000;
	sram_mem[114828] = 16'b0000000000000000;
	sram_mem[114829] = 16'b0000000000000000;
	sram_mem[114830] = 16'b0000000000000000;
	sram_mem[114831] = 16'b0000000000000000;
	sram_mem[114832] = 16'b0000000000000000;
	sram_mem[114833] = 16'b0000000000000000;
	sram_mem[114834] = 16'b0000000000000000;
	sram_mem[114835] = 16'b0000000000000000;
	sram_mem[114836] = 16'b0000000000000000;
	sram_mem[114837] = 16'b0000000000000000;
	sram_mem[114838] = 16'b0000000000000000;
	sram_mem[114839] = 16'b0000000000000000;
	sram_mem[114840] = 16'b0000000000000000;
	sram_mem[114841] = 16'b0000000000000000;
	sram_mem[114842] = 16'b0000000000000000;
	sram_mem[114843] = 16'b0000000000000000;
	sram_mem[114844] = 16'b0000000000000000;
	sram_mem[114845] = 16'b0000000000000000;
	sram_mem[114846] = 16'b0000000000000000;
	sram_mem[114847] = 16'b0000000000000000;
	sram_mem[114848] = 16'b0000000000000000;
	sram_mem[114849] = 16'b0000000000000000;
	sram_mem[114850] = 16'b0000000000000000;
	sram_mem[114851] = 16'b0000000000000000;
	sram_mem[114852] = 16'b0000000000000000;
	sram_mem[114853] = 16'b0000000000000000;
	sram_mem[114854] = 16'b0000000000000000;
	sram_mem[114855] = 16'b0000000000000000;
	sram_mem[114856] = 16'b0000000000000000;
	sram_mem[114857] = 16'b0000000000000000;
	sram_mem[114858] = 16'b0000000000000000;
	sram_mem[114859] = 16'b0000000000000000;
	sram_mem[114860] = 16'b0000000000000000;
	sram_mem[114861] = 16'b0000000000000000;
	sram_mem[114862] = 16'b0000000000000000;
	sram_mem[114863] = 16'b0000000000000000;
	sram_mem[114864] = 16'b0000000000000000;
	sram_mem[114865] = 16'b0000000000000000;
	sram_mem[114866] = 16'b0000000000000000;
	sram_mem[114867] = 16'b0000000000000000;
	sram_mem[114868] = 16'b0000000000000000;
	sram_mem[114869] = 16'b0000000000000000;
	sram_mem[114870] = 16'b0000000000000000;
	sram_mem[114871] = 16'b0000000000000000;
	sram_mem[114872] = 16'b0000000000000000;
	sram_mem[114873] = 16'b0000000000000000;
	sram_mem[114874] = 16'b0000000000000000;
	sram_mem[114875] = 16'b0000000000000000;
	sram_mem[114876] = 16'b0000000000000000;
	sram_mem[114877] = 16'b0000000000000000;
	sram_mem[114878] = 16'b0000000000000000;
	sram_mem[114879] = 16'b0000000000000000;
	sram_mem[114880] = 16'b0000000000000000;
	sram_mem[114881] = 16'b0000000000000000;
	sram_mem[114882] = 16'b0000000000000000;
	sram_mem[114883] = 16'b0000000000000000;
	sram_mem[114884] = 16'b0000000000000000;
	sram_mem[114885] = 16'b0000000000000000;
	sram_mem[114886] = 16'b0000000000000000;
	sram_mem[114887] = 16'b0000000000000000;
	sram_mem[114888] = 16'b0000000000000000;
	sram_mem[114889] = 16'b0000000000000000;
	sram_mem[114890] = 16'b0000000000000000;
	sram_mem[114891] = 16'b0000000000000000;
	sram_mem[114892] = 16'b0000000000000000;
	sram_mem[114893] = 16'b0000000000000000;
	sram_mem[114894] = 16'b0000000000000000;
	sram_mem[114895] = 16'b0000000000000000;
	sram_mem[114896] = 16'b0000000000000000;
	sram_mem[114897] = 16'b0000000000000000;
	sram_mem[114898] = 16'b0000000000000000;
	sram_mem[114899] = 16'b0000000000000000;
	sram_mem[114900] = 16'b0000000000000000;
	sram_mem[114901] = 16'b0000000000000000;
	sram_mem[114902] = 16'b0000000000000000;
	sram_mem[114903] = 16'b0000000000000000;
	sram_mem[114904] = 16'b0000000000000000;
	sram_mem[114905] = 16'b0000000000000000;
	sram_mem[114906] = 16'b0000000000000000;
	sram_mem[114907] = 16'b0000000000000000;
	sram_mem[114908] = 16'b0000000000000000;
	sram_mem[114909] = 16'b0000000000000000;
	sram_mem[114910] = 16'b0000000000000000;
	sram_mem[114911] = 16'b0000000000000000;
	sram_mem[114912] = 16'b0000000000000000;
	sram_mem[114913] = 16'b0000000000000000;
	sram_mem[114914] = 16'b0000000000000000;
	sram_mem[114915] = 16'b0000000000000000;
	sram_mem[114916] = 16'b0000000000000000;
	sram_mem[114917] = 16'b0000000000000000;
	sram_mem[114918] = 16'b0000000000000000;
	sram_mem[114919] = 16'b0000000000000000;
	sram_mem[114920] = 16'b0000000000000000;
	sram_mem[114921] = 16'b0000000000000000;
	sram_mem[114922] = 16'b0000000000000000;
	sram_mem[114923] = 16'b0000000000000000;
	sram_mem[114924] = 16'b0000000000000000;
	sram_mem[114925] = 16'b0000000000000000;
	sram_mem[114926] = 16'b0000000000000000;
	sram_mem[114927] = 16'b0000000000000000;
	sram_mem[114928] = 16'b0000000000000000;
	sram_mem[114929] = 16'b0000000000000000;
	sram_mem[114930] = 16'b0000000000000000;
	sram_mem[114931] = 16'b0000000000000000;
	sram_mem[114932] = 16'b0000000000000000;
	sram_mem[114933] = 16'b0000000000000000;
	sram_mem[114934] = 16'b0000000000000000;
	sram_mem[114935] = 16'b0000000000000000;
	sram_mem[114936] = 16'b0000000000000000;
	sram_mem[114937] = 16'b0000000000000000;
	sram_mem[114938] = 16'b0000000000000000;
	sram_mem[114939] = 16'b0000000000000000;
	sram_mem[114940] = 16'b0000000000000000;
	sram_mem[114941] = 16'b0000000000000000;
	sram_mem[114942] = 16'b0000000000000000;
	sram_mem[114943] = 16'b0000000000000000;
	sram_mem[114944] = 16'b0000000000000000;
	sram_mem[114945] = 16'b0000000000000000;
	sram_mem[114946] = 16'b0000000000000000;
	sram_mem[114947] = 16'b0000000000000000;
	sram_mem[114948] = 16'b0000000000000000;
	sram_mem[114949] = 16'b0000000000000000;
	sram_mem[114950] = 16'b0000000000000000;
	sram_mem[114951] = 16'b0000000000000000;
	sram_mem[114952] = 16'b0000000000000000;
	sram_mem[114953] = 16'b0000000000000000;
	sram_mem[114954] = 16'b0000000000000000;
	sram_mem[114955] = 16'b0000000000000000;
	sram_mem[114956] = 16'b0000000000000000;
	sram_mem[114957] = 16'b0000000000000000;
	sram_mem[114958] = 16'b0000000000000000;
	sram_mem[114959] = 16'b0000000000000000;
	sram_mem[114960] = 16'b0000000000000000;
	sram_mem[114961] = 16'b0000000000000000;
	sram_mem[114962] = 16'b0000000000000000;
	sram_mem[114963] = 16'b0000000000000000;
	sram_mem[114964] = 16'b0000000000000000;
	sram_mem[114965] = 16'b0000000000000000;
	sram_mem[114966] = 16'b0000000000000000;
	sram_mem[114967] = 16'b0000000000000000;
	sram_mem[114968] = 16'b0000000000000000;
	sram_mem[114969] = 16'b0000000000000000;
	sram_mem[114970] = 16'b0000000000000000;
	sram_mem[114971] = 16'b0000000000000000;
	sram_mem[114972] = 16'b0000000000000000;
	sram_mem[114973] = 16'b0000000000000000;
	sram_mem[114974] = 16'b0000000000000000;
	sram_mem[114975] = 16'b0000000000000000;
	sram_mem[114976] = 16'b0000000000000000;
	sram_mem[114977] = 16'b0000000000000000;
	sram_mem[114978] = 16'b0000000000000000;
	sram_mem[114979] = 16'b0000000000000000;
	sram_mem[114980] = 16'b0000000000000000;
	sram_mem[114981] = 16'b0000000000000000;
	sram_mem[114982] = 16'b0000000000000000;
	sram_mem[114983] = 16'b0000000000000000;
	sram_mem[114984] = 16'b0000000000000000;
	sram_mem[114985] = 16'b0000000000000000;
	sram_mem[114986] = 16'b0000000000000000;
	sram_mem[114987] = 16'b0000000000000000;
	sram_mem[114988] = 16'b0000000000000000;
	sram_mem[114989] = 16'b0000000000000000;
	sram_mem[114990] = 16'b0000000000000000;
	sram_mem[114991] = 16'b0000000000000000;
	sram_mem[114992] = 16'b0000000000000000;
	sram_mem[114993] = 16'b0000000000000000;
	sram_mem[114994] = 16'b0000000000000000;
	sram_mem[114995] = 16'b0000000000000000;
	sram_mem[114996] = 16'b0000000000000000;
	sram_mem[114997] = 16'b0000000000000000;
	sram_mem[114998] = 16'b0000000000000000;
	sram_mem[114999] = 16'b0000000000000000;
	sram_mem[115000] = 16'b0000000000000000;
	sram_mem[115001] = 16'b0000000000000000;
	sram_mem[115002] = 16'b0000000000000000;
	sram_mem[115003] = 16'b0000000000000000;
	sram_mem[115004] = 16'b0000000000000000;
	sram_mem[115005] = 16'b0000000000000000;
	sram_mem[115006] = 16'b0000000000000000;
	sram_mem[115007] = 16'b0000000000000000;
	sram_mem[115008] = 16'b0000000000000000;
	sram_mem[115009] = 16'b0000000000000000;
	sram_mem[115010] = 16'b0000000000000000;
	sram_mem[115011] = 16'b0000000000000000;
	sram_mem[115012] = 16'b0000000000000000;
	sram_mem[115013] = 16'b0000000000000000;
	sram_mem[115014] = 16'b0000000000000000;
	sram_mem[115015] = 16'b0000000000000000;
	sram_mem[115016] = 16'b0000000000000000;
	sram_mem[115017] = 16'b0000000000000000;
	sram_mem[115018] = 16'b0000000000000000;
	sram_mem[115019] = 16'b0000000000000000;
	sram_mem[115020] = 16'b0000000000000000;
	sram_mem[115021] = 16'b0000000000000000;
	sram_mem[115022] = 16'b0000000000000000;
	sram_mem[115023] = 16'b0000000000000000;
	sram_mem[115024] = 16'b0000000000000000;
	sram_mem[115025] = 16'b0000000000000000;
	sram_mem[115026] = 16'b0000000000000000;
	sram_mem[115027] = 16'b0000000000000000;
	sram_mem[115028] = 16'b0000000000000000;
	sram_mem[115029] = 16'b0000000000000000;
	sram_mem[115030] = 16'b0000000000000000;
	sram_mem[115031] = 16'b0000000000000000;
	sram_mem[115032] = 16'b0000000000000000;
	sram_mem[115033] = 16'b0000000000000000;
	sram_mem[115034] = 16'b0000000000000000;
	sram_mem[115035] = 16'b0000000000000000;
	sram_mem[115036] = 16'b0000000000000000;
	sram_mem[115037] = 16'b0000000000000000;
	sram_mem[115038] = 16'b0000000000000000;
	sram_mem[115039] = 16'b0000000000000000;
	sram_mem[115040] = 16'b0000000000000000;
	sram_mem[115041] = 16'b0000000000000000;
	sram_mem[115042] = 16'b0000000000000000;
	sram_mem[115043] = 16'b0000000000000000;
	sram_mem[115044] = 16'b0000000000000000;
	sram_mem[115045] = 16'b0000000000000000;
	sram_mem[115046] = 16'b0000000000000000;
	sram_mem[115047] = 16'b0000000000000000;
	sram_mem[115048] = 16'b0000000000000000;
	sram_mem[115049] = 16'b0000000000000000;
	sram_mem[115050] = 16'b0000000000000000;
	sram_mem[115051] = 16'b0000000000000000;
	sram_mem[115052] = 16'b0000000000000000;
	sram_mem[115053] = 16'b0000000000000000;
	sram_mem[115054] = 16'b0000000000000000;
	sram_mem[115055] = 16'b0000000000000000;
	sram_mem[115056] = 16'b0000000000000000;
	sram_mem[115057] = 16'b0000000000000000;
	sram_mem[115058] = 16'b0000000000000000;
	sram_mem[115059] = 16'b0000000000000000;
	sram_mem[115060] = 16'b0000000000000000;
	sram_mem[115061] = 16'b0000000000000000;
	sram_mem[115062] = 16'b0000000000000000;
	sram_mem[115063] = 16'b0000000000000000;
	sram_mem[115064] = 16'b0000000000000000;
	sram_mem[115065] = 16'b0000000000000000;
	sram_mem[115066] = 16'b0000000000000000;
	sram_mem[115067] = 16'b0000000000000000;
	sram_mem[115068] = 16'b0000000000000000;
	sram_mem[115069] = 16'b0000000000000000;
	sram_mem[115070] = 16'b0000000000000000;
	sram_mem[115071] = 16'b0000000000000000;
	sram_mem[115072] = 16'b0000000000000000;
	sram_mem[115073] = 16'b0000000000000000;
	sram_mem[115074] = 16'b0000000000000000;
	sram_mem[115075] = 16'b0000000000000000;
	sram_mem[115076] = 16'b0000000000000000;
	sram_mem[115077] = 16'b0000000000000000;
	sram_mem[115078] = 16'b0000000000000000;
	sram_mem[115079] = 16'b0000000000000000;
	sram_mem[115080] = 16'b0000000000000000;
	sram_mem[115081] = 16'b0000000000000000;
	sram_mem[115082] = 16'b0000000000000000;
	sram_mem[115083] = 16'b0000000000000000;
	sram_mem[115084] = 16'b0000000000000000;
	sram_mem[115085] = 16'b0000000000000000;
	sram_mem[115086] = 16'b0000000000000000;
	sram_mem[115087] = 16'b0000000000000000;
	sram_mem[115088] = 16'b0000000000000000;
	sram_mem[115089] = 16'b0000000000000000;
	sram_mem[115090] = 16'b0000000000000000;
	sram_mem[115091] = 16'b0000000000000000;
	sram_mem[115092] = 16'b0000000000000000;
	sram_mem[115093] = 16'b0000000000000000;
	sram_mem[115094] = 16'b0000000000000000;
	sram_mem[115095] = 16'b0000000000000000;
	sram_mem[115096] = 16'b0000000000000000;
	sram_mem[115097] = 16'b0000000000000000;
	sram_mem[115098] = 16'b0000000000000000;
	sram_mem[115099] = 16'b0000000000000000;
	sram_mem[115100] = 16'b0000000000000000;
	sram_mem[115101] = 16'b0000000000000000;
	sram_mem[115102] = 16'b0000000000000000;
	sram_mem[115103] = 16'b0000000000000000;
	sram_mem[115104] = 16'b0000000000000000;
	sram_mem[115105] = 16'b0000000000000000;
	sram_mem[115106] = 16'b0000000000000000;
	sram_mem[115107] = 16'b0000000000000000;
	sram_mem[115108] = 16'b0000000000000000;
	sram_mem[115109] = 16'b0000000000000000;
	sram_mem[115110] = 16'b0000000000000000;
	sram_mem[115111] = 16'b0000000000000000;
	sram_mem[115112] = 16'b0000000000000000;
	sram_mem[115113] = 16'b0000000000000000;
	sram_mem[115114] = 16'b0000000000000000;
	sram_mem[115115] = 16'b0000000000000000;
	sram_mem[115116] = 16'b0000000000000000;
	sram_mem[115117] = 16'b0000000000000000;
	sram_mem[115118] = 16'b0000000000000000;
	sram_mem[115119] = 16'b0000000000000000;
	sram_mem[115120] = 16'b0000000000000000;
	sram_mem[115121] = 16'b0000000000000000;
	sram_mem[115122] = 16'b0000000000000000;
	sram_mem[115123] = 16'b0000000000000000;
	sram_mem[115124] = 16'b0000000000000000;
	sram_mem[115125] = 16'b0000000000000000;
	sram_mem[115126] = 16'b0000000000000000;
	sram_mem[115127] = 16'b0000000000000000;
	sram_mem[115128] = 16'b0000000000000000;
	sram_mem[115129] = 16'b0000000000000000;
	sram_mem[115130] = 16'b0000000000000000;
	sram_mem[115131] = 16'b0000000000000000;
	sram_mem[115132] = 16'b0000000000000000;
	sram_mem[115133] = 16'b0000000000000000;
	sram_mem[115134] = 16'b0000000000000000;
	sram_mem[115135] = 16'b0000000000000000;
	sram_mem[115136] = 16'b0000000000000000;
	sram_mem[115137] = 16'b0000000000000000;
	sram_mem[115138] = 16'b0000000000000000;
	sram_mem[115139] = 16'b0000000000000000;
	sram_mem[115140] = 16'b0000000000000000;
	sram_mem[115141] = 16'b0000000000000000;
	sram_mem[115142] = 16'b0000000000000000;
	sram_mem[115143] = 16'b0000000000000000;
	sram_mem[115144] = 16'b0000000000000000;
	sram_mem[115145] = 16'b0000000000000000;
	sram_mem[115146] = 16'b0000000000000000;
	sram_mem[115147] = 16'b0000000000000000;
	sram_mem[115148] = 16'b0000000000000000;
	sram_mem[115149] = 16'b0000000000000000;
	sram_mem[115150] = 16'b0000000000000000;
	sram_mem[115151] = 16'b0000000000000000;
	sram_mem[115152] = 16'b0000000000000000;
	sram_mem[115153] = 16'b0000000000000000;
	sram_mem[115154] = 16'b0000000000000000;
	sram_mem[115155] = 16'b0000000000000000;
	sram_mem[115156] = 16'b0000000000000000;
	sram_mem[115157] = 16'b0000000000000000;
	sram_mem[115158] = 16'b0000000000000000;
	sram_mem[115159] = 16'b0000000000000000;
	sram_mem[115160] = 16'b0000000000000000;
	sram_mem[115161] = 16'b0000000000000000;
	sram_mem[115162] = 16'b0000000000000000;
	sram_mem[115163] = 16'b0000000000000000;
	sram_mem[115164] = 16'b0000000000000000;
	sram_mem[115165] = 16'b0000000000000000;
	sram_mem[115166] = 16'b0000000000000000;
	sram_mem[115167] = 16'b0000000000000000;
	sram_mem[115168] = 16'b0000000000000000;
	sram_mem[115169] = 16'b0000000000000000;
	sram_mem[115170] = 16'b0000000000000000;
	sram_mem[115171] = 16'b0000000000000000;
	sram_mem[115172] = 16'b0000000000000000;
	sram_mem[115173] = 16'b0000000000000000;
	sram_mem[115174] = 16'b0000000000000000;
	sram_mem[115175] = 16'b0000000000000000;
	sram_mem[115176] = 16'b0000000000000000;
	sram_mem[115177] = 16'b0000000000000000;
	sram_mem[115178] = 16'b0000000000000000;
	sram_mem[115179] = 16'b0000000000000000;
	sram_mem[115180] = 16'b0000000000000000;
	sram_mem[115181] = 16'b0000000000000000;
	sram_mem[115182] = 16'b0000000000000000;
	sram_mem[115183] = 16'b0000000000000000;
	sram_mem[115184] = 16'b0000000000000000;
	sram_mem[115185] = 16'b0000000000000000;
	sram_mem[115186] = 16'b0000000000000000;
	sram_mem[115187] = 16'b0000000000000000;
	sram_mem[115188] = 16'b0000000000000000;
	sram_mem[115189] = 16'b0000000000000000;
	sram_mem[115190] = 16'b0000000000000000;
	sram_mem[115191] = 16'b0000000000000000;
	sram_mem[115192] = 16'b0000000000000000;
	sram_mem[115193] = 16'b0000000000000000;
	sram_mem[115194] = 16'b0000000000000000;
	sram_mem[115195] = 16'b0000000000000000;
	sram_mem[115196] = 16'b0000000000000000;
	sram_mem[115197] = 16'b0000000000000000;
	sram_mem[115198] = 16'b0000000000000000;
	sram_mem[115199] = 16'b0000000000000000;
	sram_mem[115200] = 16'b0000000000000000;
	sram_mem[115201] = 16'b0000000000000000;
	sram_mem[115202] = 16'b0000000000000000;
	sram_mem[115203] = 16'b0000000000000000;
	sram_mem[115204] = 16'b0000000000000000;
	sram_mem[115205] = 16'b0000000000000000;
	sram_mem[115206] = 16'b0000000000000000;
	sram_mem[115207] = 16'b0000000000000000;
	sram_mem[115208] = 16'b0000000000000000;
	sram_mem[115209] = 16'b0000000000000000;
	sram_mem[115210] = 16'b0000000000000000;
	sram_mem[115211] = 16'b0000000000000000;
	sram_mem[115212] = 16'b0000000000000000;
	sram_mem[115213] = 16'b0000000000000000;
	sram_mem[115214] = 16'b0000000000000000;
	sram_mem[115215] = 16'b0000000000000000;
	sram_mem[115216] = 16'b0000000000000000;
	sram_mem[115217] = 16'b0000000000000000;
	sram_mem[115218] = 16'b0000000000000000;
	sram_mem[115219] = 16'b0000000000000000;
	sram_mem[115220] = 16'b0000000000000000;
	sram_mem[115221] = 16'b0000000000000000;
	sram_mem[115222] = 16'b0000000000000000;
	sram_mem[115223] = 16'b0000000000000000;
	sram_mem[115224] = 16'b0000000000000000;
	sram_mem[115225] = 16'b0000000000000000;
	sram_mem[115226] = 16'b0000000000000000;
	sram_mem[115227] = 16'b0000000000000000;
	sram_mem[115228] = 16'b0000000000000000;
	sram_mem[115229] = 16'b0000000000000000;
	sram_mem[115230] = 16'b0000000000000000;
	sram_mem[115231] = 16'b0000000000000000;
	sram_mem[115232] = 16'b0000000000000000;
	sram_mem[115233] = 16'b0000000000000000;
	sram_mem[115234] = 16'b0000000000000000;
	sram_mem[115235] = 16'b0000000000000000;
	sram_mem[115236] = 16'b0000000000000000;
	sram_mem[115237] = 16'b0000000000000000;
	sram_mem[115238] = 16'b0000000000000000;
	sram_mem[115239] = 16'b0000000000000000;
	sram_mem[115240] = 16'b0000000000000000;
	sram_mem[115241] = 16'b0000000000000000;
	sram_mem[115242] = 16'b0000000000000000;
	sram_mem[115243] = 16'b0000000000000000;
	sram_mem[115244] = 16'b0000000000000000;
	sram_mem[115245] = 16'b0000000000000000;
	sram_mem[115246] = 16'b0000000000000000;
	sram_mem[115247] = 16'b0000000000000000;
	sram_mem[115248] = 16'b0000000000000000;
	sram_mem[115249] = 16'b0000000000000000;
	sram_mem[115250] = 16'b0000000000000000;
	sram_mem[115251] = 16'b0000000000000000;
	sram_mem[115252] = 16'b0000000000000000;
	sram_mem[115253] = 16'b0000000000000000;
	sram_mem[115254] = 16'b0000000000000000;
	sram_mem[115255] = 16'b0000000000000000;
	sram_mem[115256] = 16'b0000000000000000;
	sram_mem[115257] = 16'b0000000000000000;
	sram_mem[115258] = 16'b0000000000000000;
	sram_mem[115259] = 16'b0000000000000000;
	sram_mem[115260] = 16'b0000000000000000;
	sram_mem[115261] = 16'b0000000000000000;
	sram_mem[115262] = 16'b0000000000000000;
	sram_mem[115263] = 16'b0000000000000000;
	sram_mem[115264] = 16'b0000000000000000;
	sram_mem[115265] = 16'b0000000000000000;
	sram_mem[115266] = 16'b0000000000000000;
	sram_mem[115267] = 16'b0000000000000000;
	sram_mem[115268] = 16'b0000000000000000;
	sram_mem[115269] = 16'b0000000000000000;
	sram_mem[115270] = 16'b0000000000000000;
	sram_mem[115271] = 16'b0000000000000000;
	sram_mem[115272] = 16'b0000000000000000;
	sram_mem[115273] = 16'b0000000000000000;
	sram_mem[115274] = 16'b0000000000000000;
	sram_mem[115275] = 16'b0000000000000000;
	sram_mem[115276] = 16'b0000000000000000;
	sram_mem[115277] = 16'b0000000000000000;
	sram_mem[115278] = 16'b0000000000000000;
	sram_mem[115279] = 16'b0000000000000000;
	sram_mem[115280] = 16'b0000000000000000;
	sram_mem[115281] = 16'b0000000000000000;
	sram_mem[115282] = 16'b0000000000000000;
	sram_mem[115283] = 16'b0000000000000000;
	sram_mem[115284] = 16'b0000000000000000;
	sram_mem[115285] = 16'b0000000000000000;
	sram_mem[115286] = 16'b0000000000000000;
	sram_mem[115287] = 16'b0000000000000000;
	sram_mem[115288] = 16'b0000000000000000;
	sram_mem[115289] = 16'b0000000000000000;
	sram_mem[115290] = 16'b0000000000000000;
	sram_mem[115291] = 16'b0000000000000000;
	sram_mem[115292] = 16'b0000000000000000;
	sram_mem[115293] = 16'b0000000000000000;
	sram_mem[115294] = 16'b0000000000000000;
	sram_mem[115295] = 16'b0000000000000000;
	sram_mem[115296] = 16'b0000000000000000;
	sram_mem[115297] = 16'b0000000000000000;
	sram_mem[115298] = 16'b0000000000000000;
	sram_mem[115299] = 16'b0000000000000000;
	sram_mem[115300] = 16'b0000000000000000;
	sram_mem[115301] = 16'b0000000000000000;
	sram_mem[115302] = 16'b0000000000000000;
	sram_mem[115303] = 16'b0000000000000000;
	sram_mem[115304] = 16'b0000000000000000;
	sram_mem[115305] = 16'b0000000000000000;
	sram_mem[115306] = 16'b0000000000000000;
	sram_mem[115307] = 16'b0000000000000000;
	sram_mem[115308] = 16'b0000000000000000;
	sram_mem[115309] = 16'b0000000000000000;
	sram_mem[115310] = 16'b0000000000000000;
	sram_mem[115311] = 16'b0000000000000000;
	sram_mem[115312] = 16'b0000000000000000;
	sram_mem[115313] = 16'b0000000000000000;
	sram_mem[115314] = 16'b0000000000000000;
	sram_mem[115315] = 16'b0000000000000000;
	sram_mem[115316] = 16'b0000000000000000;
	sram_mem[115317] = 16'b0000000000000000;
	sram_mem[115318] = 16'b0000000000000000;
	sram_mem[115319] = 16'b0000000000000000;
	sram_mem[115320] = 16'b0000000000000000;
	sram_mem[115321] = 16'b0000000000000000;
	sram_mem[115322] = 16'b0000000000000000;
	sram_mem[115323] = 16'b0000000000000000;
	sram_mem[115324] = 16'b0000000000000000;
	sram_mem[115325] = 16'b0000000000000000;
	sram_mem[115326] = 16'b0000000000000000;
	sram_mem[115327] = 16'b0000000000000000;
	sram_mem[115328] = 16'b0000000000000000;
	sram_mem[115329] = 16'b0000000000000000;
	sram_mem[115330] = 16'b0000000000000000;
	sram_mem[115331] = 16'b0000000000000000;
	sram_mem[115332] = 16'b0000000000000000;
	sram_mem[115333] = 16'b0000000000000000;
	sram_mem[115334] = 16'b0000000000000000;
	sram_mem[115335] = 16'b0000000000000000;
	sram_mem[115336] = 16'b0000000000000000;
	sram_mem[115337] = 16'b0000000000000000;
	sram_mem[115338] = 16'b0000000000000000;
	sram_mem[115339] = 16'b0000000000000000;
	sram_mem[115340] = 16'b0000000000000000;
	sram_mem[115341] = 16'b0000000000000000;
	sram_mem[115342] = 16'b0000000000000000;
	sram_mem[115343] = 16'b0000000000000000;
	sram_mem[115344] = 16'b0000000000000000;
	sram_mem[115345] = 16'b0000000000000000;
	sram_mem[115346] = 16'b0000000000000000;
	sram_mem[115347] = 16'b0000000000000000;
	sram_mem[115348] = 16'b0000000000000000;
	sram_mem[115349] = 16'b0000000000000000;
	sram_mem[115350] = 16'b0000000000000000;
	sram_mem[115351] = 16'b0000000000000000;
	sram_mem[115352] = 16'b0000000000000000;
	sram_mem[115353] = 16'b0000000000000000;
	sram_mem[115354] = 16'b0000000000000000;
	sram_mem[115355] = 16'b0000000000000000;
	sram_mem[115356] = 16'b0000000000000000;
	sram_mem[115357] = 16'b0000000000000000;
	sram_mem[115358] = 16'b0000000000000000;
	sram_mem[115359] = 16'b0000000000000000;
	sram_mem[115360] = 16'b0000000000000000;
	sram_mem[115361] = 16'b0000000000000000;
	sram_mem[115362] = 16'b0000000000000000;
	sram_mem[115363] = 16'b0000000000000000;
	sram_mem[115364] = 16'b0000000000000000;
	sram_mem[115365] = 16'b0000000000000000;
	sram_mem[115366] = 16'b0000000000000000;
	sram_mem[115367] = 16'b0000000000000000;
	sram_mem[115368] = 16'b0000000000000000;
	sram_mem[115369] = 16'b0000000000000000;
	sram_mem[115370] = 16'b0000000000000000;
	sram_mem[115371] = 16'b0000000000000000;
	sram_mem[115372] = 16'b0000000000000000;
	sram_mem[115373] = 16'b0000000000000000;
	sram_mem[115374] = 16'b0000000000000000;
	sram_mem[115375] = 16'b0000000000000000;
	sram_mem[115376] = 16'b0000000000000000;
	sram_mem[115377] = 16'b0000000000000000;
	sram_mem[115378] = 16'b0000000000000000;
	sram_mem[115379] = 16'b0000000000000000;
	sram_mem[115380] = 16'b0000000000000000;
	sram_mem[115381] = 16'b0000000000000000;
	sram_mem[115382] = 16'b0000000000000000;
	sram_mem[115383] = 16'b0000000000000000;
	sram_mem[115384] = 16'b0000000000000000;
	sram_mem[115385] = 16'b0000000000000000;
	sram_mem[115386] = 16'b0000000000000000;
	sram_mem[115387] = 16'b0000000000000000;
	sram_mem[115388] = 16'b0000000000000000;
	sram_mem[115389] = 16'b0000000000000000;
	sram_mem[115390] = 16'b0000000000000000;
	sram_mem[115391] = 16'b0000000000000000;
	sram_mem[115392] = 16'b0000000000000000;
	sram_mem[115393] = 16'b0000000000000000;
	sram_mem[115394] = 16'b0000000000000000;
	sram_mem[115395] = 16'b0000000000000000;
	sram_mem[115396] = 16'b0000000000000000;
	sram_mem[115397] = 16'b0000000000000000;
	sram_mem[115398] = 16'b0000000000000000;
	sram_mem[115399] = 16'b0000000000000000;
	sram_mem[115400] = 16'b0000000000000000;
	sram_mem[115401] = 16'b0000000000000000;
	sram_mem[115402] = 16'b0000000000000000;
	sram_mem[115403] = 16'b0000000000000000;
	sram_mem[115404] = 16'b0000000000000000;
	sram_mem[115405] = 16'b0000000000000000;
	sram_mem[115406] = 16'b0000000000000000;
	sram_mem[115407] = 16'b0000000000000000;
	sram_mem[115408] = 16'b0000000000000000;
	sram_mem[115409] = 16'b0000000000000000;
	sram_mem[115410] = 16'b0000000000000000;
	sram_mem[115411] = 16'b0000000000000000;
	sram_mem[115412] = 16'b0000000000000000;
	sram_mem[115413] = 16'b0000000000000000;
	sram_mem[115414] = 16'b0000000000000000;
	sram_mem[115415] = 16'b0000000000000000;
	sram_mem[115416] = 16'b0000000000000000;
	sram_mem[115417] = 16'b0000000000000000;
	sram_mem[115418] = 16'b0000000000000000;
	sram_mem[115419] = 16'b0000000000000000;
	sram_mem[115420] = 16'b0000000000000000;
	sram_mem[115421] = 16'b0000000000000000;
	sram_mem[115422] = 16'b0000000000000000;
	sram_mem[115423] = 16'b0000000000000000;
	sram_mem[115424] = 16'b0000000000000000;
	sram_mem[115425] = 16'b0000000000000000;
	sram_mem[115426] = 16'b0000000000000000;
	sram_mem[115427] = 16'b0000000000000000;
	sram_mem[115428] = 16'b0000000000000000;
	sram_mem[115429] = 16'b0000000000000000;
	sram_mem[115430] = 16'b0000000000000000;
	sram_mem[115431] = 16'b0000000000000000;
	sram_mem[115432] = 16'b0000000000000000;
	sram_mem[115433] = 16'b0000000000000000;
	sram_mem[115434] = 16'b0000000000000000;
	sram_mem[115435] = 16'b0000000000000000;
	sram_mem[115436] = 16'b0000000000000000;
	sram_mem[115437] = 16'b0000000000000000;
	sram_mem[115438] = 16'b0000000000000000;
	sram_mem[115439] = 16'b0000000000000000;
	sram_mem[115440] = 16'b0000000000000000;
	sram_mem[115441] = 16'b0000000000000000;
	sram_mem[115442] = 16'b0000000000000000;
	sram_mem[115443] = 16'b0000000000000000;
	sram_mem[115444] = 16'b0000000000000000;
	sram_mem[115445] = 16'b0000000000000000;
	sram_mem[115446] = 16'b0000000000000000;
	sram_mem[115447] = 16'b0000000000000000;
	sram_mem[115448] = 16'b0000000000000000;
	sram_mem[115449] = 16'b0000000000000000;
	sram_mem[115450] = 16'b0000000000000000;
	sram_mem[115451] = 16'b0000000000000000;
	sram_mem[115452] = 16'b0000000000000000;
	sram_mem[115453] = 16'b0000000000000000;
	sram_mem[115454] = 16'b0000000000000000;
	sram_mem[115455] = 16'b0000000000000000;
	sram_mem[115456] = 16'b0000000000000000;
	sram_mem[115457] = 16'b0000000000000000;
	sram_mem[115458] = 16'b0000000000000000;
	sram_mem[115459] = 16'b0000000000000000;
	sram_mem[115460] = 16'b0000000000000000;
	sram_mem[115461] = 16'b0000000000000000;
	sram_mem[115462] = 16'b0000000000000000;
	sram_mem[115463] = 16'b0000000000000000;
	sram_mem[115464] = 16'b0000000000000000;
	sram_mem[115465] = 16'b0000000000000000;
	sram_mem[115466] = 16'b0000000000000000;
	sram_mem[115467] = 16'b0000000000000000;
	sram_mem[115468] = 16'b0000000000000000;
	sram_mem[115469] = 16'b0000000000000000;
	sram_mem[115470] = 16'b0000000000000000;
	sram_mem[115471] = 16'b0000000000000000;
	sram_mem[115472] = 16'b0000000000000000;
	sram_mem[115473] = 16'b0000000000000000;
	sram_mem[115474] = 16'b0000000000000000;
	sram_mem[115475] = 16'b0000000000000000;
	sram_mem[115476] = 16'b0000000000000000;
	sram_mem[115477] = 16'b0000000000000000;
	sram_mem[115478] = 16'b0000000000000000;
	sram_mem[115479] = 16'b0000000000000000;
	sram_mem[115480] = 16'b0000000000000000;
	sram_mem[115481] = 16'b0000000000000000;
	sram_mem[115482] = 16'b0000000000000000;
	sram_mem[115483] = 16'b0000000000000000;
	sram_mem[115484] = 16'b0000000000000000;
	sram_mem[115485] = 16'b0000000000000000;
	sram_mem[115486] = 16'b0000000000000000;
	sram_mem[115487] = 16'b0000000000000000;
	sram_mem[115488] = 16'b0000000000000000;
	sram_mem[115489] = 16'b0000000000000000;
	sram_mem[115490] = 16'b0000000000000000;
	sram_mem[115491] = 16'b0000000000000000;
	sram_mem[115492] = 16'b0000000000000000;
	sram_mem[115493] = 16'b0000000000000000;
	sram_mem[115494] = 16'b0000000000000000;
	sram_mem[115495] = 16'b0000000000000000;
	sram_mem[115496] = 16'b0000000000000000;
	sram_mem[115497] = 16'b0000000000000000;
	sram_mem[115498] = 16'b0000000000000000;
	sram_mem[115499] = 16'b0000000000000000;
	sram_mem[115500] = 16'b0000000000000000;
	sram_mem[115501] = 16'b0000000000000000;
	sram_mem[115502] = 16'b0000000000000000;
	sram_mem[115503] = 16'b0000000000000000;
	sram_mem[115504] = 16'b0000000000000000;
	sram_mem[115505] = 16'b0000000000000000;
	sram_mem[115506] = 16'b0000000000000000;
	sram_mem[115507] = 16'b0000000000000000;
	sram_mem[115508] = 16'b0000000000000000;
	sram_mem[115509] = 16'b0000000000000000;
	sram_mem[115510] = 16'b0000000000000000;
	sram_mem[115511] = 16'b0000000000000000;
	sram_mem[115512] = 16'b0000000000000000;
	sram_mem[115513] = 16'b0000000000000000;
	sram_mem[115514] = 16'b0000000000000000;
	sram_mem[115515] = 16'b0000000000000000;
	sram_mem[115516] = 16'b0000000000000000;
	sram_mem[115517] = 16'b0000000000000000;
	sram_mem[115518] = 16'b0000000000000000;
	sram_mem[115519] = 16'b0000000000000000;
	sram_mem[115520] = 16'b0000000000000000;
	sram_mem[115521] = 16'b0000000000000000;
	sram_mem[115522] = 16'b0000000000000000;
	sram_mem[115523] = 16'b0000000000000000;
	sram_mem[115524] = 16'b0000000000000000;
	sram_mem[115525] = 16'b0000000000000000;
	sram_mem[115526] = 16'b0000000000000000;
	sram_mem[115527] = 16'b0000000000000000;
	sram_mem[115528] = 16'b0000000000000000;
	sram_mem[115529] = 16'b0000000000000000;
	sram_mem[115530] = 16'b0000000000000000;
	sram_mem[115531] = 16'b0000000000000000;
	sram_mem[115532] = 16'b0000000000000000;
	sram_mem[115533] = 16'b0000000000000000;
	sram_mem[115534] = 16'b0000000000000000;
	sram_mem[115535] = 16'b0000000000000000;
	sram_mem[115536] = 16'b0000000000000000;
	sram_mem[115537] = 16'b0000000000000000;
	sram_mem[115538] = 16'b0000000000000000;
	sram_mem[115539] = 16'b0000000000000000;
	sram_mem[115540] = 16'b0000000000000000;
	sram_mem[115541] = 16'b0000000000000000;
	sram_mem[115542] = 16'b0000000000000000;
	sram_mem[115543] = 16'b0000000000000000;
	sram_mem[115544] = 16'b0000000000000000;
	sram_mem[115545] = 16'b0000000000000000;
	sram_mem[115546] = 16'b0000000000000000;
	sram_mem[115547] = 16'b0000000000000000;
	sram_mem[115548] = 16'b0000000000000000;
	sram_mem[115549] = 16'b0000000000000000;
	sram_mem[115550] = 16'b0000000000000000;
	sram_mem[115551] = 16'b0000000000000000;
	sram_mem[115552] = 16'b0000000000000000;
	sram_mem[115553] = 16'b0000000000000000;
	sram_mem[115554] = 16'b0000000000000000;
	sram_mem[115555] = 16'b0000000000000000;
	sram_mem[115556] = 16'b0000000000000000;
	sram_mem[115557] = 16'b0000000000000000;
	sram_mem[115558] = 16'b0000000000000000;
	sram_mem[115559] = 16'b0000000000000000;
	sram_mem[115560] = 16'b0000000000000000;
	sram_mem[115561] = 16'b0000000000000000;
	sram_mem[115562] = 16'b0000000000000000;
	sram_mem[115563] = 16'b0000000000000000;
	sram_mem[115564] = 16'b0000000000000000;
	sram_mem[115565] = 16'b0000000000000000;
	sram_mem[115566] = 16'b0000000000000000;
	sram_mem[115567] = 16'b0000000000000000;
	sram_mem[115568] = 16'b0000000000000000;
	sram_mem[115569] = 16'b0000000000000000;
	sram_mem[115570] = 16'b0000000000000000;
	sram_mem[115571] = 16'b0000000000000000;
	sram_mem[115572] = 16'b0000000000000000;
	sram_mem[115573] = 16'b0000000000000000;
	sram_mem[115574] = 16'b0000000000000000;
	sram_mem[115575] = 16'b0000000000000000;
	sram_mem[115576] = 16'b0000000000000000;
	sram_mem[115577] = 16'b0000000000000000;
	sram_mem[115578] = 16'b0000000000000000;
	sram_mem[115579] = 16'b0000000000000000;
	sram_mem[115580] = 16'b0000000000000000;
	sram_mem[115581] = 16'b0000000000000000;
	sram_mem[115582] = 16'b0000000000000000;
	sram_mem[115583] = 16'b0000000000000000;
	sram_mem[115584] = 16'b0000000000000000;
	sram_mem[115585] = 16'b0000000000000000;
	sram_mem[115586] = 16'b0000000000000000;
	sram_mem[115587] = 16'b0000000000000000;
	sram_mem[115588] = 16'b0000000000000000;
	sram_mem[115589] = 16'b0000000000000000;
	sram_mem[115590] = 16'b0000000000000000;
	sram_mem[115591] = 16'b0000000000000000;
	sram_mem[115592] = 16'b0000000000000000;
	sram_mem[115593] = 16'b0000000000000000;
	sram_mem[115594] = 16'b0000000000000000;
	sram_mem[115595] = 16'b0000000000000000;
	sram_mem[115596] = 16'b0000000000000000;
	sram_mem[115597] = 16'b0000000000000000;
	sram_mem[115598] = 16'b0000000000000000;
	sram_mem[115599] = 16'b0000000000000000;
	sram_mem[115600] = 16'b0000000000000000;
	sram_mem[115601] = 16'b0000000000000000;
	sram_mem[115602] = 16'b0000000000000000;
	sram_mem[115603] = 16'b0000000000000000;
	sram_mem[115604] = 16'b0000000000000000;
	sram_mem[115605] = 16'b0000000000000000;
	sram_mem[115606] = 16'b0000000000000000;
	sram_mem[115607] = 16'b0000000000000000;
	sram_mem[115608] = 16'b0000000000000000;
	sram_mem[115609] = 16'b0000000000000000;
	sram_mem[115610] = 16'b0000000000000000;
	sram_mem[115611] = 16'b0000000000000000;
	sram_mem[115612] = 16'b0000000000000000;
	sram_mem[115613] = 16'b0000000000000000;
	sram_mem[115614] = 16'b0000000000000000;
	sram_mem[115615] = 16'b0000000000000000;
	sram_mem[115616] = 16'b0000000000000000;
	sram_mem[115617] = 16'b0000000000000000;
	sram_mem[115618] = 16'b0000000000000000;
	sram_mem[115619] = 16'b0000000000000000;
	sram_mem[115620] = 16'b0000000000000000;
	sram_mem[115621] = 16'b0000000000000000;
	sram_mem[115622] = 16'b0000000000000000;
	sram_mem[115623] = 16'b0000000000000000;
	sram_mem[115624] = 16'b0000000000000000;
	sram_mem[115625] = 16'b0000000000000000;
	sram_mem[115626] = 16'b0000000000000000;
	sram_mem[115627] = 16'b0000000000000000;
	sram_mem[115628] = 16'b0000000000000000;
	sram_mem[115629] = 16'b0000000000000000;
	sram_mem[115630] = 16'b0000000000000000;
	sram_mem[115631] = 16'b0000000000000000;
	sram_mem[115632] = 16'b0000000000000000;
	sram_mem[115633] = 16'b0000000000000000;
	sram_mem[115634] = 16'b0000000000000000;
	sram_mem[115635] = 16'b0000000000000000;
	sram_mem[115636] = 16'b0000000000000000;
	sram_mem[115637] = 16'b0000000000000000;
	sram_mem[115638] = 16'b0000000000000000;
	sram_mem[115639] = 16'b0000000000000000;
	sram_mem[115640] = 16'b0000000000000000;
	sram_mem[115641] = 16'b0000000000000000;
	sram_mem[115642] = 16'b0000000000000000;
	sram_mem[115643] = 16'b0000000000000000;
	sram_mem[115644] = 16'b0000000000000000;
	sram_mem[115645] = 16'b0000000000000000;
	sram_mem[115646] = 16'b0000000000000000;
	sram_mem[115647] = 16'b0000000000000000;
	sram_mem[115648] = 16'b0000000000000000;
	sram_mem[115649] = 16'b0000000000000000;
	sram_mem[115650] = 16'b0000000000000000;
	sram_mem[115651] = 16'b0000000000000000;
	sram_mem[115652] = 16'b0000000000000000;
	sram_mem[115653] = 16'b0000000000000000;
	sram_mem[115654] = 16'b0000000000000000;
	sram_mem[115655] = 16'b0000000000000000;
	sram_mem[115656] = 16'b0000000000000000;
	sram_mem[115657] = 16'b0000000000000000;
	sram_mem[115658] = 16'b0000000000000000;
	sram_mem[115659] = 16'b0000000000000000;
	sram_mem[115660] = 16'b0000000000000000;
	sram_mem[115661] = 16'b0000000000000000;
	sram_mem[115662] = 16'b0000000000000000;
	sram_mem[115663] = 16'b0000000000000000;
	sram_mem[115664] = 16'b0000000000000000;
	sram_mem[115665] = 16'b0000000000000000;
	sram_mem[115666] = 16'b0000000000000000;
	sram_mem[115667] = 16'b0000000000000000;
	sram_mem[115668] = 16'b0000000000000000;
	sram_mem[115669] = 16'b0000000000000000;
	sram_mem[115670] = 16'b0000000000000000;
	sram_mem[115671] = 16'b0000000000000000;
	sram_mem[115672] = 16'b0000000000000000;
	sram_mem[115673] = 16'b0000000000000000;
	sram_mem[115674] = 16'b0000000000000000;
	sram_mem[115675] = 16'b0000000000000000;
	sram_mem[115676] = 16'b0000000000000000;
	sram_mem[115677] = 16'b0000000000000000;
	sram_mem[115678] = 16'b0000000000000000;
	sram_mem[115679] = 16'b0000000000000000;
	sram_mem[115680] = 16'b0000000000000000;
	sram_mem[115681] = 16'b0000000000000000;
	sram_mem[115682] = 16'b0000000000000000;
	sram_mem[115683] = 16'b0000000000000000;
	sram_mem[115684] = 16'b0000000000000000;
	sram_mem[115685] = 16'b0000000000000000;
	sram_mem[115686] = 16'b0000000000000000;
	sram_mem[115687] = 16'b0000000000000000;
	sram_mem[115688] = 16'b0000000000000000;
	sram_mem[115689] = 16'b0000000000000000;
	sram_mem[115690] = 16'b0000000000000000;
	sram_mem[115691] = 16'b0000000000000000;
	sram_mem[115692] = 16'b0000000000000000;
	sram_mem[115693] = 16'b0000000000000000;
	sram_mem[115694] = 16'b0000000000000000;
	sram_mem[115695] = 16'b0000000000000000;
	sram_mem[115696] = 16'b0000000000000000;
	sram_mem[115697] = 16'b0000000000000000;
	sram_mem[115698] = 16'b0000000000000000;
	sram_mem[115699] = 16'b0000000000000000;
	sram_mem[115700] = 16'b0000000000000000;
	sram_mem[115701] = 16'b0000000000000000;
	sram_mem[115702] = 16'b0000000000000000;
	sram_mem[115703] = 16'b0000000000000000;
	sram_mem[115704] = 16'b0000000000000000;
	sram_mem[115705] = 16'b0000000000000000;
	sram_mem[115706] = 16'b0000000000000000;
	sram_mem[115707] = 16'b0000000000000000;
	sram_mem[115708] = 16'b0000000000000000;
	sram_mem[115709] = 16'b0000000000000000;
	sram_mem[115710] = 16'b0000000000000000;
	sram_mem[115711] = 16'b0000000000000000;
	sram_mem[115712] = 16'b0000000000000000;
	sram_mem[115713] = 16'b0000000000000000;
	sram_mem[115714] = 16'b0000000000000000;
	sram_mem[115715] = 16'b0000000000000000;
	sram_mem[115716] = 16'b0000000000000000;
	sram_mem[115717] = 16'b0000000000000000;
	sram_mem[115718] = 16'b0000000000000000;
	sram_mem[115719] = 16'b0000000000000000;
	sram_mem[115720] = 16'b0000000000000000;
	sram_mem[115721] = 16'b0000000000000000;
	sram_mem[115722] = 16'b0000000000000000;
	sram_mem[115723] = 16'b0000000000000000;
	sram_mem[115724] = 16'b0000000000000000;
	sram_mem[115725] = 16'b0000000000000000;
	sram_mem[115726] = 16'b0000000000000000;
	sram_mem[115727] = 16'b0000000000000000;
	sram_mem[115728] = 16'b0000000000000000;
	sram_mem[115729] = 16'b0000000000000000;
	sram_mem[115730] = 16'b0000000000000000;
	sram_mem[115731] = 16'b0000000000000000;
	sram_mem[115732] = 16'b0000000000000000;
	sram_mem[115733] = 16'b0000000000000000;
	sram_mem[115734] = 16'b0000000000000000;
	sram_mem[115735] = 16'b0000000000000000;
	sram_mem[115736] = 16'b0000000000000000;
	sram_mem[115737] = 16'b0000000000000000;
	sram_mem[115738] = 16'b0000000000000000;
	sram_mem[115739] = 16'b0000000000000000;
	sram_mem[115740] = 16'b0000000000000000;
	sram_mem[115741] = 16'b0000000000000000;
	sram_mem[115742] = 16'b0000000000000000;
	sram_mem[115743] = 16'b0000000000000000;
	sram_mem[115744] = 16'b0000000000000000;
	sram_mem[115745] = 16'b0000000000000000;
	sram_mem[115746] = 16'b0000000000000000;
	sram_mem[115747] = 16'b0000000000000000;
	sram_mem[115748] = 16'b0000000000000000;
	sram_mem[115749] = 16'b0000000000000000;
	sram_mem[115750] = 16'b0000000000000000;
	sram_mem[115751] = 16'b0000000000000000;
	sram_mem[115752] = 16'b0000000000000000;
	sram_mem[115753] = 16'b0000000000000000;
	sram_mem[115754] = 16'b0000000000000000;
	sram_mem[115755] = 16'b0000000000000000;
	sram_mem[115756] = 16'b0000000000000000;
	sram_mem[115757] = 16'b0000000000000000;
	sram_mem[115758] = 16'b0000000000000000;
	sram_mem[115759] = 16'b0000000000000000;
	sram_mem[115760] = 16'b0000000000000000;
	sram_mem[115761] = 16'b0000000000000000;
	sram_mem[115762] = 16'b0000000000000000;
	sram_mem[115763] = 16'b0000000000000000;
	sram_mem[115764] = 16'b0000000000000000;
	sram_mem[115765] = 16'b0000000000000000;
	sram_mem[115766] = 16'b0000000000000000;
	sram_mem[115767] = 16'b0000000000000000;
	sram_mem[115768] = 16'b0000000000000000;
	sram_mem[115769] = 16'b0000000000000000;
	sram_mem[115770] = 16'b0000000000000000;
	sram_mem[115771] = 16'b0000000000000000;
	sram_mem[115772] = 16'b0000000000000000;
	sram_mem[115773] = 16'b0000000000000000;
	sram_mem[115774] = 16'b0000000000000000;
	sram_mem[115775] = 16'b0000000000000000;
	sram_mem[115776] = 16'b0000000000000000;
	sram_mem[115777] = 16'b0000000000000000;
	sram_mem[115778] = 16'b0000000000000000;
	sram_mem[115779] = 16'b0000000000000000;
	sram_mem[115780] = 16'b0000000000000000;
	sram_mem[115781] = 16'b0000000000000000;
	sram_mem[115782] = 16'b0000000000000000;
	sram_mem[115783] = 16'b0000000000000000;
	sram_mem[115784] = 16'b0000000000000000;
	sram_mem[115785] = 16'b0000000000000000;
	sram_mem[115786] = 16'b0000000000000000;
	sram_mem[115787] = 16'b0000000000000000;
	sram_mem[115788] = 16'b0000000000000000;
	sram_mem[115789] = 16'b0000000000000000;
	sram_mem[115790] = 16'b0000000000000000;
	sram_mem[115791] = 16'b0000000000000000;
	sram_mem[115792] = 16'b0000000000000000;
	sram_mem[115793] = 16'b0000000000000000;
	sram_mem[115794] = 16'b0000000000000000;
	sram_mem[115795] = 16'b0000000000000000;
	sram_mem[115796] = 16'b0000000000000000;
	sram_mem[115797] = 16'b0000000000000000;
	sram_mem[115798] = 16'b0000000000000000;
	sram_mem[115799] = 16'b0000000000000000;
	sram_mem[115800] = 16'b0000000000000000;
	sram_mem[115801] = 16'b0000000000000000;
	sram_mem[115802] = 16'b0000000000000000;
	sram_mem[115803] = 16'b0000000000000000;
	sram_mem[115804] = 16'b0000000000000000;
	sram_mem[115805] = 16'b0000000000000000;
	sram_mem[115806] = 16'b0000000000000000;
	sram_mem[115807] = 16'b0000000000000000;
	sram_mem[115808] = 16'b0000000000000000;
	sram_mem[115809] = 16'b0000000000000000;
	sram_mem[115810] = 16'b0000000000000000;
	sram_mem[115811] = 16'b0000000000000000;
	sram_mem[115812] = 16'b0000000000000000;
	sram_mem[115813] = 16'b0000000000000000;
	sram_mem[115814] = 16'b0000000000000000;
	sram_mem[115815] = 16'b0000000000000000;
	sram_mem[115816] = 16'b0000000000000000;
	sram_mem[115817] = 16'b0000000000000000;
	sram_mem[115818] = 16'b0000000000000000;
	sram_mem[115819] = 16'b0000000000000000;
	sram_mem[115820] = 16'b0000000000000000;
	sram_mem[115821] = 16'b0000000000000000;
	sram_mem[115822] = 16'b0000000000000000;
	sram_mem[115823] = 16'b0000000000000000;
	sram_mem[115824] = 16'b0000000000000000;
	sram_mem[115825] = 16'b0000000000000000;
	sram_mem[115826] = 16'b0000000000000000;
	sram_mem[115827] = 16'b0000000000000000;
	sram_mem[115828] = 16'b0000000000000000;
	sram_mem[115829] = 16'b0000000000000000;
	sram_mem[115830] = 16'b0000000000000000;
	sram_mem[115831] = 16'b0000000000000000;
	sram_mem[115832] = 16'b0000000000000000;
	sram_mem[115833] = 16'b0000000000000000;
	sram_mem[115834] = 16'b0000000000000000;
	sram_mem[115835] = 16'b0000000000000000;
	sram_mem[115836] = 16'b0000000000000000;
	sram_mem[115837] = 16'b0000000000000000;
	sram_mem[115838] = 16'b0000000000000000;
	sram_mem[115839] = 16'b0000000000000000;
	sram_mem[115840] = 16'b0000000000000000;
	sram_mem[115841] = 16'b0000000000000000;
	sram_mem[115842] = 16'b0000000000000000;
	sram_mem[115843] = 16'b0000000000000000;
	sram_mem[115844] = 16'b0000000000000000;
	sram_mem[115845] = 16'b0000000000000000;
	sram_mem[115846] = 16'b0000000000000000;
	sram_mem[115847] = 16'b0000000000000000;
	sram_mem[115848] = 16'b0000000000000000;
	sram_mem[115849] = 16'b0000000000000000;
	sram_mem[115850] = 16'b0000000000000000;
	sram_mem[115851] = 16'b0000000000000000;
	sram_mem[115852] = 16'b0000000000000000;
	sram_mem[115853] = 16'b0000000000000000;
	sram_mem[115854] = 16'b0000000000000000;
	sram_mem[115855] = 16'b0000000000000000;
	sram_mem[115856] = 16'b0000000000000000;
	sram_mem[115857] = 16'b0000000000000000;
	sram_mem[115858] = 16'b0000000000000000;
	sram_mem[115859] = 16'b0000000000000000;
	sram_mem[115860] = 16'b0000000000000000;
	sram_mem[115861] = 16'b0000000000000000;
	sram_mem[115862] = 16'b0000000000000000;
	sram_mem[115863] = 16'b0000000000000000;
	sram_mem[115864] = 16'b0000000000000000;
	sram_mem[115865] = 16'b0000000000000000;
	sram_mem[115866] = 16'b0000000000000000;
	sram_mem[115867] = 16'b0000000000000000;
	sram_mem[115868] = 16'b0000000000000000;
	sram_mem[115869] = 16'b0000000000000000;
	sram_mem[115870] = 16'b0000000000000000;
	sram_mem[115871] = 16'b0000000000000000;
	sram_mem[115872] = 16'b0000000000000000;
	sram_mem[115873] = 16'b0000000000000000;
	sram_mem[115874] = 16'b0000000000000000;
	sram_mem[115875] = 16'b0000000000000000;
	sram_mem[115876] = 16'b0000000000000000;
	sram_mem[115877] = 16'b0000000000000000;
	sram_mem[115878] = 16'b0000000000000000;
	sram_mem[115879] = 16'b0000000000000000;
	sram_mem[115880] = 16'b0000000000000000;
	sram_mem[115881] = 16'b0000000000000000;
	sram_mem[115882] = 16'b0000000000000000;
	sram_mem[115883] = 16'b0000000000000000;
	sram_mem[115884] = 16'b0000000000000000;
	sram_mem[115885] = 16'b0000000000000000;
	sram_mem[115886] = 16'b0000000000000000;
	sram_mem[115887] = 16'b0000000000000000;
	sram_mem[115888] = 16'b0000000000000000;
	sram_mem[115889] = 16'b0000000000000000;
	sram_mem[115890] = 16'b0000000000000000;
	sram_mem[115891] = 16'b0000000000000000;
	sram_mem[115892] = 16'b0000000000000000;
	sram_mem[115893] = 16'b0000000000000000;
	sram_mem[115894] = 16'b0000000000000000;
	sram_mem[115895] = 16'b0000000000000000;
	sram_mem[115896] = 16'b0000000000000000;
	sram_mem[115897] = 16'b0000000000000000;
	sram_mem[115898] = 16'b0000000000000000;
	sram_mem[115899] = 16'b0000000000000000;
	sram_mem[115900] = 16'b0000000000000000;
	sram_mem[115901] = 16'b0000000000000000;
	sram_mem[115902] = 16'b0000000000000000;
	sram_mem[115903] = 16'b0000000000000000;
	sram_mem[115904] = 16'b0000000000000000;
	sram_mem[115905] = 16'b0000000000000000;
	sram_mem[115906] = 16'b0000000000000000;
	sram_mem[115907] = 16'b0000000000000000;
	sram_mem[115908] = 16'b0000000000000000;
	sram_mem[115909] = 16'b0000000000000000;
	sram_mem[115910] = 16'b0000000000000000;
	sram_mem[115911] = 16'b0000000000000000;
	sram_mem[115912] = 16'b0000000000000000;
	sram_mem[115913] = 16'b0000000000000000;
	sram_mem[115914] = 16'b0000000000000000;
	sram_mem[115915] = 16'b0000000000000000;
	sram_mem[115916] = 16'b0000000000000000;
	sram_mem[115917] = 16'b0000000000000000;
	sram_mem[115918] = 16'b0000000000000000;
	sram_mem[115919] = 16'b0000000000000000;
	sram_mem[115920] = 16'b0000000000000000;
	sram_mem[115921] = 16'b0000000000000000;
	sram_mem[115922] = 16'b0000000000000000;
	sram_mem[115923] = 16'b0000000000000000;
	sram_mem[115924] = 16'b0000000000000000;
	sram_mem[115925] = 16'b0000000000000000;
	sram_mem[115926] = 16'b0000000000000000;
	sram_mem[115927] = 16'b0000000000000000;
	sram_mem[115928] = 16'b0000000000000000;
	sram_mem[115929] = 16'b0000000000000000;
	sram_mem[115930] = 16'b0000000000000000;
	sram_mem[115931] = 16'b0000000000000000;
	sram_mem[115932] = 16'b0000000000000000;
	sram_mem[115933] = 16'b0000000000000000;
	sram_mem[115934] = 16'b0000000000000000;
	sram_mem[115935] = 16'b0000000000000000;
	sram_mem[115936] = 16'b0000000000000000;
	sram_mem[115937] = 16'b0000000000000000;
	sram_mem[115938] = 16'b0000000000000000;
	sram_mem[115939] = 16'b0000000000000000;
	sram_mem[115940] = 16'b0000000000000000;
	sram_mem[115941] = 16'b0000000000000000;
	sram_mem[115942] = 16'b0000000000000000;
	sram_mem[115943] = 16'b0000000000000000;
	sram_mem[115944] = 16'b0000000000000000;
	sram_mem[115945] = 16'b0000000000000000;
	sram_mem[115946] = 16'b0000000000000000;
	sram_mem[115947] = 16'b0000000000000000;
	sram_mem[115948] = 16'b0000000000000000;
	sram_mem[115949] = 16'b0000000000000000;
	sram_mem[115950] = 16'b0000000000000000;
	sram_mem[115951] = 16'b0000000000000000;
	sram_mem[115952] = 16'b0000000000000000;
	sram_mem[115953] = 16'b0000000000000000;
	sram_mem[115954] = 16'b0000000000000000;
	sram_mem[115955] = 16'b0000000000000000;
	sram_mem[115956] = 16'b0000000000000000;
	sram_mem[115957] = 16'b0000000000000000;
	sram_mem[115958] = 16'b0000000000000000;
	sram_mem[115959] = 16'b0000000000000000;
	sram_mem[115960] = 16'b0000000000000000;
	sram_mem[115961] = 16'b0000000000000000;
	sram_mem[115962] = 16'b0000000000000000;
	sram_mem[115963] = 16'b0000000000000000;
	sram_mem[115964] = 16'b0000000000000000;
	sram_mem[115965] = 16'b0000000000000000;
	sram_mem[115966] = 16'b0000000000000000;
	sram_mem[115967] = 16'b0000000000000000;
	sram_mem[115968] = 16'b0000000000000000;
	sram_mem[115969] = 16'b0000000000000000;
	sram_mem[115970] = 16'b0000000000000000;
	sram_mem[115971] = 16'b0000000000000000;
	sram_mem[115972] = 16'b0000000000000000;
	sram_mem[115973] = 16'b0000000000000000;
	sram_mem[115974] = 16'b0000000000000000;
	sram_mem[115975] = 16'b0000000000000000;
	sram_mem[115976] = 16'b0000000000000000;
	sram_mem[115977] = 16'b0000000000000000;
	sram_mem[115978] = 16'b0000000000000000;
	sram_mem[115979] = 16'b0000000000000000;
	sram_mem[115980] = 16'b0000000000000000;
	sram_mem[115981] = 16'b0000000000000000;
	sram_mem[115982] = 16'b0000000000000000;
	sram_mem[115983] = 16'b0000000000000000;
	sram_mem[115984] = 16'b0000000000000000;
	sram_mem[115985] = 16'b0000000000000000;
	sram_mem[115986] = 16'b0000000000000000;
	sram_mem[115987] = 16'b0000000000000000;
	sram_mem[115988] = 16'b0000000000000000;
	sram_mem[115989] = 16'b0000000000000000;
	sram_mem[115990] = 16'b0000000000000000;
	sram_mem[115991] = 16'b0000000000000000;
	sram_mem[115992] = 16'b0000000000000000;
	sram_mem[115993] = 16'b0000000000000000;
	sram_mem[115994] = 16'b0000000000000000;
	sram_mem[115995] = 16'b0000000000000000;
	sram_mem[115996] = 16'b0000000000000000;
	sram_mem[115997] = 16'b0000000000000000;
	sram_mem[115998] = 16'b0000000000000000;
	sram_mem[115999] = 16'b0000000000000000;
	sram_mem[116000] = 16'b0000000000000000;
	sram_mem[116001] = 16'b0000000000000000;
	sram_mem[116002] = 16'b0000000000000000;
	sram_mem[116003] = 16'b0000000000000000;
	sram_mem[116004] = 16'b0000000000000000;
	sram_mem[116005] = 16'b0000000000000000;
	sram_mem[116006] = 16'b0000000000000000;
	sram_mem[116007] = 16'b0000000000000000;
	sram_mem[116008] = 16'b0000000000000000;
	sram_mem[116009] = 16'b0000000000000000;
	sram_mem[116010] = 16'b0000000000000000;
	sram_mem[116011] = 16'b0000000000000000;
	sram_mem[116012] = 16'b0000000000000000;
	sram_mem[116013] = 16'b0000000000000000;
	sram_mem[116014] = 16'b0000000000000000;
	sram_mem[116015] = 16'b0000000000000000;
	sram_mem[116016] = 16'b0000000000000000;
	sram_mem[116017] = 16'b0000000000000000;
	sram_mem[116018] = 16'b0000000000000000;
	sram_mem[116019] = 16'b0000000000000000;
	sram_mem[116020] = 16'b0000000000000000;
	sram_mem[116021] = 16'b0000000000000000;
	sram_mem[116022] = 16'b0000000000000000;
	sram_mem[116023] = 16'b0000000000000000;
	sram_mem[116024] = 16'b0000000000000000;
	sram_mem[116025] = 16'b0000000000000000;
	sram_mem[116026] = 16'b0000000000000000;
	sram_mem[116027] = 16'b0000000000000000;
	sram_mem[116028] = 16'b0000000000000000;
	sram_mem[116029] = 16'b0000000000000000;
	sram_mem[116030] = 16'b0000000000000000;
	sram_mem[116031] = 16'b0000000000000000;
	sram_mem[116032] = 16'b0000000000000000;
	sram_mem[116033] = 16'b0000000000000000;
	sram_mem[116034] = 16'b0000000000000000;
	sram_mem[116035] = 16'b0000000000000000;
	sram_mem[116036] = 16'b0000000000000000;
	sram_mem[116037] = 16'b0000000000000000;
	sram_mem[116038] = 16'b0000000000000000;
	sram_mem[116039] = 16'b0000000000000000;
	sram_mem[116040] = 16'b0000000000000000;
	sram_mem[116041] = 16'b0000000000000000;
	sram_mem[116042] = 16'b0000000000000000;
	sram_mem[116043] = 16'b0000000000000000;
	sram_mem[116044] = 16'b0000000000000000;
	sram_mem[116045] = 16'b0000000000000000;
	sram_mem[116046] = 16'b0000000000000000;
	sram_mem[116047] = 16'b0000000000000000;
	sram_mem[116048] = 16'b0000000000000000;
	sram_mem[116049] = 16'b0000000000000000;
	sram_mem[116050] = 16'b0000000000000000;
	sram_mem[116051] = 16'b0000000000000000;
	sram_mem[116052] = 16'b0000000000000000;
	sram_mem[116053] = 16'b0000000000000000;
	sram_mem[116054] = 16'b0000000000000000;
	sram_mem[116055] = 16'b0000000000000000;
	sram_mem[116056] = 16'b0000000000000000;
	sram_mem[116057] = 16'b0000000000000000;
	sram_mem[116058] = 16'b0000000000000000;
	sram_mem[116059] = 16'b0000000000000000;
	sram_mem[116060] = 16'b0000000000000000;
	sram_mem[116061] = 16'b0000000000000000;
	sram_mem[116062] = 16'b0000000000000000;
	sram_mem[116063] = 16'b0000000000000000;
	sram_mem[116064] = 16'b0000000000000000;
	sram_mem[116065] = 16'b0000000000000000;
	sram_mem[116066] = 16'b0000000000000000;
	sram_mem[116067] = 16'b0000000000000000;
	sram_mem[116068] = 16'b0000000000000000;
	sram_mem[116069] = 16'b0000000000000000;
	sram_mem[116070] = 16'b0000000000000000;
	sram_mem[116071] = 16'b0000000000000000;
	sram_mem[116072] = 16'b0000000000000000;
	sram_mem[116073] = 16'b0000000000000000;
	sram_mem[116074] = 16'b0000000000000000;
	sram_mem[116075] = 16'b0000000000000000;
	sram_mem[116076] = 16'b0000000000000000;
	sram_mem[116077] = 16'b0000000000000000;
	sram_mem[116078] = 16'b0000000000000000;
	sram_mem[116079] = 16'b0000000000000000;
	sram_mem[116080] = 16'b0000000000000000;
	sram_mem[116081] = 16'b0000000000000000;
	sram_mem[116082] = 16'b0000000000000000;
	sram_mem[116083] = 16'b0000000000000000;
	sram_mem[116084] = 16'b0000000000000000;
	sram_mem[116085] = 16'b0000000000000000;
	sram_mem[116086] = 16'b0000000000000000;
	sram_mem[116087] = 16'b0000000000000000;
	sram_mem[116088] = 16'b0000000000000000;
	sram_mem[116089] = 16'b0000000000000000;
	sram_mem[116090] = 16'b0000000000000000;
	sram_mem[116091] = 16'b0000000000000000;
	sram_mem[116092] = 16'b0000000000000000;
	sram_mem[116093] = 16'b0000000000000000;
	sram_mem[116094] = 16'b0000000000000000;
	sram_mem[116095] = 16'b0000000000000000;
	sram_mem[116096] = 16'b0000000000000000;
	sram_mem[116097] = 16'b0000000000000000;
	sram_mem[116098] = 16'b0000000000000000;
	sram_mem[116099] = 16'b0000000000000000;
	sram_mem[116100] = 16'b0000000000000000;
	sram_mem[116101] = 16'b0000000000000000;
	sram_mem[116102] = 16'b0000000000000000;
	sram_mem[116103] = 16'b0000000000000000;
	sram_mem[116104] = 16'b0000000000000000;
	sram_mem[116105] = 16'b0000000000000000;
	sram_mem[116106] = 16'b0000000000000000;
	sram_mem[116107] = 16'b0000000000000000;
	sram_mem[116108] = 16'b0000000000000000;
	sram_mem[116109] = 16'b0000000000000000;
	sram_mem[116110] = 16'b0000000000000000;
	sram_mem[116111] = 16'b0000000000000000;
	sram_mem[116112] = 16'b0000000000000000;
	sram_mem[116113] = 16'b0000000000000000;
	sram_mem[116114] = 16'b0000000000000000;
	sram_mem[116115] = 16'b0000000000000000;
	sram_mem[116116] = 16'b0000000000000000;
	sram_mem[116117] = 16'b0000000000000000;
	sram_mem[116118] = 16'b0000000000000000;
	sram_mem[116119] = 16'b0000000000000000;
	sram_mem[116120] = 16'b0000000000000000;
	sram_mem[116121] = 16'b0000000000000000;
	sram_mem[116122] = 16'b0000000000000000;
	sram_mem[116123] = 16'b0000000000000000;
	sram_mem[116124] = 16'b0000000000000000;
	sram_mem[116125] = 16'b0000000000000000;
	sram_mem[116126] = 16'b0000000000000000;
	sram_mem[116127] = 16'b0000000000000000;
	sram_mem[116128] = 16'b0000000000000000;
	sram_mem[116129] = 16'b0000000000000000;
	sram_mem[116130] = 16'b0000000000000000;
	sram_mem[116131] = 16'b0000000000000000;
	sram_mem[116132] = 16'b0000000000000000;
	sram_mem[116133] = 16'b0000000000000000;
	sram_mem[116134] = 16'b0000000000000000;
	sram_mem[116135] = 16'b0000000000000000;
	sram_mem[116136] = 16'b0000000000000000;
	sram_mem[116137] = 16'b0000000000000000;
	sram_mem[116138] = 16'b0000000000000000;
	sram_mem[116139] = 16'b0000000000000000;
	sram_mem[116140] = 16'b0000000000000000;
	sram_mem[116141] = 16'b0000000000000000;
	sram_mem[116142] = 16'b0000000000000000;
	sram_mem[116143] = 16'b0000000000000000;
	sram_mem[116144] = 16'b0000000000000000;
	sram_mem[116145] = 16'b0000000000000000;
	sram_mem[116146] = 16'b0000000000000000;
	sram_mem[116147] = 16'b0000000000000000;
	sram_mem[116148] = 16'b0000000000000000;
	sram_mem[116149] = 16'b0000000000000000;
	sram_mem[116150] = 16'b0000000000000000;
	sram_mem[116151] = 16'b0000000000000000;
	sram_mem[116152] = 16'b0000000000000000;
	sram_mem[116153] = 16'b0000000000000000;
	sram_mem[116154] = 16'b0000000000000000;
	sram_mem[116155] = 16'b0000000000000000;
	sram_mem[116156] = 16'b0000000000000000;
	sram_mem[116157] = 16'b0000000000000000;
	sram_mem[116158] = 16'b0000000000000000;
	sram_mem[116159] = 16'b0000000000000000;
	sram_mem[116160] = 16'b0000000000000000;
	sram_mem[116161] = 16'b0000000000000000;
	sram_mem[116162] = 16'b0000000000000000;
	sram_mem[116163] = 16'b0000000000000000;
	sram_mem[116164] = 16'b0000000000000000;
	sram_mem[116165] = 16'b0000000000000000;
	sram_mem[116166] = 16'b0000000000000000;
	sram_mem[116167] = 16'b0000000000000000;
	sram_mem[116168] = 16'b0000000000000000;
	sram_mem[116169] = 16'b0000000000000000;
	sram_mem[116170] = 16'b0000000000000000;
	sram_mem[116171] = 16'b0000000000000000;
	sram_mem[116172] = 16'b0000000000000000;
	sram_mem[116173] = 16'b0000000000000000;
	sram_mem[116174] = 16'b0000000000000000;
	sram_mem[116175] = 16'b0000000000000000;
	sram_mem[116176] = 16'b0000000000000000;
	sram_mem[116177] = 16'b0000000000000000;
	sram_mem[116178] = 16'b0000000000000000;
	sram_mem[116179] = 16'b0000000000000000;
	sram_mem[116180] = 16'b0000000000000000;
	sram_mem[116181] = 16'b0000000000000000;
	sram_mem[116182] = 16'b0000000000000000;
	sram_mem[116183] = 16'b0000000000000000;
	sram_mem[116184] = 16'b0000000000000000;
	sram_mem[116185] = 16'b0000000000000000;
	sram_mem[116186] = 16'b0000000000000000;
	sram_mem[116187] = 16'b0000000000000000;
	sram_mem[116188] = 16'b0000000000000000;
	sram_mem[116189] = 16'b0000000000000000;
	sram_mem[116190] = 16'b0000000000000000;
	sram_mem[116191] = 16'b0000000000000000;
	sram_mem[116192] = 16'b0000000000000000;
	sram_mem[116193] = 16'b0000000000000000;
	sram_mem[116194] = 16'b0000000000000000;
	sram_mem[116195] = 16'b0000000000000000;
	sram_mem[116196] = 16'b0000000000000000;
	sram_mem[116197] = 16'b0000000000000000;
	sram_mem[116198] = 16'b0000000000000000;
	sram_mem[116199] = 16'b0000000000000000;
	sram_mem[116200] = 16'b0000000000000000;
	sram_mem[116201] = 16'b0000000000000000;
	sram_mem[116202] = 16'b0000000000000000;
	sram_mem[116203] = 16'b0000000000000000;
	sram_mem[116204] = 16'b0000000000000000;
	sram_mem[116205] = 16'b0000000000000000;
	sram_mem[116206] = 16'b0000000000000000;
	sram_mem[116207] = 16'b0000000000000000;
	sram_mem[116208] = 16'b0000000000000000;
	sram_mem[116209] = 16'b0000000000000000;
	sram_mem[116210] = 16'b0000000000000000;
	sram_mem[116211] = 16'b0000000000000000;
	sram_mem[116212] = 16'b0000000000000000;
	sram_mem[116213] = 16'b0000000000000000;
	sram_mem[116214] = 16'b0000000000000000;
	sram_mem[116215] = 16'b0000000000000000;
	sram_mem[116216] = 16'b0000000000000000;
	sram_mem[116217] = 16'b0000000000000000;
	sram_mem[116218] = 16'b0000000000000000;
	sram_mem[116219] = 16'b0000000000000000;
	sram_mem[116220] = 16'b0000000000000000;
	sram_mem[116221] = 16'b0000000000000000;
	sram_mem[116222] = 16'b0000000000000000;
	sram_mem[116223] = 16'b0000000000000000;
	sram_mem[116224] = 16'b0000000000000000;
	sram_mem[116225] = 16'b0000000000000000;
	sram_mem[116226] = 16'b0000000000000000;
	sram_mem[116227] = 16'b0000000000000000;
	sram_mem[116228] = 16'b0000000000000000;
	sram_mem[116229] = 16'b0000000000000000;
	sram_mem[116230] = 16'b0000000000000000;
	sram_mem[116231] = 16'b0000000000000000;
	sram_mem[116232] = 16'b0000000000000000;
	sram_mem[116233] = 16'b0000000000000000;
	sram_mem[116234] = 16'b0000000000000000;
	sram_mem[116235] = 16'b0000000000000000;
	sram_mem[116236] = 16'b0000000000000000;
	sram_mem[116237] = 16'b0000000000000000;
	sram_mem[116238] = 16'b0000000000000000;
	sram_mem[116239] = 16'b0000000000000000;
	sram_mem[116240] = 16'b0000000000000000;
	sram_mem[116241] = 16'b0000000000000000;
	sram_mem[116242] = 16'b0000000000000000;
	sram_mem[116243] = 16'b0000000000000000;
	sram_mem[116244] = 16'b0000000000000000;
	sram_mem[116245] = 16'b0000000000000000;
	sram_mem[116246] = 16'b0000000000000000;
	sram_mem[116247] = 16'b0000000000000000;
	sram_mem[116248] = 16'b0000000000000000;
	sram_mem[116249] = 16'b0000000000000000;
	sram_mem[116250] = 16'b0000000000000000;
	sram_mem[116251] = 16'b0000000000000000;
	sram_mem[116252] = 16'b0000000000000000;
	sram_mem[116253] = 16'b0000000000000000;
	sram_mem[116254] = 16'b0000000000000000;
	sram_mem[116255] = 16'b0000000000000000;
	sram_mem[116256] = 16'b0000000000000000;
	sram_mem[116257] = 16'b0000000000000000;
	sram_mem[116258] = 16'b0000000000000000;
	sram_mem[116259] = 16'b0000000000000000;
	sram_mem[116260] = 16'b0000000000000000;
	sram_mem[116261] = 16'b0000000000000000;
	sram_mem[116262] = 16'b0000000000000000;
	sram_mem[116263] = 16'b0000000000000000;
	sram_mem[116264] = 16'b0000000000000000;
	sram_mem[116265] = 16'b0000000000000000;
	sram_mem[116266] = 16'b0000000000000000;
	sram_mem[116267] = 16'b0000000000000000;
	sram_mem[116268] = 16'b0000000000000000;
	sram_mem[116269] = 16'b0000000000000000;
	sram_mem[116270] = 16'b0000000000000000;
	sram_mem[116271] = 16'b0000000000000000;
	sram_mem[116272] = 16'b0000000000000000;
	sram_mem[116273] = 16'b0000000000000000;
	sram_mem[116274] = 16'b0000000000000000;
	sram_mem[116275] = 16'b0000000000000000;
	sram_mem[116276] = 16'b0000000000000000;
	sram_mem[116277] = 16'b0000000000000000;
	sram_mem[116278] = 16'b0000000000000000;
	sram_mem[116279] = 16'b0000000000000000;
	sram_mem[116280] = 16'b0000000000000000;
	sram_mem[116281] = 16'b0000000000000000;
	sram_mem[116282] = 16'b0000000000000000;
	sram_mem[116283] = 16'b0000000000000000;
	sram_mem[116284] = 16'b0000000000000000;
	sram_mem[116285] = 16'b0000000000000000;
	sram_mem[116286] = 16'b0000000000000000;
	sram_mem[116287] = 16'b0000000000000000;
	sram_mem[116288] = 16'b0000000000000000;
	sram_mem[116289] = 16'b0000000000000000;
	sram_mem[116290] = 16'b0000000000000000;
	sram_mem[116291] = 16'b0000000000000000;
	sram_mem[116292] = 16'b0000000000000000;
	sram_mem[116293] = 16'b0000000000000000;
	sram_mem[116294] = 16'b0000000000000000;
	sram_mem[116295] = 16'b0000000000000000;
	sram_mem[116296] = 16'b0000000000000000;
	sram_mem[116297] = 16'b0000000000000000;
	sram_mem[116298] = 16'b0000000000000000;
	sram_mem[116299] = 16'b0000000000000000;
	sram_mem[116300] = 16'b0000000000000000;
	sram_mem[116301] = 16'b0000000000000000;
	sram_mem[116302] = 16'b0000000000000000;
	sram_mem[116303] = 16'b0000000000000000;
	sram_mem[116304] = 16'b0000000000000000;
	sram_mem[116305] = 16'b0000000000000000;
	sram_mem[116306] = 16'b0000000000000000;
	sram_mem[116307] = 16'b0000000000000000;
	sram_mem[116308] = 16'b0000000000000000;
	sram_mem[116309] = 16'b0000000000000000;
	sram_mem[116310] = 16'b0000000000000000;
	sram_mem[116311] = 16'b0000000000000000;
	sram_mem[116312] = 16'b0000000000000000;
	sram_mem[116313] = 16'b0000000000000000;
	sram_mem[116314] = 16'b0000000000000000;
	sram_mem[116315] = 16'b0000000000000000;
	sram_mem[116316] = 16'b0000000000000000;
	sram_mem[116317] = 16'b0000000000000000;
	sram_mem[116318] = 16'b0000000000000000;
	sram_mem[116319] = 16'b0000000000000000;
	sram_mem[116320] = 16'b0000000000000000;
	sram_mem[116321] = 16'b0000000000000000;
	sram_mem[116322] = 16'b0000000000000000;
	sram_mem[116323] = 16'b0000000000000000;
	sram_mem[116324] = 16'b0000000000000000;
	sram_mem[116325] = 16'b0000000000000000;
	sram_mem[116326] = 16'b0000000000000000;
	sram_mem[116327] = 16'b0000000000000000;
	sram_mem[116328] = 16'b0000000000000000;
	sram_mem[116329] = 16'b0000000000000000;
	sram_mem[116330] = 16'b0000000000000000;
	sram_mem[116331] = 16'b0000000000000000;
	sram_mem[116332] = 16'b0000000000000000;
	sram_mem[116333] = 16'b0000000000000000;
	sram_mem[116334] = 16'b0000000000000000;
	sram_mem[116335] = 16'b0000000000000000;
	sram_mem[116336] = 16'b0000000000000000;
	sram_mem[116337] = 16'b0000000000000000;
	sram_mem[116338] = 16'b0000000000000000;
	sram_mem[116339] = 16'b0000000000000000;
	sram_mem[116340] = 16'b0000000000000000;
	sram_mem[116341] = 16'b0000000000000000;
	sram_mem[116342] = 16'b0000000000000000;
	sram_mem[116343] = 16'b0000000000000000;
	sram_mem[116344] = 16'b0000000000000000;
	sram_mem[116345] = 16'b0000000000000000;
	sram_mem[116346] = 16'b0000000000000000;
	sram_mem[116347] = 16'b0000000000000000;
	sram_mem[116348] = 16'b0000000000000000;
	sram_mem[116349] = 16'b0000000000000000;
	sram_mem[116350] = 16'b0000000000000000;
	sram_mem[116351] = 16'b0000000000000000;
	sram_mem[116352] = 16'b0000000000000000;
	sram_mem[116353] = 16'b0000000000000000;
	sram_mem[116354] = 16'b0000000000000000;
	sram_mem[116355] = 16'b0000000000000000;
	sram_mem[116356] = 16'b0000000000000000;
	sram_mem[116357] = 16'b0000000000000000;
	sram_mem[116358] = 16'b0000000000000000;
	sram_mem[116359] = 16'b0000000000000000;
	sram_mem[116360] = 16'b0000000000000000;
	sram_mem[116361] = 16'b0000000000000000;
	sram_mem[116362] = 16'b0000000000000000;
	sram_mem[116363] = 16'b0000000000000000;
	sram_mem[116364] = 16'b0000000000000000;
	sram_mem[116365] = 16'b0000000000000000;
	sram_mem[116366] = 16'b0000000000000000;
	sram_mem[116367] = 16'b0000000000000000;
	sram_mem[116368] = 16'b0000000000000000;
	sram_mem[116369] = 16'b0000000000000000;
	sram_mem[116370] = 16'b0000000000000000;
	sram_mem[116371] = 16'b0000000000000000;
	sram_mem[116372] = 16'b0000000000000000;
	sram_mem[116373] = 16'b0000000000000000;
	sram_mem[116374] = 16'b0000000000000000;
	sram_mem[116375] = 16'b0000000000000000;
	sram_mem[116376] = 16'b0000000000000000;
	sram_mem[116377] = 16'b0000000000000000;
	sram_mem[116378] = 16'b0000000000000000;
	sram_mem[116379] = 16'b0000000000000000;
	sram_mem[116380] = 16'b0000000000000000;
	sram_mem[116381] = 16'b0000000000000000;
	sram_mem[116382] = 16'b0000000000000000;
	sram_mem[116383] = 16'b0000000000000000;
	sram_mem[116384] = 16'b0000000000000000;
	sram_mem[116385] = 16'b0000000000000000;
	sram_mem[116386] = 16'b0000000000000000;
	sram_mem[116387] = 16'b0000000000000000;
	sram_mem[116388] = 16'b0000000000000000;
	sram_mem[116389] = 16'b0000000000000000;
	sram_mem[116390] = 16'b0000000000000000;
	sram_mem[116391] = 16'b0000000000000000;
	sram_mem[116392] = 16'b0000000000000000;
	sram_mem[116393] = 16'b0000000000000000;
	sram_mem[116394] = 16'b0000000000000000;
	sram_mem[116395] = 16'b0000000000000000;
	sram_mem[116396] = 16'b0000000000000000;
	sram_mem[116397] = 16'b0000000000000000;
	sram_mem[116398] = 16'b0000000000000000;
	sram_mem[116399] = 16'b0000000000000000;
	sram_mem[116400] = 16'b0000000000000000;
	sram_mem[116401] = 16'b0000000000000000;
	sram_mem[116402] = 16'b0000000000000000;
	sram_mem[116403] = 16'b0000000000000000;
	sram_mem[116404] = 16'b0000000000000000;
	sram_mem[116405] = 16'b0000000000000000;
	sram_mem[116406] = 16'b0000000000000000;
	sram_mem[116407] = 16'b0000000000000000;
	sram_mem[116408] = 16'b0000000000000000;
	sram_mem[116409] = 16'b0000000000000000;
	sram_mem[116410] = 16'b0000000000000000;
	sram_mem[116411] = 16'b0000000000000000;
	sram_mem[116412] = 16'b0000000000000000;
	sram_mem[116413] = 16'b0000000000000000;
	sram_mem[116414] = 16'b0000000000000000;
	sram_mem[116415] = 16'b0000000000000000;
	sram_mem[116416] = 16'b0000000000000000;
	sram_mem[116417] = 16'b0000000000000000;
	sram_mem[116418] = 16'b0000000000000000;
	sram_mem[116419] = 16'b0000000000000000;
	sram_mem[116420] = 16'b0000000000000000;
	sram_mem[116421] = 16'b0000000000000000;
	sram_mem[116422] = 16'b0000000000000000;
	sram_mem[116423] = 16'b0000000000000000;
	sram_mem[116424] = 16'b0000000000000000;
	sram_mem[116425] = 16'b0000000000000000;
	sram_mem[116426] = 16'b0000000000000000;
	sram_mem[116427] = 16'b0000000000000000;
	sram_mem[116428] = 16'b0000000000000000;
	sram_mem[116429] = 16'b0000000000000000;
	sram_mem[116430] = 16'b0000000000000000;
	sram_mem[116431] = 16'b0000000000000000;
	sram_mem[116432] = 16'b0000000000000000;
	sram_mem[116433] = 16'b0000000000000000;
	sram_mem[116434] = 16'b0000000000000000;
	sram_mem[116435] = 16'b0000000000000000;
	sram_mem[116436] = 16'b0000000000000000;
	sram_mem[116437] = 16'b0000000000000000;
	sram_mem[116438] = 16'b0000000000000000;
	sram_mem[116439] = 16'b0000000000000000;
	sram_mem[116440] = 16'b0000000000000000;
	sram_mem[116441] = 16'b0000000000000000;
	sram_mem[116442] = 16'b0000000000000000;
	sram_mem[116443] = 16'b0000000000000000;
	sram_mem[116444] = 16'b0000000000000000;
	sram_mem[116445] = 16'b0000000000000000;
	sram_mem[116446] = 16'b0000000000000000;
	sram_mem[116447] = 16'b0000000000000000;
	sram_mem[116448] = 16'b0000000000000000;
	sram_mem[116449] = 16'b0000000000000000;
	sram_mem[116450] = 16'b0000000000000000;
	sram_mem[116451] = 16'b0000000000000000;
	sram_mem[116452] = 16'b0000000000000000;
	sram_mem[116453] = 16'b0000000000000000;
	sram_mem[116454] = 16'b0000000000000000;
	sram_mem[116455] = 16'b0000000000000000;
	sram_mem[116456] = 16'b0000000000000000;
	sram_mem[116457] = 16'b0000000000000000;
	sram_mem[116458] = 16'b0000000000000000;
	sram_mem[116459] = 16'b0000000000000000;
	sram_mem[116460] = 16'b0000000000000000;
	sram_mem[116461] = 16'b0000000000000000;
	sram_mem[116462] = 16'b0000000000000000;
	sram_mem[116463] = 16'b0000000000000000;
	sram_mem[116464] = 16'b0000000000000000;
	sram_mem[116465] = 16'b0000000000000000;
	sram_mem[116466] = 16'b0000000000000000;
	sram_mem[116467] = 16'b0000000000000000;
	sram_mem[116468] = 16'b0000000000000000;
	sram_mem[116469] = 16'b0000000000000000;
	sram_mem[116470] = 16'b0000000000000000;
	sram_mem[116471] = 16'b0000000000000000;
	sram_mem[116472] = 16'b0000000000000000;
	sram_mem[116473] = 16'b0000000000000000;
	sram_mem[116474] = 16'b0000000000000000;
	sram_mem[116475] = 16'b0000000000000000;
	sram_mem[116476] = 16'b0000000000000000;
	sram_mem[116477] = 16'b0000000000000000;
	sram_mem[116478] = 16'b0000000000000000;
	sram_mem[116479] = 16'b0000000000000000;
	sram_mem[116480] = 16'b0000000000000000;
	sram_mem[116481] = 16'b0000000000000000;
	sram_mem[116482] = 16'b0000000000000000;
	sram_mem[116483] = 16'b0000000000000000;
	sram_mem[116484] = 16'b0000000000000000;
	sram_mem[116485] = 16'b0000000000000000;
	sram_mem[116486] = 16'b0000000000000000;
	sram_mem[116487] = 16'b0000000000000000;
	sram_mem[116488] = 16'b0000000000000000;
	sram_mem[116489] = 16'b0000000000000000;
	sram_mem[116490] = 16'b0000000000000000;
	sram_mem[116491] = 16'b0000000000000000;
	sram_mem[116492] = 16'b0000000000000000;
	sram_mem[116493] = 16'b0000000000000000;
	sram_mem[116494] = 16'b0000000000000000;
	sram_mem[116495] = 16'b0000000000000000;
	sram_mem[116496] = 16'b0000000000000000;
	sram_mem[116497] = 16'b0000000000000000;
	sram_mem[116498] = 16'b0000000000000000;
	sram_mem[116499] = 16'b0000000000000000;
	sram_mem[116500] = 16'b0000000000000000;
	sram_mem[116501] = 16'b0000000000000000;
	sram_mem[116502] = 16'b0000000000000000;
	sram_mem[116503] = 16'b0000000000000000;
	sram_mem[116504] = 16'b0000000000000000;
	sram_mem[116505] = 16'b0000000000000000;
	sram_mem[116506] = 16'b0000000000000000;
	sram_mem[116507] = 16'b0000000000000000;
	sram_mem[116508] = 16'b0000000000000000;
	sram_mem[116509] = 16'b0000000000000000;
	sram_mem[116510] = 16'b0000000000000000;
	sram_mem[116511] = 16'b0000000000000000;
	sram_mem[116512] = 16'b0000000000000000;
	sram_mem[116513] = 16'b0000000000000000;
	sram_mem[116514] = 16'b0000000000000000;
	sram_mem[116515] = 16'b0000000000000000;
	sram_mem[116516] = 16'b0000000000000000;
	sram_mem[116517] = 16'b0000000000000000;
	sram_mem[116518] = 16'b0000000000000000;
	sram_mem[116519] = 16'b0000000000000000;
	sram_mem[116520] = 16'b0000000000000000;
	sram_mem[116521] = 16'b0000000000000000;
	sram_mem[116522] = 16'b0000000000000000;
	sram_mem[116523] = 16'b0000000000000000;
	sram_mem[116524] = 16'b0000000000000000;
	sram_mem[116525] = 16'b0000000000000000;
	sram_mem[116526] = 16'b0000000000000000;
	sram_mem[116527] = 16'b0000000000000000;
	sram_mem[116528] = 16'b0000000000000000;
	sram_mem[116529] = 16'b0000000000000000;
	sram_mem[116530] = 16'b0000000000000000;
	sram_mem[116531] = 16'b0000000000000000;
	sram_mem[116532] = 16'b0000000000000000;
	sram_mem[116533] = 16'b0000000000000000;
	sram_mem[116534] = 16'b0000000000000000;
	sram_mem[116535] = 16'b0000000000000000;
	sram_mem[116536] = 16'b0000000000000000;
	sram_mem[116537] = 16'b0000000000000000;
	sram_mem[116538] = 16'b0000000000000000;
	sram_mem[116539] = 16'b0000000000000000;
	sram_mem[116540] = 16'b0000000000000000;
	sram_mem[116541] = 16'b0000000000000000;
	sram_mem[116542] = 16'b0000000000000000;
	sram_mem[116543] = 16'b0000000000000000;
	sram_mem[116544] = 16'b0000000000000000;
	sram_mem[116545] = 16'b0000000000000000;
	sram_mem[116546] = 16'b0000000000000000;
	sram_mem[116547] = 16'b0000000000000000;
	sram_mem[116548] = 16'b0000000000000000;
	sram_mem[116549] = 16'b0000000000000000;
	sram_mem[116550] = 16'b0000000000000000;
	sram_mem[116551] = 16'b0000000000000000;
	sram_mem[116552] = 16'b0000000000000000;
	sram_mem[116553] = 16'b0000000000000000;
	sram_mem[116554] = 16'b0000000000000000;
	sram_mem[116555] = 16'b0000000000000000;
	sram_mem[116556] = 16'b0000000000000000;
	sram_mem[116557] = 16'b0000000000000000;
	sram_mem[116558] = 16'b0000000000000000;
	sram_mem[116559] = 16'b0000000000000000;
	sram_mem[116560] = 16'b0000000000000000;
	sram_mem[116561] = 16'b0000000000000000;
	sram_mem[116562] = 16'b0000000000000000;
	sram_mem[116563] = 16'b0000000000000000;
	sram_mem[116564] = 16'b0000000000000000;
	sram_mem[116565] = 16'b0000000000000000;
	sram_mem[116566] = 16'b0000000000000000;
	sram_mem[116567] = 16'b0000000000000000;
	sram_mem[116568] = 16'b0000000000000000;
	sram_mem[116569] = 16'b0000000000000000;
	sram_mem[116570] = 16'b0000000000000000;
	sram_mem[116571] = 16'b0000000000000000;
	sram_mem[116572] = 16'b0000000000000000;
	sram_mem[116573] = 16'b0000000000000000;
	sram_mem[116574] = 16'b0000000000000000;
	sram_mem[116575] = 16'b0000000000000000;
	sram_mem[116576] = 16'b0000000000000000;
	sram_mem[116577] = 16'b0000000000000000;
	sram_mem[116578] = 16'b0000000000000000;
	sram_mem[116579] = 16'b0000000000000000;
	sram_mem[116580] = 16'b0000000000000000;
	sram_mem[116581] = 16'b0000000000000000;
	sram_mem[116582] = 16'b0000000000000000;
	sram_mem[116583] = 16'b0000000000000000;
	sram_mem[116584] = 16'b0000000000000000;
	sram_mem[116585] = 16'b0000000000000000;
	sram_mem[116586] = 16'b0000000000000000;
	sram_mem[116587] = 16'b0000000000000000;
	sram_mem[116588] = 16'b0000000000000000;
	sram_mem[116589] = 16'b0000000000000000;
	sram_mem[116590] = 16'b0000000000000000;
	sram_mem[116591] = 16'b0000000000000000;
	sram_mem[116592] = 16'b0000000000000000;
	sram_mem[116593] = 16'b0000000000000000;
	sram_mem[116594] = 16'b0000000000000000;
	sram_mem[116595] = 16'b0000000000000000;
	sram_mem[116596] = 16'b0000000000000000;
	sram_mem[116597] = 16'b0000000000000000;
	sram_mem[116598] = 16'b0000000000000000;
	sram_mem[116599] = 16'b0000000000000000;
	sram_mem[116600] = 16'b0000000000000000;
	sram_mem[116601] = 16'b0000000000000000;
	sram_mem[116602] = 16'b0000000000000000;
	sram_mem[116603] = 16'b0000000000000000;
	sram_mem[116604] = 16'b0000000000000000;
	sram_mem[116605] = 16'b0000000000000000;
	sram_mem[116606] = 16'b0000000000000000;
	sram_mem[116607] = 16'b0000000000000000;
	sram_mem[116608] = 16'b0000000000000000;
	sram_mem[116609] = 16'b0000000000000000;
	sram_mem[116610] = 16'b0000000000000000;
	sram_mem[116611] = 16'b0000000000000000;
	sram_mem[116612] = 16'b0000000000000000;
	sram_mem[116613] = 16'b0000000000000000;
	sram_mem[116614] = 16'b0000000000000000;
	sram_mem[116615] = 16'b0000000000000000;
	sram_mem[116616] = 16'b0000000000000000;
	sram_mem[116617] = 16'b0000000000000000;
	sram_mem[116618] = 16'b0000000000000000;
	sram_mem[116619] = 16'b0000000000000000;
	sram_mem[116620] = 16'b0000000000000000;
	sram_mem[116621] = 16'b0000000000000000;
	sram_mem[116622] = 16'b0000000000000000;
	sram_mem[116623] = 16'b0000000000000000;
	sram_mem[116624] = 16'b0000000000000000;
	sram_mem[116625] = 16'b0000000000000000;
	sram_mem[116626] = 16'b0000000000000000;
	sram_mem[116627] = 16'b0000000000000000;
	sram_mem[116628] = 16'b0000000000000000;
	sram_mem[116629] = 16'b0000000000000000;
	sram_mem[116630] = 16'b0000000000000000;
	sram_mem[116631] = 16'b0000000000000000;
	sram_mem[116632] = 16'b0000000000000000;
	sram_mem[116633] = 16'b0000000000000000;
	sram_mem[116634] = 16'b0000000000000000;
	sram_mem[116635] = 16'b0000000000000000;
	sram_mem[116636] = 16'b0000000000000000;
	sram_mem[116637] = 16'b0000000000000000;
	sram_mem[116638] = 16'b0000000000000000;
	sram_mem[116639] = 16'b0000000000000000;
	sram_mem[116640] = 16'b0000000000000000;
	sram_mem[116641] = 16'b0000000000000000;
	sram_mem[116642] = 16'b0000000000000000;
	sram_mem[116643] = 16'b0000000000000000;
	sram_mem[116644] = 16'b0000000000000000;
	sram_mem[116645] = 16'b0000000000000000;
	sram_mem[116646] = 16'b0000000000000000;
	sram_mem[116647] = 16'b0000000000000000;
	sram_mem[116648] = 16'b0000000000000000;
	sram_mem[116649] = 16'b0000000000000000;
	sram_mem[116650] = 16'b0000000000000000;
	sram_mem[116651] = 16'b0000000000000000;
	sram_mem[116652] = 16'b0000000000000000;
	sram_mem[116653] = 16'b0000000000000000;
	sram_mem[116654] = 16'b0000000000000000;
	sram_mem[116655] = 16'b0000000000000000;
	sram_mem[116656] = 16'b0000000000000000;
	sram_mem[116657] = 16'b0000000000000000;
	sram_mem[116658] = 16'b0000000000000000;
	sram_mem[116659] = 16'b0000000000000000;
	sram_mem[116660] = 16'b0000000000000000;
	sram_mem[116661] = 16'b0000000000000000;
	sram_mem[116662] = 16'b0000000000000000;
	sram_mem[116663] = 16'b0000000000000000;
	sram_mem[116664] = 16'b0000000000000000;
	sram_mem[116665] = 16'b0000000000000000;
	sram_mem[116666] = 16'b0000000000000000;
	sram_mem[116667] = 16'b0000000000000000;
	sram_mem[116668] = 16'b0000000000000000;
	sram_mem[116669] = 16'b0000000000000000;
	sram_mem[116670] = 16'b0000000000000000;
	sram_mem[116671] = 16'b0000000000000000;
	sram_mem[116672] = 16'b0000000000000000;
	sram_mem[116673] = 16'b0000000000000000;
	sram_mem[116674] = 16'b0000000000000000;
	sram_mem[116675] = 16'b0000000000000000;
	sram_mem[116676] = 16'b0000000000000000;
	sram_mem[116677] = 16'b0000000000000000;
	sram_mem[116678] = 16'b0000000000000000;
	sram_mem[116679] = 16'b0000000000000000;
	sram_mem[116680] = 16'b0000000000000000;
	sram_mem[116681] = 16'b0000000000000000;
	sram_mem[116682] = 16'b0000000000000000;
	sram_mem[116683] = 16'b0000000000000000;
	sram_mem[116684] = 16'b0000000000000000;
	sram_mem[116685] = 16'b0000000000000000;
	sram_mem[116686] = 16'b0000000000000000;
	sram_mem[116687] = 16'b0000000000000000;
	sram_mem[116688] = 16'b0000000000000000;
	sram_mem[116689] = 16'b0000000000000000;
	sram_mem[116690] = 16'b0000000000000000;
	sram_mem[116691] = 16'b0000000000000000;
	sram_mem[116692] = 16'b0000000000000000;
	sram_mem[116693] = 16'b0000000000000000;
	sram_mem[116694] = 16'b0000000000000000;
	sram_mem[116695] = 16'b0000000000000000;
	sram_mem[116696] = 16'b0000000000000000;
	sram_mem[116697] = 16'b0000000000000000;
	sram_mem[116698] = 16'b0000000000000000;
	sram_mem[116699] = 16'b0000000000000000;
	sram_mem[116700] = 16'b0000000000000000;
	sram_mem[116701] = 16'b0000000000000000;
	sram_mem[116702] = 16'b0000000000000000;
	sram_mem[116703] = 16'b0000000000000000;
	sram_mem[116704] = 16'b0000000000000000;
	sram_mem[116705] = 16'b0000000000000000;
	sram_mem[116706] = 16'b0000000000000000;
	sram_mem[116707] = 16'b0000000000000000;
	sram_mem[116708] = 16'b0000000000000000;
	sram_mem[116709] = 16'b0000000000000000;
	sram_mem[116710] = 16'b0000000000000000;
	sram_mem[116711] = 16'b0000000000000000;
	sram_mem[116712] = 16'b0000000000000000;
	sram_mem[116713] = 16'b0000000000000000;
	sram_mem[116714] = 16'b0000000000000000;
	sram_mem[116715] = 16'b0000000000000000;
	sram_mem[116716] = 16'b0000000000000000;
	sram_mem[116717] = 16'b0000000000000000;
	sram_mem[116718] = 16'b0000000000000000;
	sram_mem[116719] = 16'b0000000000000000;
	sram_mem[116720] = 16'b0000000000000000;
	sram_mem[116721] = 16'b0000000000000000;
	sram_mem[116722] = 16'b0000000000000000;
	sram_mem[116723] = 16'b0000000000000000;
	sram_mem[116724] = 16'b0000000000000000;
	sram_mem[116725] = 16'b0000000000000000;
	sram_mem[116726] = 16'b0000000000000000;
	sram_mem[116727] = 16'b0000000000000000;
	sram_mem[116728] = 16'b0000000000000000;
	sram_mem[116729] = 16'b0000000000000000;
	sram_mem[116730] = 16'b0000000000000000;
	sram_mem[116731] = 16'b0000000000000000;
	sram_mem[116732] = 16'b0000000000000000;
	sram_mem[116733] = 16'b0000000000000000;
	sram_mem[116734] = 16'b0000000000000000;
	sram_mem[116735] = 16'b0000000000000000;
	sram_mem[116736] = 16'b0000000000000000;
	sram_mem[116737] = 16'b0000000000000000;
	sram_mem[116738] = 16'b0000000000000000;
	sram_mem[116739] = 16'b0000000000000000;
	sram_mem[116740] = 16'b0000000000000000;
	sram_mem[116741] = 16'b0000000000000000;
	sram_mem[116742] = 16'b0000000000000000;
	sram_mem[116743] = 16'b0000000000000000;
	sram_mem[116744] = 16'b0000000000000000;
	sram_mem[116745] = 16'b0000000000000000;
	sram_mem[116746] = 16'b0000000000000000;
	sram_mem[116747] = 16'b0000000000000000;
	sram_mem[116748] = 16'b0000000000000000;
	sram_mem[116749] = 16'b0000000000000000;
	sram_mem[116750] = 16'b0000000000000000;
	sram_mem[116751] = 16'b0000000000000000;
	sram_mem[116752] = 16'b0000000000000000;
	sram_mem[116753] = 16'b0000000000000000;
	sram_mem[116754] = 16'b0000000000000000;
	sram_mem[116755] = 16'b0000000000000000;
	sram_mem[116756] = 16'b0000000000000000;
	sram_mem[116757] = 16'b0000000000000000;
	sram_mem[116758] = 16'b0000000000000000;
	sram_mem[116759] = 16'b0000000000000000;
	sram_mem[116760] = 16'b0000000000000000;
	sram_mem[116761] = 16'b0000000000000000;
	sram_mem[116762] = 16'b0000000000000000;
	sram_mem[116763] = 16'b0000000000000000;
	sram_mem[116764] = 16'b0000000000000000;
	sram_mem[116765] = 16'b0000000000000000;
	sram_mem[116766] = 16'b0000000000000000;
	sram_mem[116767] = 16'b0000000000000000;
	sram_mem[116768] = 16'b0000000000000000;
	sram_mem[116769] = 16'b0000000000000000;
	sram_mem[116770] = 16'b0000000000000000;
	sram_mem[116771] = 16'b0000000000000000;
	sram_mem[116772] = 16'b0000000000000000;
	sram_mem[116773] = 16'b0000000000000000;
	sram_mem[116774] = 16'b0000000000000000;
	sram_mem[116775] = 16'b0000000000000000;
	sram_mem[116776] = 16'b0000000000000000;
	sram_mem[116777] = 16'b0000000000000000;
	sram_mem[116778] = 16'b0000000000000000;
	sram_mem[116779] = 16'b0000000000000000;
	sram_mem[116780] = 16'b0000000000000000;
	sram_mem[116781] = 16'b0000000000000000;
	sram_mem[116782] = 16'b0000000000000000;
	sram_mem[116783] = 16'b0000000000000000;
	sram_mem[116784] = 16'b0000000000000000;
	sram_mem[116785] = 16'b0000000000000000;
	sram_mem[116786] = 16'b0000000000000000;
	sram_mem[116787] = 16'b0000000000000000;
	sram_mem[116788] = 16'b0000000000000000;
	sram_mem[116789] = 16'b0000000000000000;
	sram_mem[116790] = 16'b0000000000000000;
	sram_mem[116791] = 16'b0000000000000000;
	sram_mem[116792] = 16'b0000000000000000;
	sram_mem[116793] = 16'b0000000000000000;
	sram_mem[116794] = 16'b0000000000000000;
	sram_mem[116795] = 16'b0000000000000000;
	sram_mem[116796] = 16'b0000000000000000;
	sram_mem[116797] = 16'b0000000000000000;
	sram_mem[116798] = 16'b0000000000000000;
	sram_mem[116799] = 16'b0000000000000000;
	sram_mem[116800] = 16'b0000000000000000;
	sram_mem[116801] = 16'b0000000000000000;
	sram_mem[116802] = 16'b0000000000000000;
	sram_mem[116803] = 16'b0000000000000000;
	sram_mem[116804] = 16'b0000000000000000;
	sram_mem[116805] = 16'b0000000000000000;
	sram_mem[116806] = 16'b0000000000000000;
	sram_mem[116807] = 16'b0000000000000000;
	sram_mem[116808] = 16'b0000000000000000;
	sram_mem[116809] = 16'b0000000000000000;
	sram_mem[116810] = 16'b0000000000000000;
	sram_mem[116811] = 16'b0000000000000000;
	sram_mem[116812] = 16'b0000000000000000;
	sram_mem[116813] = 16'b0000000000000000;
	sram_mem[116814] = 16'b0000000000000000;
	sram_mem[116815] = 16'b0000000000000000;
	sram_mem[116816] = 16'b0000000000000000;
	sram_mem[116817] = 16'b0000000000000000;
	sram_mem[116818] = 16'b0000000000000000;
	sram_mem[116819] = 16'b0000000000000000;
	sram_mem[116820] = 16'b0000000000000000;
	sram_mem[116821] = 16'b0000000000000000;
	sram_mem[116822] = 16'b0000000000000000;
	sram_mem[116823] = 16'b0000000000000000;
	sram_mem[116824] = 16'b0000000000000000;
	sram_mem[116825] = 16'b0000000000000000;
	sram_mem[116826] = 16'b0000000000000000;
	sram_mem[116827] = 16'b0000000000000000;
	sram_mem[116828] = 16'b0000000000000000;
	sram_mem[116829] = 16'b0000000000000000;
	sram_mem[116830] = 16'b0000000000000000;
	sram_mem[116831] = 16'b0000000000000000;
	sram_mem[116832] = 16'b0000000000000000;
	sram_mem[116833] = 16'b0000000000000000;
	sram_mem[116834] = 16'b0000000000000000;
	sram_mem[116835] = 16'b0000000000000000;
	sram_mem[116836] = 16'b0000000000000000;
	sram_mem[116837] = 16'b0000000000000000;
	sram_mem[116838] = 16'b0000000000000000;
	sram_mem[116839] = 16'b0000000000000000;
	sram_mem[116840] = 16'b0000000000000000;
	sram_mem[116841] = 16'b0000000000000000;
	sram_mem[116842] = 16'b0000000000000000;
	sram_mem[116843] = 16'b0000000000000000;
	sram_mem[116844] = 16'b0000000000000000;
	sram_mem[116845] = 16'b0000000000000000;
	sram_mem[116846] = 16'b0000000000000000;
	sram_mem[116847] = 16'b0000000000000000;
	sram_mem[116848] = 16'b0000000000000000;
	sram_mem[116849] = 16'b0000000000000000;
	sram_mem[116850] = 16'b0000000000000000;
	sram_mem[116851] = 16'b0000000000000000;
	sram_mem[116852] = 16'b0000000000000000;
	sram_mem[116853] = 16'b0000000000000000;
	sram_mem[116854] = 16'b0000000000000000;
	sram_mem[116855] = 16'b0000000000000000;
	sram_mem[116856] = 16'b0000000000000000;
	sram_mem[116857] = 16'b0000000000000000;
	sram_mem[116858] = 16'b0000000000000000;
	sram_mem[116859] = 16'b0000000000000000;
	sram_mem[116860] = 16'b0000000000000000;
	sram_mem[116861] = 16'b0000000000000000;
	sram_mem[116862] = 16'b0000000000000000;
	sram_mem[116863] = 16'b0000000000000000;
	sram_mem[116864] = 16'b0000000000000000;
	sram_mem[116865] = 16'b0000000000000000;
	sram_mem[116866] = 16'b0000000000000000;
	sram_mem[116867] = 16'b0000000000000000;
	sram_mem[116868] = 16'b0000000000000000;
	sram_mem[116869] = 16'b0000000000000000;
	sram_mem[116870] = 16'b0000000000000000;
	sram_mem[116871] = 16'b0000000000000000;
	sram_mem[116872] = 16'b0000000000000000;
	sram_mem[116873] = 16'b0000000000000000;
	sram_mem[116874] = 16'b0000000000000000;
	sram_mem[116875] = 16'b0000000000000000;
	sram_mem[116876] = 16'b0000000000000000;
	sram_mem[116877] = 16'b0000000000000000;
	sram_mem[116878] = 16'b0000000000000000;
	sram_mem[116879] = 16'b0000000000000000;
	sram_mem[116880] = 16'b0000000000000000;
	sram_mem[116881] = 16'b0000000000000000;
	sram_mem[116882] = 16'b0000000000000000;
	sram_mem[116883] = 16'b0000000000000000;
	sram_mem[116884] = 16'b0000000000000000;
	sram_mem[116885] = 16'b0000000000000000;
	sram_mem[116886] = 16'b0000000000000000;
	sram_mem[116887] = 16'b0000000000000000;
	sram_mem[116888] = 16'b0000000000000000;
	sram_mem[116889] = 16'b0000000000000000;
	sram_mem[116890] = 16'b0000000000000000;
	sram_mem[116891] = 16'b0000000000000000;
	sram_mem[116892] = 16'b0000000000000000;
	sram_mem[116893] = 16'b0000000000000000;
	sram_mem[116894] = 16'b0000000000000000;
	sram_mem[116895] = 16'b0000000000000000;
	sram_mem[116896] = 16'b0000000000000000;
	sram_mem[116897] = 16'b0000000000000000;
	sram_mem[116898] = 16'b0000000000000000;
	sram_mem[116899] = 16'b0000000000000000;
	sram_mem[116900] = 16'b0000000000000000;
	sram_mem[116901] = 16'b0000000000000000;
	sram_mem[116902] = 16'b0000000000000000;
	sram_mem[116903] = 16'b0000000000000000;
	sram_mem[116904] = 16'b0000000000000000;
	sram_mem[116905] = 16'b0000000000000000;
	sram_mem[116906] = 16'b0000000000000000;
	sram_mem[116907] = 16'b0000000000000000;
	sram_mem[116908] = 16'b0000000000000000;
	sram_mem[116909] = 16'b0000000000000000;
	sram_mem[116910] = 16'b0000000000000000;
	sram_mem[116911] = 16'b0000000000000000;
	sram_mem[116912] = 16'b0000000000000000;
	sram_mem[116913] = 16'b0000000000000000;
	sram_mem[116914] = 16'b0000000000000000;
	sram_mem[116915] = 16'b0000000000000000;
	sram_mem[116916] = 16'b0000000000000000;
	sram_mem[116917] = 16'b0000000000000000;
	sram_mem[116918] = 16'b0000000000000000;
	sram_mem[116919] = 16'b0000000000000000;
	sram_mem[116920] = 16'b0000000000000000;
	sram_mem[116921] = 16'b0000000000000000;
	sram_mem[116922] = 16'b0000000000000000;
	sram_mem[116923] = 16'b0000000000000000;
	sram_mem[116924] = 16'b0000000000000000;
	sram_mem[116925] = 16'b0000000000000000;
	sram_mem[116926] = 16'b0000000000000000;
	sram_mem[116927] = 16'b0000000000000000;
	sram_mem[116928] = 16'b0000000000000000;
	sram_mem[116929] = 16'b0000000000000000;
	sram_mem[116930] = 16'b0000000000000000;
	sram_mem[116931] = 16'b0000000000000000;
	sram_mem[116932] = 16'b0000000000000000;
	sram_mem[116933] = 16'b0000000000000000;
	sram_mem[116934] = 16'b0000000000000000;
	sram_mem[116935] = 16'b0000000000000000;
	sram_mem[116936] = 16'b0000000000000000;
	sram_mem[116937] = 16'b0000000000000000;
	sram_mem[116938] = 16'b0000000000000000;
	sram_mem[116939] = 16'b0000000000000000;
	sram_mem[116940] = 16'b0000000000000000;
	sram_mem[116941] = 16'b0000000000000000;
	sram_mem[116942] = 16'b0000000000000000;
	sram_mem[116943] = 16'b0000000000000000;
	sram_mem[116944] = 16'b0000000000000000;
	sram_mem[116945] = 16'b0000000000000000;
	sram_mem[116946] = 16'b0000000000000000;
	sram_mem[116947] = 16'b0000000000000000;
	sram_mem[116948] = 16'b0000000000000000;
	sram_mem[116949] = 16'b0000000000000000;
	sram_mem[116950] = 16'b0000000000000000;
	sram_mem[116951] = 16'b0000000000000000;
	sram_mem[116952] = 16'b0000000000000000;
	sram_mem[116953] = 16'b0000000000000000;
	sram_mem[116954] = 16'b0000000000000000;
	sram_mem[116955] = 16'b0000000000000000;
	sram_mem[116956] = 16'b0000000000000000;
	sram_mem[116957] = 16'b0000000000000000;
	sram_mem[116958] = 16'b0000000000000000;
	sram_mem[116959] = 16'b0000000000000000;
	sram_mem[116960] = 16'b0000000000000000;
	sram_mem[116961] = 16'b0000000000000000;
	sram_mem[116962] = 16'b0000000000000000;
	sram_mem[116963] = 16'b0000000000000000;
	sram_mem[116964] = 16'b0000000000000000;
	sram_mem[116965] = 16'b0000000000000000;
	sram_mem[116966] = 16'b0000000000000000;
	sram_mem[116967] = 16'b0000000000000000;
	sram_mem[116968] = 16'b0000000000000000;
	sram_mem[116969] = 16'b0000000000000000;
	sram_mem[116970] = 16'b0000000000000000;
	sram_mem[116971] = 16'b0000000000000000;
	sram_mem[116972] = 16'b0000000000000000;
	sram_mem[116973] = 16'b0000000000000000;
	sram_mem[116974] = 16'b0000000000000000;
	sram_mem[116975] = 16'b0000000000000000;
	sram_mem[116976] = 16'b0000000000000000;
	sram_mem[116977] = 16'b0000000000000000;
	sram_mem[116978] = 16'b0000000000000000;
	sram_mem[116979] = 16'b0000000000000000;
	sram_mem[116980] = 16'b0000000000000000;
	sram_mem[116981] = 16'b0000000000000000;
	sram_mem[116982] = 16'b0000000000000000;
	sram_mem[116983] = 16'b0000000000000000;
	sram_mem[116984] = 16'b0000000000000000;
	sram_mem[116985] = 16'b0000000000000000;
	sram_mem[116986] = 16'b0000000000000000;
	sram_mem[116987] = 16'b0000000000000000;
	sram_mem[116988] = 16'b0000000000000000;
	sram_mem[116989] = 16'b0000000000000000;
	sram_mem[116990] = 16'b0000000000000000;
	sram_mem[116991] = 16'b0000000000000000;
	sram_mem[116992] = 16'b0000000000000000;
	sram_mem[116993] = 16'b0000000000000000;
	sram_mem[116994] = 16'b0000000000000000;
	sram_mem[116995] = 16'b0000000000000000;
	sram_mem[116996] = 16'b0000000000000000;
	sram_mem[116997] = 16'b0000000000000000;
	sram_mem[116998] = 16'b0000000000000000;
	sram_mem[116999] = 16'b0000000000000000;
	sram_mem[117000] = 16'b0000000000000000;
	sram_mem[117001] = 16'b0000000000000000;
	sram_mem[117002] = 16'b0000000000000000;
	sram_mem[117003] = 16'b0000000000000000;
	sram_mem[117004] = 16'b0000000000000000;
	sram_mem[117005] = 16'b0000000000000000;
	sram_mem[117006] = 16'b0000000000000000;
	sram_mem[117007] = 16'b0000000000000000;
	sram_mem[117008] = 16'b0000000000000000;
	sram_mem[117009] = 16'b0000000000000000;
	sram_mem[117010] = 16'b0000000000000000;
	sram_mem[117011] = 16'b0000000000000000;
	sram_mem[117012] = 16'b0000000000000000;
	sram_mem[117013] = 16'b0000000000000000;
	sram_mem[117014] = 16'b0000000000000000;
	sram_mem[117015] = 16'b0000000000000000;
	sram_mem[117016] = 16'b0000000000000000;
	sram_mem[117017] = 16'b0000000000000000;
	sram_mem[117018] = 16'b0000000000000000;
	sram_mem[117019] = 16'b0000000000000000;
	sram_mem[117020] = 16'b0000000000000000;
	sram_mem[117021] = 16'b0000000000000000;
	sram_mem[117022] = 16'b0000000000000000;
	sram_mem[117023] = 16'b0000000000000000;
	sram_mem[117024] = 16'b0000000000000000;
	sram_mem[117025] = 16'b0000000000000000;
	sram_mem[117026] = 16'b0000000000000000;
	sram_mem[117027] = 16'b0000000000000000;
	sram_mem[117028] = 16'b0000000000000000;
	sram_mem[117029] = 16'b0000000000000000;
	sram_mem[117030] = 16'b0000000000000000;
	sram_mem[117031] = 16'b0000000000000000;
	sram_mem[117032] = 16'b0000000000000000;
	sram_mem[117033] = 16'b0000000000000000;
	sram_mem[117034] = 16'b0000000000000000;
	sram_mem[117035] = 16'b0000000000000000;
	sram_mem[117036] = 16'b0000000000000000;
	sram_mem[117037] = 16'b0000000000000000;
	sram_mem[117038] = 16'b0000000000000000;
	sram_mem[117039] = 16'b0000000000000000;
	sram_mem[117040] = 16'b0000000000000000;
	sram_mem[117041] = 16'b0000000000000000;
	sram_mem[117042] = 16'b0000000000000000;
	sram_mem[117043] = 16'b0000000000000000;
	sram_mem[117044] = 16'b0000000000000000;
	sram_mem[117045] = 16'b0000000000000000;
	sram_mem[117046] = 16'b0000000000000000;
	sram_mem[117047] = 16'b0000000000000000;
	sram_mem[117048] = 16'b0000000000000000;
	sram_mem[117049] = 16'b0000000000000000;
	sram_mem[117050] = 16'b0000000000000000;
	sram_mem[117051] = 16'b0000000000000000;
	sram_mem[117052] = 16'b0000000000000000;
	sram_mem[117053] = 16'b0000000000000000;
	sram_mem[117054] = 16'b0000000000000000;
	sram_mem[117055] = 16'b0000000000000000;
	sram_mem[117056] = 16'b0000000000000000;
	sram_mem[117057] = 16'b0000000000000000;
	sram_mem[117058] = 16'b0000000000000000;
	sram_mem[117059] = 16'b0000000000000000;
	sram_mem[117060] = 16'b0000000000000000;
	sram_mem[117061] = 16'b0000000000000000;
	sram_mem[117062] = 16'b0000000000000000;
	sram_mem[117063] = 16'b0000000000000000;
	sram_mem[117064] = 16'b0000000000000000;
	sram_mem[117065] = 16'b0000000000000000;
	sram_mem[117066] = 16'b0000000000000000;
	sram_mem[117067] = 16'b0000000000000000;
	sram_mem[117068] = 16'b0000000000000000;
	sram_mem[117069] = 16'b0000000000000000;
	sram_mem[117070] = 16'b0000000000000000;
	sram_mem[117071] = 16'b0000000000000000;
	sram_mem[117072] = 16'b0000000000000000;
	sram_mem[117073] = 16'b0000000000000000;
	sram_mem[117074] = 16'b0000000000000000;
	sram_mem[117075] = 16'b0000000000000000;
	sram_mem[117076] = 16'b0000000000000000;
	sram_mem[117077] = 16'b0000000000000000;
	sram_mem[117078] = 16'b0000000000000000;
	sram_mem[117079] = 16'b0000000000000000;
	sram_mem[117080] = 16'b0000000000000000;
	sram_mem[117081] = 16'b0000000000000000;
	sram_mem[117082] = 16'b0000000000000000;
	sram_mem[117083] = 16'b0000000000000000;
	sram_mem[117084] = 16'b0000000000000000;
	sram_mem[117085] = 16'b0000000000000000;
	sram_mem[117086] = 16'b0000000000000000;
	sram_mem[117087] = 16'b0000000000000000;
	sram_mem[117088] = 16'b0000000000000000;
	sram_mem[117089] = 16'b0000000000000000;
	sram_mem[117090] = 16'b0000000000000000;
	sram_mem[117091] = 16'b0000000000000000;
	sram_mem[117092] = 16'b0000000000000000;
	sram_mem[117093] = 16'b0000000000000000;
	sram_mem[117094] = 16'b0000000000000000;
	sram_mem[117095] = 16'b0000000000000000;
	sram_mem[117096] = 16'b0000000000000000;
	sram_mem[117097] = 16'b0000000000000000;
	sram_mem[117098] = 16'b0000000000000000;
	sram_mem[117099] = 16'b0000000000000000;
	sram_mem[117100] = 16'b0000000000000000;
	sram_mem[117101] = 16'b0000000000000000;
	sram_mem[117102] = 16'b0000000000000000;
	sram_mem[117103] = 16'b0000000000000000;
	sram_mem[117104] = 16'b0000000000000000;
	sram_mem[117105] = 16'b0000000000000000;
	sram_mem[117106] = 16'b0000000000000000;
	sram_mem[117107] = 16'b0000000000000000;
	sram_mem[117108] = 16'b0000000000000000;
	sram_mem[117109] = 16'b0000000000000000;
	sram_mem[117110] = 16'b0000000000000000;
	sram_mem[117111] = 16'b0000000000000000;
	sram_mem[117112] = 16'b0000000000000000;
	sram_mem[117113] = 16'b0000000000000000;
	sram_mem[117114] = 16'b0000000000000000;
	sram_mem[117115] = 16'b0000000000000000;
	sram_mem[117116] = 16'b0000000000000000;
	sram_mem[117117] = 16'b0000000000000000;
	sram_mem[117118] = 16'b0000000000000000;
	sram_mem[117119] = 16'b0000000000000000;
	sram_mem[117120] = 16'b0000000000000000;
	sram_mem[117121] = 16'b0000000000000000;
	sram_mem[117122] = 16'b0000000000000000;
	sram_mem[117123] = 16'b0000000000000000;
	sram_mem[117124] = 16'b0000000000000000;
	sram_mem[117125] = 16'b0000000000000000;
	sram_mem[117126] = 16'b0000000000000000;
	sram_mem[117127] = 16'b0000000000000000;
	sram_mem[117128] = 16'b0000000000000000;
	sram_mem[117129] = 16'b0000000000000000;
	sram_mem[117130] = 16'b0000000000000000;
	sram_mem[117131] = 16'b0000000000000000;
	sram_mem[117132] = 16'b0000000000000000;
	sram_mem[117133] = 16'b0000000000000000;
	sram_mem[117134] = 16'b0000000000000000;
	sram_mem[117135] = 16'b0000000000000000;
	sram_mem[117136] = 16'b0000000000000000;
	sram_mem[117137] = 16'b0000000000000000;
	sram_mem[117138] = 16'b0000000000000000;
	sram_mem[117139] = 16'b0000000000000000;
	sram_mem[117140] = 16'b0000000000000000;
	sram_mem[117141] = 16'b0000000000000000;
	sram_mem[117142] = 16'b0000000000000000;
	sram_mem[117143] = 16'b0000000000000000;
	sram_mem[117144] = 16'b0000000000000000;
	sram_mem[117145] = 16'b0000000000000000;
	sram_mem[117146] = 16'b0000000000000000;
	sram_mem[117147] = 16'b0000000000000000;
	sram_mem[117148] = 16'b0000000000000000;
	sram_mem[117149] = 16'b0000000000000000;
	sram_mem[117150] = 16'b0000000000000000;
	sram_mem[117151] = 16'b0000000000000000;
	sram_mem[117152] = 16'b0000000000000000;
	sram_mem[117153] = 16'b0000000000000000;
	sram_mem[117154] = 16'b0000000000000000;
	sram_mem[117155] = 16'b0000000000000000;
	sram_mem[117156] = 16'b0000000000000000;
	sram_mem[117157] = 16'b0000000000000000;
	sram_mem[117158] = 16'b0000000000000000;
	sram_mem[117159] = 16'b0000000000000000;
	sram_mem[117160] = 16'b0000000000000000;
	sram_mem[117161] = 16'b0000000000000000;
	sram_mem[117162] = 16'b0000000000000000;
	sram_mem[117163] = 16'b0000000000000000;
	sram_mem[117164] = 16'b0000000000000000;
	sram_mem[117165] = 16'b0000000000000000;
	sram_mem[117166] = 16'b0000000000000000;
	sram_mem[117167] = 16'b0000000000000000;
	sram_mem[117168] = 16'b0000000000000000;
	sram_mem[117169] = 16'b0000000000000000;
	sram_mem[117170] = 16'b0000000000000000;
	sram_mem[117171] = 16'b0000000000000000;
	sram_mem[117172] = 16'b0000000000000000;
	sram_mem[117173] = 16'b0000000000000000;
	sram_mem[117174] = 16'b0000000000000000;
	sram_mem[117175] = 16'b0000000000000000;
	sram_mem[117176] = 16'b0000000000000000;
	sram_mem[117177] = 16'b0000000000000000;
	sram_mem[117178] = 16'b0000000000000000;
	sram_mem[117179] = 16'b0000000000000000;
	sram_mem[117180] = 16'b0000000000000000;
	sram_mem[117181] = 16'b0000000000000000;
	sram_mem[117182] = 16'b0000000000000000;
	sram_mem[117183] = 16'b0000000000000000;
	sram_mem[117184] = 16'b0000000000000000;
	sram_mem[117185] = 16'b0000000000000000;
	sram_mem[117186] = 16'b0000000000000000;
	sram_mem[117187] = 16'b0000000000000000;
	sram_mem[117188] = 16'b0000000000000000;
	sram_mem[117189] = 16'b0000000000000000;
	sram_mem[117190] = 16'b0000000000000000;
	sram_mem[117191] = 16'b0000000000000000;
	sram_mem[117192] = 16'b0000000000000000;
	sram_mem[117193] = 16'b0000000000000000;
	sram_mem[117194] = 16'b0000000000000000;
	sram_mem[117195] = 16'b0000000000000000;
	sram_mem[117196] = 16'b0000000000000000;
	sram_mem[117197] = 16'b0000000000000000;
	sram_mem[117198] = 16'b0000000000000000;
	sram_mem[117199] = 16'b0000000000000000;
	sram_mem[117200] = 16'b0000000000000000;
	sram_mem[117201] = 16'b0000000000000000;
	sram_mem[117202] = 16'b0000000000000000;
	sram_mem[117203] = 16'b0000000000000000;
	sram_mem[117204] = 16'b0000000000000000;
	sram_mem[117205] = 16'b0000000000000000;
	sram_mem[117206] = 16'b0000000000000000;
	sram_mem[117207] = 16'b0000000000000000;
	sram_mem[117208] = 16'b0000000000000000;
	sram_mem[117209] = 16'b0000000000000000;
	sram_mem[117210] = 16'b0000000000000000;
	sram_mem[117211] = 16'b0000000000000000;
	sram_mem[117212] = 16'b0000000000000000;
	sram_mem[117213] = 16'b0000000000000000;
	sram_mem[117214] = 16'b0000000000000000;
	sram_mem[117215] = 16'b0000000000000000;
	sram_mem[117216] = 16'b0000000000000000;
	sram_mem[117217] = 16'b0000000000000000;
	sram_mem[117218] = 16'b0000000000000000;
	sram_mem[117219] = 16'b0000000000000000;
	sram_mem[117220] = 16'b0000000000000000;
	sram_mem[117221] = 16'b0000000000000000;
	sram_mem[117222] = 16'b0000000000000000;
	sram_mem[117223] = 16'b0000000000000000;
	sram_mem[117224] = 16'b0000000000000000;
	sram_mem[117225] = 16'b0000000000000000;
	sram_mem[117226] = 16'b0000000000000000;
	sram_mem[117227] = 16'b0000000000000000;
	sram_mem[117228] = 16'b0000000000000000;
	sram_mem[117229] = 16'b0000000000000000;
	sram_mem[117230] = 16'b0000000000000000;
	sram_mem[117231] = 16'b0000000000000000;
	sram_mem[117232] = 16'b0000000000000000;
	sram_mem[117233] = 16'b0000000000000000;
	sram_mem[117234] = 16'b0000000000000000;
	sram_mem[117235] = 16'b0000000000000000;
	sram_mem[117236] = 16'b0000000000000000;
	sram_mem[117237] = 16'b0000000000000000;
	sram_mem[117238] = 16'b0000000000000000;
	sram_mem[117239] = 16'b0000000000000000;
	sram_mem[117240] = 16'b0000000000000000;
	sram_mem[117241] = 16'b0000000000000000;
	sram_mem[117242] = 16'b0000000000000000;
	sram_mem[117243] = 16'b0000000000000000;
	sram_mem[117244] = 16'b0000000000000000;
	sram_mem[117245] = 16'b0000000000000000;
	sram_mem[117246] = 16'b0000000000000000;
	sram_mem[117247] = 16'b0000000000000000;
	sram_mem[117248] = 16'b0000000000000000;
	sram_mem[117249] = 16'b0000000000000000;
	sram_mem[117250] = 16'b0000000000000000;
	sram_mem[117251] = 16'b0000000000000000;
	sram_mem[117252] = 16'b0000000000000000;
	sram_mem[117253] = 16'b0000000000000000;
	sram_mem[117254] = 16'b0000000000000000;
	sram_mem[117255] = 16'b0000000000000000;
	sram_mem[117256] = 16'b0000000000000000;
	sram_mem[117257] = 16'b0000000000000000;
	sram_mem[117258] = 16'b0000000000000000;
	sram_mem[117259] = 16'b0000000000000000;
	sram_mem[117260] = 16'b0000000000000000;
	sram_mem[117261] = 16'b0000000000000000;
	sram_mem[117262] = 16'b0000000000000000;
	sram_mem[117263] = 16'b0000000000000000;
	sram_mem[117264] = 16'b0000000000000000;
	sram_mem[117265] = 16'b0000000000000000;
	sram_mem[117266] = 16'b0000000000000000;
	sram_mem[117267] = 16'b0000000000000000;
	sram_mem[117268] = 16'b0000000000000000;
	sram_mem[117269] = 16'b0000000000000000;
	sram_mem[117270] = 16'b0000000000000000;
	sram_mem[117271] = 16'b0000000000000000;
	sram_mem[117272] = 16'b0000000000000000;
	sram_mem[117273] = 16'b0000000000000000;
	sram_mem[117274] = 16'b0000000000000000;
	sram_mem[117275] = 16'b0000000000000000;
	sram_mem[117276] = 16'b0000000000000000;
	sram_mem[117277] = 16'b0000000000000000;
	sram_mem[117278] = 16'b0000000000000000;
	sram_mem[117279] = 16'b0000000000000000;
	sram_mem[117280] = 16'b0000000000000000;
	sram_mem[117281] = 16'b0000000000000000;
	sram_mem[117282] = 16'b0000000000000000;
	sram_mem[117283] = 16'b0000000000000000;
	sram_mem[117284] = 16'b0000000000000000;
	sram_mem[117285] = 16'b0000000000000000;
	sram_mem[117286] = 16'b0000000000000000;
	sram_mem[117287] = 16'b0000000000000000;
	sram_mem[117288] = 16'b0000000000000000;
	sram_mem[117289] = 16'b0000000000000000;
	sram_mem[117290] = 16'b0000000000000000;
	sram_mem[117291] = 16'b0000000000000000;
	sram_mem[117292] = 16'b0000000000000000;
	sram_mem[117293] = 16'b0000000000000000;
	sram_mem[117294] = 16'b0000000000000000;
	sram_mem[117295] = 16'b0000000000000000;
	sram_mem[117296] = 16'b0000000000000000;
	sram_mem[117297] = 16'b0000000000000000;
	sram_mem[117298] = 16'b0000000000000000;
	sram_mem[117299] = 16'b0000000000000000;
	sram_mem[117300] = 16'b0000000000000000;
	sram_mem[117301] = 16'b0000000000000000;
	sram_mem[117302] = 16'b0000000000000000;
	sram_mem[117303] = 16'b0000000000000000;
	sram_mem[117304] = 16'b0000000000000000;
	sram_mem[117305] = 16'b0000000000000000;
	sram_mem[117306] = 16'b0000000000000000;
	sram_mem[117307] = 16'b0000000000000000;
	sram_mem[117308] = 16'b0000000000000000;
	sram_mem[117309] = 16'b0000000000000000;
	sram_mem[117310] = 16'b0000000000000000;
	sram_mem[117311] = 16'b0000000000000000;
	sram_mem[117312] = 16'b0000000000000000;
	sram_mem[117313] = 16'b0000000000000000;
	sram_mem[117314] = 16'b0000000000000000;
	sram_mem[117315] = 16'b0000000000000000;
	sram_mem[117316] = 16'b0000000000000000;
	sram_mem[117317] = 16'b0000000000000000;
	sram_mem[117318] = 16'b0000000000000000;
	sram_mem[117319] = 16'b0000000000000000;
	sram_mem[117320] = 16'b0000000000000000;
	sram_mem[117321] = 16'b0000000000000000;
	sram_mem[117322] = 16'b0000000000000000;
	sram_mem[117323] = 16'b0000000000000000;
	sram_mem[117324] = 16'b0000000000000000;
	sram_mem[117325] = 16'b0000000000000000;
	sram_mem[117326] = 16'b0000000000000000;
	sram_mem[117327] = 16'b0000000000000000;
	sram_mem[117328] = 16'b0000000000000000;
	sram_mem[117329] = 16'b0000000000000000;
	sram_mem[117330] = 16'b0000000000000000;
	sram_mem[117331] = 16'b0000000000000000;
	sram_mem[117332] = 16'b0000000000000000;
	sram_mem[117333] = 16'b0000000000000000;
	sram_mem[117334] = 16'b0000000000000000;
	sram_mem[117335] = 16'b0000000000000000;
	sram_mem[117336] = 16'b0000000000000000;
	sram_mem[117337] = 16'b0000000000000000;
	sram_mem[117338] = 16'b0000000000000000;
	sram_mem[117339] = 16'b0000000000000000;
	sram_mem[117340] = 16'b0000000000000000;
	sram_mem[117341] = 16'b0000000000000000;
	sram_mem[117342] = 16'b0000000000000000;
	sram_mem[117343] = 16'b0000000000000000;
	sram_mem[117344] = 16'b0000000000000000;
	sram_mem[117345] = 16'b0000000000000000;
	sram_mem[117346] = 16'b0000000000000000;
	sram_mem[117347] = 16'b0000000000000000;
	sram_mem[117348] = 16'b0000000000000000;
	sram_mem[117349] = 16'b0000000000000000;
	sram_mem[117350] = 16'b0000000000000000;
	sram_mem[117351] = 16'b0000000000000000;
	sram_mem[117352] = 16'b0000000000000000;
	sram_mem[117353] = 16'b0000000000000000;
	sram_mem[117354] = 16'b0000000000000000;
	sram_mem[117355] = 16'b0000000000000000;
	sram_mem[117356] = 16'b0000000000000000;
	sram_mem[117357] = 16'b0000000000000000;
	sram_mem[117358] = 16'b0000000000000000;
	sram_mem[117359] = 16'b0000000000000000;
	sram_mem[117360] = 16'b0000000000000000;
	sram_mem[117361] = 16'b0000000000000000;
	sram_mem[117362] = 16'b0000000000000000;
	sram_mem[117363] = 16'b0000000000000000;
	sram_mem[117364] = 16'b0000000000000000;
	sram_mem[117365] = 16'b0000000000000000;
	sram_mem[117366] = 16'b0000000000000000;
	sram_mem[117367] = 16'b0000000000000000;
	sram_mem[117368] = 16'b0000000000000000;
	sram_mem[117369] = 16'b0000000000000000;
	sram_mem[117370] = 16'b0000000000000000;
	sram_mem[117371] = 16'b0000000000000000;
	sram_mem[117372] = 16'b0000000000000000;
	sram_mem[117373] = 16'b0000000000000000;
	sram_mem[117374] = 16'b0000000000000000;
	sram_mem[117375] = 16'b0000000000000000;
	sram_mem[117376] = 16'b0000000000000000;
	sram_mem[117377] = 16'b0000000000000000;
	sram_mem[117378] = 16'b0000000000000000;
	sram_mem[117379] = 16'b0000000000000000;
	sram_mem[117380] = 16'b0000000000000000;
	sram_mem[117381] = 16'b0000000000000000;
	sram_mem[117382] = 16'b0000000000000000;
	sram_mem[117383] = 16'b0000000000000000;
	sram_mem[117384] = 16'b0000000000000000;
	sram_mem[117385] = 16'b0000000000000000;
	sram_mem[117386] = 16'b0000000000000000;
	sram_mem[117387] = 16'b0000000000000000;
	sram_mem[117388] = 16'b0000000000000000;
	sram_mem[117389] = 16'b0000000000000000;
	sram_mem[117390] = 16'b0000000000000000;
	sram_mem[117391] = 16'b0000000000000000;
	sram_mem[117392] = 16'b0000000000000000;
	sram_mem[117393] = 16'b0000000000000000;
	sram_mem[117394] = 16'b0000000000000000;
	sram_mem[117395] = 16'b0000000000000000;
	sram_mem[117396] = 16'b0000000000000000;
	sram_mem[117397] = 16'b0000000000000000;
	sram_mem[117398] = 16'b0000000000000000;
	sram_mem[117399] = 16'b0000000000000000;
	sram_mem[117400] = 16'b0000000000000000;
	sram_mem[117401] = 16'b0000000000000000;
	sram_mem[117402] = 16'b0000000000000000;
	sram_mem[117403] = 16'b0000000000000000;
	sram_mem[117404] = 16'b0000000000000000;
	sram_mem[117405] = 16'b0000000000000000;
	sram_mem[117406] = 16'b0000000000000000;
	sram_mem[117407] = 16'b0000000000000000;
	sram_mem[117408] = 16'b0000000000000000;
	sram_mem[117409] = 16'b0000000000000000;
	sram_mem[117410] = 16'b0000000000000000;
	sram_mem[117411] = 16'b0000000000000000;
	sram_mem[117412] = 16'b0000000000000000;
	sram_mem[117413] = 16'b0000000000000000;
	sram_mem[117414] = 16'b0000000000000000;
	sram_mem[117415] = 16'b0000000000000000;
	sram_mem[117416] = 16'b0000000000000000;
	sram_mem[117417] = 16'b0000000000000000;
	sram_mem[117418] = 16'b0000000000000000;
	sram_mem[117419] = 16'b0000000000000000;
	sram_mem[117420] = 16'b0000000000000000;
	sram_mem[117421] = 16'b0000000000000000;
	sram_mem[117422] = 16'b0000000000000000;
	sram_mem[117423] = 16'b0000000000000000;
	sram_mem[117424] = 16'b0000000000000000;
	sram_mem[117425] = 16'b0000000000000000;
	sram_mem[117426] = 16'b0000000000000000;
	sram_mem[117427] = 16'b0000000000000000;
	sram_mem[117428] = 16'b0000000000000000;
	sram_mem[117429] = 16'b0000000000000000;
	sram_mem[117430] = 16'b0000000000000000;
	sram_mem[117431] = 16'b0000000000000000;
	sram_mem[117432] = 16'b0000000000000000;
	sram_mem[117433] = 16'b0000000000000000;
	sram_mem[117434] = 16'b0000000000000000;
	sram_mem[117435] = 16'b0000000000000000;
	sram_mem[117436] = 16'b0000000000000000;
	sram_mem[117437] = 16'b0000000000000000;
	sram_mem[117438] = 16'b0000000000000000;
	sram_mem[117439] = 16'b0000000000000000;
	sram_mem[117440] = 16'b0000000000000000;
	sram_mem[117441] = 16'b0000000000000000;
	sram_mem[117442] = 16'b0000000000000000;
	sram_mem[117443] = 16'b0000000000000000;
	sram_mem[117444] = 16'b0000000000000000;
	sram_mem[117445] = 16'b0000000000000000;
	sram_mem[117446] = 16'b0000000000000000;
	sram_mem[117447] = 16'b0000000000000000;
	sram_mem[117448] = 16'b0000000000000000;
	sram_mem[117449] = 16'b0000000000000000;
	sram_mem[117450] = 16'b0000000000000000;
	sram_mem[117451] = 16'b0000000000000000;
	sram_mem[117452] = 16'b0000000000000000;
	sram_mem[117453] = 16'b0000000000000000;
	sram_mem[117454] = 16'b0000000000000000;
	sram_mem[117455] = 16'b0000000000000000;
	sram_mem[117456] = 16'b0000000000000000;
	sram_mem[117457] = 16'b0000000000000000;
	sram_mem[117458] = 16'b0000000000000000;
	sram_mem[117459] = 16'b0000000000000000;
	sram_mem[117460] = 16'b0000000000000000;
	sram_mem[117461] = 16'b0000000000000000;
	sram_mem[117462] = 16'b0000000000000000;
	sram_mem[117463] = 16'b0000000000000000;
	sram_mem[117464] = 16'b0000000000000000;
	sram_mem[117465] = 16'b0000000000000000;
	sram_mem[117466] = 16'b0000000000000000;
	sram_mem[117467] = 16'b0000000000000000;
	sram_mem[117468] = 16'b0000000000000000;
	sram_mem[117469] = 16'b0000000000000000;
	sram_mem[117470] = 16'b0000000000000000;
	sram_mem[117471] = 16'b0000000000000000;
	sram_mem[117472] = 16'b0000000000000000;
	sram_mem[117473] = 16'b0000000000000000;
	sram_mem[117474] = 16'b0000000000000000;
	sram_mem[117475] = 16'b0000000000000000;
	sram_mem[117476] = 16'b0000000000000000;
	sram_mem[117477] = 16'b0000000000000000;
	sram_mem[117478] = 16'b0000000000000000;
	sram_mem[117479] = 16'b0000000000000000;
	sram_mem[117480] = 16'b0000000000000000;
	sram_mem[117481] = 16'b0000000000000000;
	sram_mem[117482] = 16'b0000000000000000;
	sram_mem[117483] = 16'b0000000000000000;
	sram_mem[117484] = 16'b0000000000000000;
	sram_mem[117485] = 16'b0000000000000000;
	sram_mem[117486] = 16'b0000000000000000;
	sram_mem[117487] = 16'b0000000000000000;
	sram_mem[117488] = 16'b0000000000000000;
	sram_mem[117489] = 16'b0000000000000000;
	sram_mem[117490] = 16'b0000000000000000;
	sram_mem[117491] = 16'b0000000000000000;
	sram_mem[117492] = 16'b0000000000000000;
	sram_mem[117493] = 16'b0000000000000000;
	sram_mem[117494] = 16'b0000000000000000;
	sram_mem[117495] = 16'b0000000000000000;
	sram_mem[117496] = 16'b0000000000000000;
	sram_mem[117497] = 16'b0000000000000000;
	sram_mem[117498] = 16'b0000000000000000;
	sram_mem[117499] = 16'b0000000000000000;
	sram_mem[117500] = 16'b0000000000000000;
	sram_mem[117501] = 16'b0000000000000000;
	sram_mem[117502] = 16'b0000000000000000;
	sram_mem[117503] = 16'b0000000000000000;
	sram_mem[117504] = 16'b0000000000000000;
	sram_mem[117505] = 16'b0000000000000000;
	sram_mem[117506] = 16'b0000000000000000;
	sram_mem[117507] = 16'b0000000000000000;
	sram_mem[117508] = 16'b0000000000000000;
	sram_mem[117509] = 16'b0000000000000000;
	sram_mem[117510] = 16'b0000000000000000;
	sram_mem[117511] = 16'b0000000000000000;
	sram_mem[117512] = 16'b0000000000000000;
	sram_mem[117513] = 16'b0000000000000000;
	sram_mem[117514] = 16'b0000000000000000;
	sram_mem[117515] = 16'b0000000000000000;
	sram_mem[117516] = 16'b0000000000000000;
	sram_mem[117517] = 16'b0000000000000000;
	sram_mem[117518] = 16'b0000000000000000;
	sram_mem[117519] = 16'b0000000000000000;
	sram_mem[117520] = 16'b0000000000000000;
	sram_mem[117521] = 16'b0000000000000000;
	sram_mem[117522] = 16'b0000000000000000;
	sram_mem[117523] = 16'b0000000000000000;
	sram_mem[117524] = 16'b0000000000000000;
	sram_mem[117525] = 16'b0000000000000000;
	sram_mem[117526] = 16'b0000000000000000;
	sram_mem[117527] = 16'b0000000000000000;
	sram_mem[117528] = 16'b0000000000000000;
	sram_mem[117529] = 16'b0000000000000000;
	sram_mem[117530] = 16'b0000000000000000;
	sram_mem[117531] = 16'b0000000000000000;
	sram_mem[117532] = 16'b0000000000000000;
	sram_mem[117533] = 16'b0000000000000000;
	sram_mem[117534] = 16'b0000000000000000;
	sram_mem[117535] = 16'b0000000000000000;
	sram_mem[117536] = 16'b0000000000000000;
	sram_mem[117537] = 16'b0000000000000000;
	sram_mem[117538] = 16'b0000000000000000;
	sram_mem[117539] = 16'b0000000000000000;
	sram_mem[117540] = 16'b0000000000000000;
	sram_mem[117541] = 16'b0000000000000000;
	sram_mem[117542] = 16'b0000000000000000;
	sram_mem[117543] = 16'b0000000000000000;
	sram_mem[117544] = 16'b0000000000000000;
	sram_mem[117545] = 16'b0000000000000000;
	sram_mem[117546] = 16'b0000000000000000;
	sram_mem[117547] = 16'b0000000000000000;
	sram_mem[117548] = 16'b0000000000000000;
	sram_mem[117549] = 16'b0000000000000000;
	sram_mem[117550] = 16'b0000000000000000;
	sram_mem[117551] = 16'b0000000000000000;
	sram_mem[117552] = 16'b0000000000000000;
	sram_mem[117553] = 16'b0000000000000000;
	sram_mem[117554] = 16'b0000000000000000;
	sram_mem[117555] = 16'b0000000000000000;
	sram_mem[117556] = 16'b0000000000000000;
	sram_mem[117557] = 16'b0000000000000000;
	sram_mem[117558] = 16'b0000000000000000;
	sram_mem[117559] = 16'b0000000000000000;
	sram_mem[117560] = 16'b0000000000000000;
	sram_mem[117561] = 16'b0000000000000000;
	sram_mem[117562] = 16'b0000000000000000;
	sram_mem[117563] = 16'b0000000000000000;
	sram_mem[117564] = 16'b0000000000000000;
	sram_mem[117565] = 16'b0000000000000000;
	sram_mem[117566] = 16'b0000000000000000;
	sram_mem[117567] = 16'b0000000000000000;
	sram_mem[117568] = 16'b0000000000000000;
	sram_mem[117569] = 16'b0000000000000000;
	sram_mem[117570] = 16'b0000000000000000;
	sram_mem[117571] = 16'b0000000000000000;
	sram_mem[117572] = 16'b0000000000000000;
	sram_mem[117573] = 16'b0000000000000000;
	sram_mem[117574] = 16'b0000000000000000;
	sram_mem[117575] = 16'b0000000000000000;
	sram_mem[117576] = 16'b0000000000000000;
	sram_mem[117577] = 16'b0000000000000000;
	sram_mem[117578] = 16'b0000000000000000;
	sram_mem[117579] = 16'b0000000000000000;
	sram_mem[117580] = 16'b0000000000000000;
	sram_mem[117581] = 16'b0000000000000000;
	sram_mem[117582] = 16'b0000000000000000;
	sram_mem[117583] = 16'b0000000000000000;
	sram_mem[117584] = 16'b0000000000000000;
	sram_mem[117585] = 16'b0000000000000000;
	sram_mem[117586] = 16'b0000000000000000;
	sram_mem[117587] = 16'b0000000000000000;
	sram_mem[117588] = 16'b0000000000000000;
	sram_mem[117589] = 16'b0000000000000000;
	sram_mem[117590] = 16'b0000000000000000;
	sram_mem[117591] = 16'b0000000000000000;
	sram_mem[117592] = 16'b0000000000000000;
	sram_mem[117593] = 16'b0000000000000000;
	sram_mem[117594] = 16'b0000000000000000;
	sram_mem[117595] = 16'b0000000000000000;
	sram_mem[117596] = 16'b0000000000000000;
	sram_mem[117597] = 16'b0000000000000000;
	sram_mem[117598] = 16'b0000000000000000;
	sram_mem[117599] = 16'b0000000000000000;
	sram_mem[117600] = 16'b0000000000000000;
	sram_mem[117601] = 16'b0000000000000000;
	sram_mem[117602] = 16'b0000000000000000;
	sram_mem[117603] = 16'b0000000000000000;
	sram_mem[117604] = 16'b0000000000000000;
	sram_mem[117605] = 16'b0000000000000000;
	sram_mem[117606] = 16'b0000000000000000;
	sram_mem[117607] = 16'b0000000000000000;
	sram_mem[117608] = 16'b0000000000000000;
	sram_mem[117609] = 16'b0000000000000000;
	sram_mem[117610] = 16'b0000000000000000;
	sram_mem[117611] = 16'b0000000000000000;
	sram_mem[117612] = 16'b0000000000000000;
	sram_mem[117613] = 16'b0000000000000000;
	sram_mem[117614] = 16'b0000000000000000;
	sram_mem[117615] = 16'b0000000000000000;
	sram_mem[117616] = 16'b0000000000000000;
	sram_mem[117617] = 16'b0000000000000000;
	sram_mem[117618] = 16'b0000000000000000;
	sram_mem[117619] = 16'b0000000000000000;
	sram_mem[117620] = 16'b0000000000000000;
	sram_mem[117621] = 16'b0000000000000000;
	sram_mem[117622] = 16'b0000000000000000;
	sram_mem[117623] = 16'b0000000000000000;
	sram_mem[117624] = 16'b0000000000000000;
	sram_mem[117625] = 16'b0000000000000000;
	sram_mem[117626] = 16'b0000000000000000;
	sram_mem[117627] = 16'b0000000000000000;
	sram_mem[117628] = 16'b0000000000000000;
	sram_mem[117629] = 16'b0000000000000000;
	sram_mem[117630] = 16'b0000000000000000;
	sram_mem[117631] = 16'b0000000000000000;
	sram_mem[117632] = 16'b0000000000000000;
	sram_mem[117633] = 16'b0000000000000000;
	sram_mem[117634] = 16'b0000000000000000;
	sram_mem[117635] = 16'b0000000000000000;
	sram_mem[117636] = 16'b0000000000000000;
	sram_mem[117637] = 16'b0000000000000000;
	sram_mem[117638] = 16'b0000000000000000;
	sram_mem[117639] = 16'b0000000000000000;
	sram_mem[117640] = 16'b0000000000000000;
	sram_mem[117641] = 16'b0000000000000000;
	sram_mem[117642] = 16'b0000000000000000;
	sram_mem[117643] = 16'b0000000000000000;
	sram_mem[117644] = 16'b0000000000000000;
	sram_mem[117645] = 16'b0000000000000000;
	sram_mem[117646] = 16'b0000000000000000;
	sram_mem[117647] = 16'b0000000000000000;
	sram_mem[117648] = 16'b0000000000000000;
	sram_mem[117649] = 16'b0000000000000000;
	sram_mem[117650] = 16'b0000000000000000;
	sram_mem[117651] = 16'b0000000000000000;
	sram_mem[117652] = 16'b0000000000000000;
	sram_mem[117653] = 16'b0000000000000000;
	sram_mem[117654] = 16'b0000000000000000;
	sram_mem[117655] = 16'b0000000000000000;
	sram_mem[117656] = 16'b0000000000000000;
	sram_mem[117657] = 16'b0000000000000000;
	sram_mem[117658] = 16'b0000000000000000;
	sram_mem[117659] = 16'b0000000000000000;
	sram_mem[117660] = 16'b0000000000000000;
	sram_mem[117661] = 16'b0000000000000000;
	sram_mem[117662] = 16'b0000000000000000;
	sram_mem[117663] = 16'b0000000000000000;
	sram_mem[117664] = 16'b0000000000000000;
	sram_mem[117665] = 16'b0000000000000000;
	sram_mem[117666] = 16'b0000000000000000;
	sram_mem[117667] = 16'b0000000000000000;
	sram_mem[117668] = 16'b0000000000000000;
	sram_mem[117669] = 16'b0000000000000000;
	sram_mem[117670] = 16'b0000000000000000;
	sram_mem[117671] = 16'b0000000000000000;
	sram_mem[117672] = 16'b0000000000000000;
	sram_mem[117673] = 16'b0000000000000000;
	sram_mem[117674] = 16'b0000000000000000;
	sram_mem[117675] = 16'b0000000000000000;
	sram_mem[117676] = 16'b0000000000000000;
	sram_mem[117677] = 16'b0000000000000000;
	sram_mem[117678] = 16'b0000000000000000;
	sram_mem[117679] = 16'b0000000000000000;
	sram_mem[117680] = 16'b0000000000000000;
	sram_mem[117681] = 16'b0000000000000000;
	sram_mem[117682] = 16'b0000000000000000;
	sram_mem[117683] = 16'b0000000000000000;
	sram_mem[117684] = 16'b0000000000000000;
	sram_mem[117685] = 16'b0000000000000000;
	sram_mem[117686] = 16'b0000000000000000;
	sram_mem[117687] = 16'b0000000000000000;
	sram_mem[117688] = 16'b0000000000000000;
	sram_mem[117689] = 16'b0000000000000000;
	sram_mem[117690] = 16'b0000000000000000;
	sram_mem[117691] = 16'b0000000000000000;
	sram_mem[117692] = 16'b0000000000000000;
	sram_mem[117693] = 16'b0000000000000000;
	sram_mem[117694] = 16'b0000000000000000;
	sram_mem[117695] = 16'b0000000000000000;
	sram_mem[117696] = 16'b0000000000000000;
	sram_mem[117697] = 16'b0000000000000000;
	sram_mem[117698] = 16'b0000000000000000;
	sram_mem[117699] = 16'b0000000000000000;
	sram_mem[117700] = 16'b0000000000000000;
	sram_mem[117701] = 16'b0000000000000000;
	sram_mem[117702] = 16'b0000000000000000;
	sram_mem[117703] = 16'b0000000000000000;
	sram_mem[117704] = 16'b0000000000000000;
	sram_mem[117705] = 16'b0000000000000000;
	sram_mem[117706] = 16'b0000000000000000;
	sram_mem[117707] = 16'b0000000000000000;
	sram_mem[117708] = 16'b0000000000000000;
	sram_mem[117709] = 16'b0000000000000000;
	sram_mem[117710] = 16'b0000000000000000;
	sram_mem[117711] = 16'b0000000000000000;
	sram_mem[117712] = 16'b0000000000000000;
	sram_mem[117713] = 16'b0000000000000000;
	sram_mem[117714] = 16'b0000000000000000;
	sram_mem[117715] = 16'b0000000000000000;
	sram_mem[117716] = 16'b0000000000000000;
	sram_mem[117717] = 16'b0000000000000000;
	sram_mem[117718] = 16'b0000000000000000;
	sram_mem[117719] = 16'b0000000000000000;
	sram_mem[117720] = 16'b0000000000000000;
	sram_mem[117721] = 16'b0000000000000000;
	sram_mem[117722] = 16'b0000000000000000;
	sram_mem[117723] = 16'b0000000000000000;
	sram_mem[117724] = 16'b0000000000000000;
	sram_mem[117725] = 16'b0000000000000000;
	sram_mem[117726] = 16'b0000000000000000;
	sram_mem[117727] = 16'b0000000000000000;
	sram_mem[117728] = 16'b0000000000000000;
	sram_mem[117729] = 16'b0000000000000000;
	sram_mem[117730] = 16'b0000000000000000;
	sram_mem[117731] = 16'b0000000000000000;
	sram_mem[117732] = 16'b0000000000000000;
	sram_mem[117733] = 16'b0000000000000000;
	sram_mem[117734] = 16'b0000000000000000;
	sram_mem[117735] = 16'b0000000000000000;
	sram_mem[117736] = 16'b0000000000000000;
	sram_mem[117737] = 16'b0000000000000000;
	sram_mem[117738] = 16'b0000000000000000;
	sram_mem[117739] = 16'b0000000000000000;
	sram_mem[117740] = 16'b0000000000000000;
	sram_mem[117741] = 16'b0000000000000000;
	sram_mem[117742] = 16'b0000000000000000;
	sram_mem[117743] = 16'b0000000000000000;
	sram_mem[117744] = 16'b0000000000000000;
	sram_mem[117745] = 16'b0000000000000000;
	sram_mem[117746] = 16'b0000000000000000;
	sram_mem[117747] = 16'b0000000000000000;
	sram_mem[117748] = 16'b0000000000000000;
	sram_mem[117749] = 16'b0000000000000000;
	sram_mem[117750] = 16'b0000000000000000;
	sram_mem[117751] = 16'b0000000000000000;
	sram_mem[117752] = 16'b0000000000000000;
	sram_mem[117753] = 16'b0000000000000000;
	sram_mem[117754] = 16'b0000000000000000;
	sram_mem[117755] = 16'b0000000000000000;
	sram_mem[117756] = 16'b0000000000000000;
	sram_mem[117757] = 16'b0000000000000000;
	sram_mem[117758] = 16'b0000000000000000;
	sram_mem[117759] = 16'b0000000000000000;
	sram_mem[117760] = 16'b0000000000000000;
	sram_mem[117761] = 16'b0000000000000000;
	sram_mem[117762] = 16'b0000000000000000;
	sram_mem[117763] = 16'b0000000000000000;
	sram_mem[117764] = 16'b0000000000000000;
	sram_mem[117765] = 16'b0000000000000000;
	sram_mem[117766] = 16'b0000000000000000;
	sram_mem[117767] = 16'b0000000000000000;
	sram_mem[117768] = 16'b0000000000000000;
	sram_mem[117769] = 16'b0000000000000000;
	sram_mem[117770] = 16'b0000000000000000;
	sram_mem[117771] = 16'b0000000000000000;
	sram_mem[117772] = 16'b0000000000000000;
	sram_mem[117773] = 16'b0000000000000000;
	sram_mem[117774] = 16'b0000000000000000;
	sram_mem[117775] = 16'b0000000000000000;
	sram_mem[117776] = 16'b0000000000000000;
	sram_mem[117777] = 16'b0000000000000000;
	sram_mem[117778] = 16'b0000000000000000;
	sram_mem[117779] = 16'b0000000000000000;
	sram_mem[117780] = 16'b0000000000000000;
	sram_mem[117781] = 16'b0000000000000000;
	sram_mem[117782] = 16'b0000000000000000;
	sram_mem[117783] = 16'b0000000000000000;
	sram_mem[117784] = 16'b0000000000000000;
	sram_mem[117785] = 16'b0000000000000000;
	sram_mem[117786] = 16'b0000000000000000;
	sram_mem[117787] = 16'b0000000000000000;
	sram_mem[117788] = 16'b0000000000000000;
	sram_mem[117789] = 16'b0000000000000000;
	sram_mem[117790] = 16'b0000000000000000;
	sram_mem[117791] = 16'b0000000000000000;
	sram_mem[117792] = 16'b0000000000000000;
	sram_mem[117793] = 16'b0000000000000000;
	sram_mem[117794] = 16'b0000000000000000;
	sram_mem[117795] = 16'b0000000000000000;
	sram_mem[117796] = 16'b0000000000000000;
	sram_mem[117797] = 16'b0000000000000000;
	sram_mem[117798] = 16'b0000000000000000;
	sram_mem[117799] = 16'b0000000000000000;
	sram_mem[117800] = 16'b0000000000000000;
	sram_mem[117801] = 16'b0000000000000000;
	sram_mem[117802] = 16'b0000000000000000;
	sram_mem[117803] = 16'b0000000000000000;
	sram_mem[117804] = 16'b0000000000000000;
	sram_mem[117805] = 16'b0000000000000000;
	sram_mem[117806] = 16'b0000000000000000;
	sram_mem[117807] = 16'b0000000000000000;
	sram_mem[117808] = 16'b0000000000000000;
	sram_mem[117809] = 16'b0000000000000000;
	sram_mem[117810] = 16'b0000000000000000;
	sram_mem[117811] = 16'b0000000000000000;
	sram_mem[117812] = 16'b0000000000000000;
	sram_mem[117813] = 16'b0000000000000000;
	sram_mem[117814] = 16'b0000000000000000;
	sram_mem[117815] = 16'b0000000000000000;
	sram_mem[117816] = 16'b0000000000000000;
	sram_mem[117817] = 16'b0000000000000000;
	sram_mem[117818] = 16'b0000000000000000;
	sram_mem[117819] = 16'b0000000000000000;
	sram_mem[117820] = 16'b0000000000000000;
	sram_mem[117821] = 16'b0000000000000000;
	sram_mem[117822] = 16'b0000000000000000;
	sram_mem[117823] = 16'b0000000000000000;
	sram_mem[117824] = 16'b0000000000000000;
	sram_mem[117825] = 16'b0000000000000000;
	sram_mem[117826] = 16'b0000000000000000;
	sram_mem[117827] = 16'b0000000000000000;
	sram_mem[117828] = 16'b0000000000000000;
	sram_mem[117829] = 16'b0000000000000000;
	sram_mem[117830] = 16'b0000000000000000;
	sram_mem[117831] = 16'b0000000000000000;
	sram_mem[117832] = 16'b0000000000000000;
	sram_mem[117833] = 16'b0000000000000000;
	sram_mem[117834] = 16'b0000000000000000;
	sram_mem[117835] = 16'b0000000000000000;
	sram_mem[117836] = 16'b0000000000000000;
	sram_mem[117837] = 16'b0000000000000000;
	sram_mem[117838] = 16'b0000000000000000;
	sram_mem[117839] = 16'b0000000000000000;
	sram_mem[117840] = 16'b0000000000000000;
	sram_mem[117841] = 16'b0000000000000000;
	sram_mem[117842] = 16'b0000000000000000;
	sram_mem[117843] = 16'b0000000000000000;
	sram_mem[117844] = 16'b0000000000000000;
	sram_mem[117845] = 16'b0000000000000000;
	sram_mem[117846] = 16'b0000000000000000;
	sram_mem[117847] = 16'b0000000000000000;
	sram_mem[117848] = 16'b0000000000000000;
	sram_mem[117849] = 16'b0000000000000000;
	sram_mem[117850] = 16'b0000000000000000;
	sram_mem[117851] = 16'b0000000000000000;
	sram_mem[117852] = 16'b0000000000000000;
	sram_mem[117853] = 16'b0000000000000000;
	sram_mem[117854] = 16'b0000000000000000;
	sram_mem[117855] = 16'b0000000000000000;
	sram_mem[117856] = 16'b0000000000000000;
	sram_mem[117857] = 16'b0000000000000000;
	sram_mem[117858] = 16'b0000000000000000;
	sram_mem[117859] = 16'b0000000000000000;
	sram_mem[117860] = 16'b0000000000000000;
	sram_mem[117861] = 16'b0000000000000000;
	sram_mem[117862] = 16'b0000000000000000;
	sram_mem[117863] = 16'b0000000000000000;
	sram_mem[117864] = 16'b0000000000000000;
	sram_mem[117865] = 16'b0000000000000000;
	sram_mem[117866] = 16'b0000000000000000;
	sram_mem[117867] = 16'b0000000000000000;
	sram_mem[117868] = 16'b0000000000000000;
	sram_mem[117869] = 16'b0000000000000000;
	sram_mem[117870] = 16'b0000000000000000;
	sram_mem[117871] = 16'b0000000000000000;
	sram_mem[117872] = 16'b0000000000000000;
	sram_mem[117873] = 16'b0000000000000000;
	sram_mem[117874] = 16'b0000000000000000;
	sram_mem[117875] = 16'b0000000000000000;
	sram_mem[117876] = 16'b0000000000000000;
	sram_mem[117877] = 16'b0000000000000000;
	sram_mem[117878] = 16'b0000000000000000;
	sram_mem[117879] = 16'b0000000000000000;
	sram_mem[117880] = 16'b0000000000000000;
	sram_mem[117881] = 16'b0000000000000000;
	sram_mem[117882] = 16'b0000000000000000;
	sram_mem[117883] = 16'b0000000000000000;
	sram_mem[117884] = 16'b0000000000000000;
	sram_mem[117885] = 16'b0000000000000000;
	sram_mem[117886] = 16'b0000000000000000;
	sram_mem[117887] = 16'b0000000000000000;
	sram_mem[117888] = 16'b0000000000000000;
	sram_mem[117889] = 16'b0000000000000000;
	sram_mem[117890] = 16'b0000000000000000;
	sram_mem[117891] = 16'b0000000000000000;
	sram_mem[117892] = 16'b0000000000000000;
	sram_mem[117893] = 16'b0000000000000000;
	sram_mem[117894] = 16'b0000000000000000;
	sram_mem[117895] = 16'b0000000000000000;
	sram_mem[117896] = 16'b0000000000000000;
	sram_mem[117897] = 16'b0000000000000000;
	sram_mem[117898] = 16'b0000000000000000;
	sram_mem[117899] = 16'b0000000000000000;
	sram_mem[117900] = 16'b0000000000000000;
	sram_mem[117901] = 16'b0000000000000000;
	sram_mem[117902] = 16'b0000000000000000;
	sram_mem[117903] = 16'b0000000000000000;
	sram_mem[117904] = 16'b0000000000000000;
	sram_mem[117905] = 16'b0000000000000000;
	sram_mem[117906] = 16'b0000000000000000;
	sram_mem[117907] = 16'b0000000000000000;
	sram_mem[117908] = 16'b0000000000000000;
	sram_mem[117909] = 16'b0000000000000000;
	sram_mem[117910] = 16'b0000000000000000;
	sram_mem[117911] = 16'b0000000000000000;
	sram_mem[117912] = 16'b0000000000000000;
	sram_mem[117913] = 16'b0000000000000000;
	sram_mem[117914] = 16'b0000000000000000;
	sram_mem[117915] = 16'b0000000000000000;
	sram_mem[117916] = 16'b0000000000000000;
	sram_mem[117917] = 16'b0000000000000000;
	sram_mem[117918] = 16'b0000000000000000;
	sram_mem[117919] = 16'b0000000000000000;
	sram_mem[117920] = 16'b0000000000000000;
	sram_mem[117921] = 16'b0000000000000000;
	sram_mem[117922] = 16'b0000000000000000;
	sram_mem[117923] = 16'b0000000000000000;
	sram_mem[117924] = 16'b0000000000000000;
	sram_mem[117925] = 16'b0000000000000000;
	sram_mem[117926] = 16'b0000000000000000;
	sram_mem[117927] = 16'b0000000000000000;
	sram_mem[117928] = 16'b0000000000000000;
	sram_mem[117929] = 16'b0000000000000000;
	sram_mem[117930] = 16'b0000000000000000;
	sram_mem[117931] = 16'b0000000000000000;
	sram_mem[117932] = 16'b0000000000000000;
	sram_mem[117933] = 16'b0000000000000000;
	sram_mem[117934] = 16'b0000000000000000;
	sram_mem[117935] = 16'b0000000000000000;
	sram_mem[117936] = 16'b0000000000000000;
	sram_mem[117937] = 16'b0000000000000000;
	sram_mem[117938] = 16'b0000000000000000;
	sram_mem[117939] = 16'b0000000000000000;
	sram_mem[117940] = 16'b0000000000000000;
	sram_mem[117941] = 16'b0000000000000000;
	sram_mem[117942] = 16'b0000000000000000;
	sram_mem[117943] = 16'b0000000000000000;
	sram_mem[117944] = 16'b0000000000000000;
	sram_mem[117945] = 16'b0000000000000000;
	sram_mem[117946] = 16'b0000000000000000;
	sram_mem[117947] = 16'b0000000000000000;
	sram_mem[117948] = 16'b0000000000000000;
	sram_mem[117949] = 16'b0000000000000000;
	sram_mem[117950] = 16'b0000000000000000;
	sram_mem[117951] = 16'b0000000000000000;
	sram_mem[117952] = 16'b0000000000000000;
	sram_mem[117953] = 16'b0000000000000000;
	sram_mem[117954] = 16'b0000000000000000;
	sram_mem[117955] = 16'b0000000000000000;
	sram_mem[117956] = 16'b0000000000000000;
	sram_mem[117957] = 16'b0000000000000000;
	sram_mem[117958] = 16'b0000000000000000;
	sram_mem[117959] = 16'b0000000000000000;
	sram_mem[117960] = 16'b0000000000000000;
	sram_mem[117961] = 16'b0000000000000000;
	sram_mem[117962] = 16'b0000000000000000;
	sram_mem[117963] = 16'b0000000000000000;
	sram_mem[117964] = 16'b0000000000000000;
	sram_mem[117965] = 16'b0000000000000000;
	sram_mem[117966] = 16'b0000000000000000;
	sram_mem[117967] = 16'b0000000000000000;
	sram_mem[117968] = 16'b0000000000000000;
	sram_mem[117969] = 16'b0000000000000000;
	sram_mem[117970] = 16'b0000000000000000;
	sram_mem[117971] = 16'b0000000000000000;
	sram_mem[117972] = 16'b0000000000000000;
	sram_mem[117973] = 16'b0000000000000000;
	sram_mem[117974] = 16'b0000000000000000;
	sram_mem[117975] = 16'b0000000000000000;
	sram_mem[117976] = 16'b0000000000000000;
	sram_mem[117977] = 16'b0000000000000000;
	sram_mem[117978] = 16'b0000000000000000;
	sram_mem[117979] = 16'b0000000000000000;
	sram_mem[117980] = 16'b0000000000000000;
	sram_mem[117981] = 16'b0000000000000000;
	sram_mem[117982] = 16'b0000000000000000;
	sram_mem[117983] = 16'b0000000000000000;
	sram_mem[117984] = 16'b0000000000000000;
	sram_mem[117985] = 16'b0000000000000000;
	sram_mem[117986] = 16'b0000000000000000;
	sram_mem[117987] = 16'b0000000000000000;
	sram_mem[117988] = 16'b0000000000000000;
	sram_mem[117989] = 16'b0000000000000000;
	sram_mem[117990] = 16'b0000000000000000;
	sram_mem[117991] = 16'b0000000000000000;
	sram_mem[117992] = 16'b0000000000000000;
	sram_mem[117993] = 16'b0000000000000000;
	sram_mem[117994] = 16'b0000000000000000;
	sram_mem[117995] = 16'b0000000000000000;
	sram_mem[117996] = 16'b0000000000000000;
	sram_mem[117997] = 16'b0000000000000000;
	sram_mem[117998] = 16'b0000000000000000;
	sram_mem[117999] = 16'b0000000000000000;
	sram_mem[118000] = 16'b0000000000000000;
	sram_mem[118001] = 16'b0000000000000000;
	sram_mem[118002] = 16'b0000000000000000;
	sram_mem[118003] = 16'b0000000000000000;
	sram_mem[118004] = 16'b0000000000000000;
	sram_mem[118005] = 16'b0000000000000000;
	sram_mem[118006] = 16'b0000000000000000;
	sram_mem[118007] = 16'b0000000000000000;
	sram_mem[118008] = 16'b0000000000000000;
	sram_mem[118009] = 16'b0000000000000000;
	sram_mem[118010] = 16'b0000000000000000;
	sram_mem[118011] = 16'b0000000000000000;
	sram_mem[118012] = 16'b0000000000000000;
	sram_mem[118013] = 16'b0000000000000000;
	sram_mem[118014] = 16'b0000000000000000;
	sram_mem[118015] = 16'b0000000000000000;
	sram_mem[118016] = 16'b0000000000000000;
	sram_mem[118017] = 16'b0000000000000000;
	sram_mem[118018] = 16'b0000000000000000;
	sram_mem[118019] = 16'b0000000000000000;
	sram_mem[118020] = 16'b0000000000000000;
	sram_mem[118021] = 16'b0000000000000000;
	sram_mem[118022] = 16'b0000000000000000;
	sram_mem[118023] = 16'b0000000000000000;
	sram_mem[118024] = 16'b0000000000000000;
	sram_mem[118025] = 16'b0000000000000000;
	sram_mem[118026] = 16'b0000000000000000;
	sram_mem[118027] = 16'b0000000000000000;
	sram_mem[118028] = 16'b0000000000000000;
	sram_mem[118029] = 16'b0000000000000000;
	sram_mem[118030] = 16'b0000000000000000;
	sram_mem[118031] = 16'b0000000000000000;
	sram_mem[118032] = 16'b0000000000000000;
	sram_mem[118033] = 16'b0000000000000000;
	sram_mem[118034] = 16'b0000000000000000;
	sram_mem[118035] = 16'b0000000000000000;
	sram_mem[118036] = 16'b0000000000000000;
	sram_mem[118037] = 16'b0000000000000000;
	sram_mem[118038] = 16'b0000000000000000;
	sram_mem[118039] = 16'b0000000000000000;
	sram_mem[118040] = 16'b0000000000000000;
	sram_mem[118041] = 16'b0000000000000000;
	sram_mem[118042] = 16'b0000000000000000;
	sram_mem[118043] = 16'b0000000000000000;
	sram_mem[118044] = 16'b0000000000000000;
	sram_mem[118045] = 16'b0000000000000000;
	sram_mem[118046] = 16'b0000000000000000;
	sram_mem[118047] = 16'b0000000000000000;
	sram_mem[118048] = 16'b0000000000000000;
	sram_mem[118049] = 16'b0000000000000000;
	sram_mem[118050] = 16'b0000000000000000;
	sram_mem[118051] = 16'b0000000000000000;
	sram_mem[118052] = 16'b0000000000000000;
	sram_mem[118053] = 16'b0000000000000000;
	sram_mem[118054] = 16'b0000000000000000;
	sram_mem[118055] = 16'b0000000000000000;
	sram_mem[118056] = 16'b0000000000000000;
	sram_mem[118057] = 16'b0000000000000000;
	sram_mem[118058] = 16'b0000000000000000;
	sram_mem[118059] = 16'b0000000000000000;
	sram_mem[118060] = 16'b0000000000000000;
	sram_mem[118061] = 16'b0000000000000000;
	sram_mem[118062] = 16'b0000000000000000;
	sram_mem[118063] = 16'b0000000000000000;
	sram_mem[118064] = 16'b0000000000000000;
	sram_mem[118065] = 16'b0000000000000000;
	sram_mem[118066] = 16'b0000000000000000;
	sram_mem[118067] = 16'b0000000000000000;
	sram_mem[118068] = 16'b0000000000000000;
	sram_mem[118069] = 16'b0000000000000000;
	sram_mem[118070] = 16'b0000000000000000;
	sram_mem[118071] = 16'b0000000000000000;
	sram_mem[118072] = 16'b0000000000000000;
	sram_mem[118073] = 16'b0000000000000000;
	sram_mem[118074] = 16'b0000000000000000;
	sram_mem[118075] = 16'b0000000000000000;
	sram_mem[118076] = 16'b0000000000000000;
	sram_mem[118077] = 16'b0000000000000000;
	sram_mem[118078] = 16'b0000000000000000;
	sram_mem[118079] = 16'b0000000000000000;
	sram_mem[118080] = 16'b0000000000000000;
	sram_mem[118081] = 16'b0000000000000000;
	sram_mem[118082] = 16'b0000000000000000;
	sram_mem[118083] = 16'b0000000000000000;
	sram_mem[118084] = 16'b0000000000000000;
	sram_mem[118085] = 16'b0000000000000000;
	sram_mem[118086] = 16'b0000000000000000;
	sram_mem[118087] = 16'b0000000000000000;
	sram_mem[118088] = 16'b0000000000000000;
	sram_mem[118089] = 16'b0000000000000000;
	sram_mem[118090] = 16'b0000000000000000;
	sram_mem[118091] = 16'b0000000000000000;
	sram_mem[118092] = 16'b0000000000000000;
	sram_mem[118093] = 16'b0000000000000000;
	sram_mem[118094] = 16'b0000000000000000;
	sram_mem[118095] = 16'b0000000000000000;
	sram_mem[118096] = 16'b0000000000000000;
	sram_mem[118097] = 16'b0000000000000000;
	sram_mem[118098] = 16'b0000000000000000;
	sram_mem[118099] = 16'b0000000000000000;
	sram_mem[118100] = 16'b0000000000000000;
	sram_mem[118101] = 16'b0000000000000000;
	sram_mem[118102] = 16'b0000000000000000;
	sram_mem[118103] = 16'b0000000000000000;
	sram_mem[118104] = 16'b0000000000000000;
	sram_mem[118105] = 16'b0000000000000000;
	sram_mem[118106] = 16'b0000000000000000;
	sram_mem[118107] = 16'b0000000000000000;
	sram_mem[118108] = 16'b0000000000000000;
	sram_mem[118109] = 16'b0000000000000000;
	sram_mem[118110] = 16'b0000000000000000;
	sram_mem[118111] = 16'b0000000000000000;
	sram_mem[118112] = 16'b0000000000000000;
	sram_mem[118113] = 16'b0000000000000000;
	sram_mem[118114] = 16'b0000000000000000;
	sram_mem[118115] = 16'b0000000000000000;
	sram_mem[118116] = 16'b0000000000000000;
	sram_mem[118117] = 16'b0000000000000000;
	sram_mem[118118] = 16'b0000000000000000;
	sram_mem[118119] = 16'b0000000000000000;
	sram_mem[118120] = 16'b0000000000000000;
	sram_mem[118121] = 16'b0000000000000000;
	sram_mem[118122] = 16'b0000000000000000;
	sram_mem[118123] = 16'b0000000000000000;
	sram_mem[118124] = 16'b0000000000000000;
	sram_mem[118125] = 16'b0000000000000000;
	sram_mem[118126] = 16'b0000000000000000;
	sram_mem[118127] = 16'b0000000000000000;
	sram_mem[118128] = 16'b0000000000000000;
	sram_mem[118129] = 16'b0000000000000000;
	sram_mem[118130] = 16'b0000000000000000;
	sram_mem[118131] = 16'b0000000000000000;
	sram_mem[118132] = 16'b0000000000000000;
	sram_mem[118133] = 16'b0000000000000000;
	sram_mem[118134] = 16'b0000000000000000;
	sram_mem[118135] = 16'b0000000000000000;
	sram_mem[118136] = 16'b0000000000000000;
	sram_mem[118137] = 16'b0000000000000000;
	sram_mem[118138] = 16'b0000000000000000;
	sram_mem[118139] = 16'b0000000000000000;
	sram_mem[118140] = 16'b0000000000000000;
	sram_mem[118141] = 16'b0000000000000000;
	sram_mem[118142] = 16'b0000000000000000;
	sram_mem[118143] = 16'b0000000000000000;
	sram_mem[118144] = 16'b0000000000000000;
	sram_mem[118145] = 16'b0000000000000000;
	sram_mem[118146] = 16'b0000000000000000;
	sram_mem[118147] = 16'b0000000000000000;
	sram_mem[118148] = 16'b0000000000000000;
	sram_mem[118149] = 16'b0000000000000000;
	sram_mem[118150] = 16'b0000000000000000;
	sram_mem[118151] = 16'b0000000000000000;
	sram_mem[118152] = 16'b0000000000000000;
	sram_mem[118153] = 16'b0000000000000000;
	sram_mem[118154] = 16'b0000000000000000;
	sram_mem[118155] = 16'b0000000000000000;
	sram_mem[118156] = 16'b0000000000000000;
	sram_mem[118157] = 16'b0000000000000000;
	sram_mem[118158] = 16'b0000000000000000;
	sram_mem[118159] = 16'b0000000000000000;
	sram_mem[118160] = 16'b0000000000000000;
	sram_mem[118161] = 16'b0000000000000000;
	sram_mem[118162] = 16'b0000000000000000;
	sram_mem[118163] = 16'b0000000000000000;
	sram_mem[118164] = 16'b0000000000000000;
	sram_mem[118165] = 16'b0000000000000000;
	sram_mem[118166] = 16'b0000000000000000;
	sram_mem[118167] = 16'b0000000000000000;
	sram_mem[118168] = 16'b0000000000000000;
	sram_mem[118169] = 16'b0000000000000000;
	sram_mem[118170] = 16'b0000000000000000;
	sram_mem[118171] = 16'b0000000000000000;
	sram_mem[118172] = 16'b0000000000000000;
	sram_mem[118173] = 16'b0000000000000000;
	sram_mem[118174] = 16'b0000000000000000;
	sram_mem[118175] = 16'b0000000000000000;
	sram_mem[118176] = 16'b0000000000000000;
	sram_mem[118177] = 16'b0000000000000000;
	sram_mem[118178] = 16'b0000000000000000;
	sram_mem[118179] = 16'b0000000000000000;
	sram_mem[118180] = 16'b0000000000000000;
	sram_mem[118181] = 16'b0000000000000000;
	sram_mem[118182] = 16'b0000000000000000;
	sram_mem[118183] = 16'b0000000000000000;
	sram_mem[118184] = 16'b0000000000000000;
	sram_mem[118185] = 16'b0000000000000000;
	sram_mem[118186] = 16'b0000000000000000;
	sram_mem[118187] = 16'b0000000000000000;
	sram_mem[118188] = 16'b0000000000000000;
	sram_mem[118189] = 16'b0000000000000000;
	sram_mem[118190] = 16'b0000000000000000;
	sram_mem[118191] = 16'b0000000000000000;
	sram_mem[118192] = 16'b0000000000000000;
	sram_mem[118193] = 16'b0000000000000000;
	sram_mem[118194] = 16'b0000000000000000;
	sram_mem[118195] = 16'b0000000000000000;
	sram_mem[118196] = 16'b0000000000000000;
	sram_mem[118197] = 16'b0000000000000000;
	sram_mem[118198] = 16'b0000000000000000;
	sram_mem[118199] = 16'b0000000000000000;
	sram_mem[118200] = 16'b0000000000000000;
	sram_mem[118201] = 16'b0000000000000000;
	sram_mem[118202] = 16'b0000000000000000;
	sram_mem[118203] = 16'b0000000000000000;
	sram_mem[118204] = 16'b0000000000000000;
	sram_mem[118205] = 16'b0000000000000000;
	sram_mem[118206] = 16'b0000000000000000;
	sram_mem[118207] = 16'b0000000000000000;
	sram_mem[118208] = 16'b0000000000000000;
	sram_mem[118209] = 16'b0000000000000000;
	sram_mem[118210] = 16'b0000000000000000;
	sram_mem[118211] = 16'b0000000000000000;
	sram_mem[118212] = 16'b0000000000000000;
	sram_mem[118213] = 16'b0000000000000000;
	sram_mem[118214] = 16'b0000000000000000;
	sram_mem[118215] = 16'b0000000000000000;
	sram_mem[118216] = 16'b0000000000000000;
	sram_mem[118217] = 16'b0000000000000000;
	sram_mem[118218] = 16'b0000000000000000;
	sram_mem[118219] = 16'b0000000000000000;
	sram_mem[118220] = 16'b0000000000000000;
	sram_mem[118221] = 16'b0000000000000000;
	sram_mem[118222] = 16'b0000000000000000;
	sram_mem[118223] = 16'b0000000000000000;
	sram_mem[118224] = 16'b0000000000000000;
	sram_mem[118225] = 16'b0000000000000000;
	sram_mem[118226] = 16'b0000000000000000;
	sram_mem[118227] = 16'b0000000000000000;
	sram_mem[118228] = 16'b0000000000000000;
	sram_mem[118229] = 16'b0000000000000000;
	sram_mem[118230] = 16'b0000000000000000;
	sram_mem[118231] = 16'b0000000000000000;
	sram_mem[118232] = 16'b0000000000000000;
	sram_mem[118233] = 16'b0000000000000000;
	sram_mem[118234] = 16'b0000000000000000;
	sram_mem[118235] = 16'b0000000000000000;
	sram_mem[118236] = 16'b0000000000000000;
	sram_mem[118237] = 16'b0000000000000000;
	sram_mem[118238] = 16'b0000000000000000;
	sram_mem[118239] = 16'b0000000000000000;
	sram_mem[118240] = 16'b0000000000000000;
	sram_mem[118241] = 16'b0000000000000000;
	sram_mem[118242] = 16'b0000000000000000;
	sram_mem[118243] = 16'b0000000000000000;
	sram_mem[118244] = 16'b0000000000000000;
	sram_mem[118245] = 16'b0000000000000000;
	sram_mem[118246] = 16'b0000000000000000;
	sram_mem[118247] = 16'b0000000000000000;
	sram_mem[118248] = 16'b0000000000000000;
	sram_mem[118249] = 16'b0000000000000000;
	sram_mem[118250] = 16'b0000000000000000;
	sram_mem[118251] = 16'b0000000000000000;
	sram_mem[118252] = 16'b0000000000000000;
	sram_mem[118253] = 16'b0000000000000000;
	sram_mem[118254] = 16'b0000000000000000;
	sram_mem[118255] = 16'b0000000000000000;
	sram_mem[118256] = 16'b0000000000000000;
	sram_mem[118257] = 16'b0000000000000000;
	sram_mem[118258] = 16'b0000000000000000;
	sram_mem[118259] = 16'b0000000000000000;
	sram_mem[118260] = 16'b0000000000000000;
	sram_mem[118261] = 16'b0000000000000000;
	sram_mem[118262] = 16'b0000000000000000;
	sram_mem[118263] = 16'b0000000000000000;
	sram_mem[118264] = 16'b0000000000000000;
	sram_mem[118265] = 16'b0000000000000000;
	sram_mem[118266] = 16'b0000000000000000;
	sram_mem[118267] = 16'b0000000000000000;
	sram_mem[118268] = 16'b0000000000000000;
	sram_mem[118269] = 16'b0000000000000000;
	sram_mem[118270] = 16'b0000000000000000;
	sram_mem[118271] = 16'b0000000000000000;
	sram_mem[118272] = 16'b0000000000000000;
	sram_mem[118273] = 16'b0000000000000000;
	sram_mem[118274] = 16'b0000000000000000;
	sram_mem[118275] = 16'b0000000000000000;
	sram_mem[118276] = 16'b0000000000000000;
	sram_mem[118277] = 16'b0000000000000000;
	sram_mem[118278] = 16'b0000000000000000;
	sram_mem[118279] = 16'b0000000000000000;
	sram_mem[118280] = 16'b0000000000000000;
	sram_mem[118281] = 16'b0000000000000000;
	sram_mem[118282] = 16'b0000000000000000;
	sram_mem[118283] = 16'b0000000000000000;
	sram_mem[118284] = 16'b0000000000000000;
	sram_mem[118285] = 16'b0000000000000000;
	sram_mem[118286] = 16'b0000000000000000;
	sram_mem[118287] = 16'b0000000000000000;
	sram_mem[118288] = 16'b0000000000000000;
	sram_mem[118289] = 16'b0000000000000000;
	sram_mem[118290] = 16'b0000000000000000;
	sram_mem[118291] = 16'b0000000000000000;
	sram_mem[118292] = 16'b0000000000000000;
	sram_mem[118293] = 16'b0000000000000000;
	sram_mem[118294] = 16'b0000000000000000;
	sram_mem[118295] = 16'b0000000000000000;
	sram_mem[118296] = 16'b0000000000000000;
	sram_mem[118297] = 16'b0000000000000000;
	sram_mem[118298] = 16'b0000000000000000;
	sram_mem[118299] = 16'b0000000000000000;
	sram_mem[118300] = 16'b0000000000000000;
	sram_mem[118301] = 16'b0000000000000000;
	sram_mem[118302] = 16'b0000000000000000;
	sram_mem[118303] = 16'b0000000000000000;
	sram_mem[118304] = 16'b0000000000000000;
	sram_mem[118305] = 16'b0000000000000000;
	sram_mem[118306] = 16'b0000000000000000;
	sram_mem[118307] = 16'b0000000000000000;
	sram_mem[118308] = 16'b0000000000000000;
	sram_mem[118309] = 16'b0000000000000000;
	sram_mem[118310] = 16'b0000000000000000;
	sram_mem[118311] = 16'b0000000000000000;
	sram_mem[118312] = 16'b0000000000000000;
	sram_mem[118313] = 16'b0000000000000000;
	sram_mem[118314] = 16'b0000000000000000;
	sram_mem[118315] = 16'b0000000000000000;
	sram_mem[118316] = 16'b0000000000000000;
	sram_mem[118317] = 16'b0000000000000000;
	sram_mem[118318] = 16'b0000000000000000;
	sram_mem[118319] = 16'b0000000000000000;
	sram_mem[118320] = 16'b0000000000000000;
	sram_mem[118321] = 16'b0000000000000000;
	sram_mem[118322] = 16'b0000000000000000;
	sram_mem[118323] = 16'b0000000000000000;
	sram_mem[118324] = 16'b0000000000000000;
	sram_mem[118325] = 16'b0000000000000000;
	sram_mem[118326] = 16'b0000000000000000;
	sram_mem[118327] = 16'b0000000000000000;
	sram_mem[118328] = 16'b0000000000000000;
	sram_mem[118329] = 16'b0000000000000000;
	sram_mem[118330] = 16'b0000000000000000;
	sram_mem[118331] = 16'b0000000000000000;
	sram_mem[118332] = 16'b0000000000000000;
	sram_mem[118333] = 16'b0000000000000000;
	sram_mem[118334] = 16'b0000000000000000;
	sram_mem[118335] = 16'b0000000000000000;
	sram_mem[118336] = 16'b0000000000000000;
	sram_mem[118337] = 16'b0000000000000000;
	sram_mem[118338] = 16'b0000000000000000;
	sram_mem[118339] = 16'b0000000000000000;
	sram_mem[118340] = 16'b0000000000000000;
	sram_mem[118341] = 16'b0000000000000000;
	sram_mem[118342] = 16'b0000000000000000;
	sram_mem[118343] = 16'b0000000000000000;
	sram_mem[118344] = 16'b0000000000000000;
	sram_mem[118345] = 16'b0000000000000000;
	sram_mem[118346] = 16'b0000000000000000;
	sram_mem[118347] = 16'b0000000000000000;
	sram_mem[118348] = 16'b0000000000000000;
	sram_mem[118349] = 16'b0000000000000000;
	sram_mem[118350] = 16'b0000000000000000;
	sram_mem[118351] = 16'b0000000000000000;
	sram_mem[118352] = 16'b0000000000000000;
	sram_mem[118353] = 16'b0000000000000000;
	sram_mem[118354] = 16'b0000000000000000;
	sram_mem[118355] = 16'b0000000000000000;
	sram_mem[118356] = 16'b0000000000000000;
	sram_mem[118357] = 16'b0000000000000000;
	sram_mem[118358] = 16'b0000000000000000;
	sram_mem[118359] = 16'b0000000000000000;
	sram_mem[118360] = 16'b0000000000000000;
	sram_mem[118361] = 16'b0000000000000000;
	sram_mem[118362] = 16'b0000000000000000;
	sram_mem[118363] = 16'b0000000000000000;
	sram_mem[118364] = 16'b0000000000000000;
	sram_mem[118365] = 16'b0000000000000000;
	sram_mem[118366] = 16'b0000000000000000;
	sram_mem[118367] = 16'b0000000000000000;
	sram_mem[118368] = 16'b0000000000000000;
	sram_mem[118369] = 16'b0000000000000000;
	sram_mem[118370] = 16'b0000000000000000;
	sram_mem[118371] = 16'b0000000000000000;
	sram_mem[118372] = 16'b0000000000000000;
	sram_mem[118373] = 16'b0000000000000000;
	sram_mem[118374] = 16'b0000000000000000;
	sram_mem[118375] = 16'b0000000000000000;
	sram_mem[118376] = 16'b0000000000000000;
	sram_mem[118377] = 16'b0000000000000000;
	sram_mem[118378] = 16'b0000000000000000;
	sram_mem[118379] = 16'b0000000000000000;
	sram_mem[118380] = 16'b0000000000000000;
	sram_mem[118381] = 16'b0000000000000000;
	sram_mem[118382] = 16'b0000000000000000;
	sram_mem[118383] = 16'b0000000000000000;
	sram_mem[118384] = 16'b0000000000000000;
	sram_mem[118385] = 16'b0000000000000000;
	sram_mem[118386] = 16'b0000000000000000;
	sram_mem[118387] = 16'b0000000000000000;
	sram_mem[118388] = 16'b0000000000000000;
	sram_mem[118389] = 16'b0000000000000000;
	sram_mem[118390] = 16'b0000000000000000;
	sram_mem[118391] = 16'b0000000000000000;
	sram_mem[118392] = 16'b0000000000000000;
	sram_mem[118393] = 16'b0000000000000000;
	sram_mem[118394] = 16'b0000000000000000;
	sram_mem[118395] = 16'b0000000000000000;
	sram_mem[118396] = 16'b0000000000000000;
	sram_mem[118397] = 16'b0000000000000000;
	sram_mem[118398] = 16'b0000000000000000;
	sram_mem[118399] = 16'b0000000000000000;
	sram_mem[118400] = 16'b0000000000000000;
	sram_mem[118401] = 16'b0000000000000000;
	sram_mem[118402] = 16'b0000000000000000;
	sram_mem[118403] = 16'b0000000000000000;
	sram_mem[118404] = 16'b0000000000000000;
	sram_mem[118405] = 16'b0000000000000000;
	sram_mem[118406] = 16'b0000000000000000;
	sram_mem[118407] = 16'b0000000000000000;
	sram_mem[118408] = 16'b0000000000000000;
	sram_mem[118409] = 16'b0000000000000000;
	sram_mem[118410] = 16'b0000000000000000;
	sram_mem[118411] = 16'b0000000000000000;
	sram_mem[118412] = 16'b0000000000000000;
	sram_mem[118413] = 16'b0000000000000000;
	sram_mem[118414] = 16'b0000000000000000;
	sram_mem[118415] = 16'b0000000000000000;
	sram_mem[118416] = 16'b0000000000000000;
	sram_mem[118417] = 16'b0000000000000000;
	sram_mem[118418] = 16'b0000000000000000;
	sram_mem[118419] = 16'b0000000000000000;
	sram_mem[118420] = 16'b0000000000000000;
	sram_mem[118421] = 16'b0000000000000000;
	sram_mem[118422] = 16'b0000000000000000;
	sram_mem[118423] = 16'b0000000000000000;
	sram_mem[118424] = 16'b0000000000000000;
	sram_mem[118425] = 16'b0000000000000000;
	sram_mem[118426] = 16'b0000000000000000;
	sram_mem[118427] = 16'b0000000000000000;
	sram_mem[118428] = 16'b0000000000000000;
	sram_mem[118429] = 16'b0000000000000000;
	sram_mem[118430] = 16'b0000000000000000;
	sram_mem[118431] = 16'b0000000000000000;
	sram_mem[118432] = 16'b0000000000000000;
	sram_mem[118433] = 16'b0000000000000000;
	sram_mem[118434] = 16'b0000000000000000;
	sram_mem[118435] = 16'b0000000000000000;
	sram_mem[118436] = 16'b0000000000000000;
	sram_mem[118437] = 16'b0000000000000000;
	sram_mem[118438] = 16'b0000000000000000;
	sram_mem[118439] = 16'b0000000000000000;
	sram_mem[118440] = 16'b0000000000000000;
	sram_mem[118441] = 16'b0000000000000000;
	sram_mem[118442] = 16'b0000000000000000;
	sram_mem[118443] = 16'b0000000000000000;
	sram_mem[118444] = 16'b0000000000000000;
	sram_mem[118445] = 16'b0000000000000000;
	sram_mem[118446] = 16'b0000000000000000;
	sram_mem[118447] = 16'b0000000000000000;
	sram_mem[118448] = 16'b0000000000000000;
	sram_mem[118449] = 16'b0000000000000000;
	sram_mem[118450] = 16'b0000000000000000;
	sram_mem[118451] = 16'b0000000000000000;
	sram_mem[118452] = 16'b0000000000000000;
	sram_mem[118453] = 16'b0000000000000000;
	sram_mem[118454] = 16'b0000000000000000;
	sram_mem[118455] = 16'b0000000000000000;
	sram_mem[118456] = 16'b0000000000000000;
	sram_mem[118457] = 16'b0000000000000000;
	sram_mem[118458] = 16'b0000000000000000;
	sram_mem[118459] = 16'b0000000000000000;
	sram_mem[118460] = 16'b0000000000000000;
	sram_mem[118461] = 16'b0000000000000000;
	sram_mem[118462] = 16'b0000000000000000;
	sram_mem[118463] = 16'b0000000000000000;
	sram_mem[118464] = 16'b0000000000000000;
	sram_mem[118465] = 16'b0000000000000000;
	sram_mem[118466] = 16'b0000000000000000;
	sram_mem[118467] = 16'b0000000000000000;
	sram_mem[118468] = 16'b0000000000000000;
	sram_mem[118469] = 16'b0000000000000000;
	sram_mem[118470] = 16'b0000000000000000;
	sram_mem[118471] = 16'b0000000000000000;
	sram_mem[118472] = 16'b0000000000000000;
	sram_mem[118473] = 16'b0000000000000000;
	sram_mem[118474] = 16'b0000000000000000;
	sram_mem[118475] = 16'b0000000000000000;
	sram_mem[118476] = 16'b0000000000000000;
	sram_mem[118477] = 16'b0000000000000000;
	sram_mem[118478] = 16'b0000000000000000;
	sram_mem[118479] = 16'b0000000000000000;
	sram_mem[118480] = 16'b0000000000000000;
	sram_mem[118481] = 16'b0000000000000000;
	sram_mem[118482] = 16'b0000000000000000;
	sram_mem[118483] = 16'b0000000000000000;
	sram_mem[118484] = 16'b0000000000000000;
	sram_mem[118485] = 16'b0000000000000000;
	sram_mem[118486] = 16'b0000000000000000;
	sram_mem[118487] = 16'b0000000000000000;
	sram_mem[118488] = 16'b0000000000000000;
	sram_mem[118489] = 16'b0000000000000000;
	sram_mem[118490] = 16'b0000000000000000;
	sram_mem[118491] = 16'b0000000000000000;
	sram_mem[118492] = 16'b0000000000000000;
	sram_mem[118493] = 16'b0000000000000000;
	sram_mem[118494] = 16'b0000000000000000;
	sram_mem[118495] = 16'b0000000000000000;
	sram_mem[118496] = 16'b0000000000000000;
	sram_mem[118497] = 16'b0000000000000000;
	sram_mem[118498] = 16'b0000000000000000;
	sram_mem[118499] = 16'b0000000000000000;
	sram_mem[118500] = 16'b0000000000000000;
	sram_mem[118501] = 16'b0000000000000000;
	sram_mem[118502] = 16'b0000000000000000;
	sram_mem[118503] = 16'b0000000000000000;
	sram_mem[118504] = 16'b0000000000000000;
	sram_mem[118505] = 16'b0000000000000000;
	sram_mem[118506] = 16'b0000000000000000;
	sram_mem[118507] = 16'b0000000000000000;
	sram_mem[118508] = 16'b0000000000000000;
	sram_mem[118509] = 16'b0000000000000000;
	sram_mem[118510] = 16'b0000000000000000;
	sram_mem[118511] = 16'b0000000000000000;
	sram_mem[118512] = 16'b0000000000000000;
	sram_mem[118513] = 16'b0000000000000000;
	sram_mem[118514] = 16'b0000000000000000;
	sram_mem[118515] = 16'b0000000000000000;
	sram_mem[118516] = 16'b0000000000000000;
	sram_mem[118517] = 16'b0000000000000000;
	sram_mem[118518] = 16'b0000000000000000;
	sram_mem[118519] = 16'b0000000000000000;
	sram_mem[118520] = 16'b0000000000000000;
	sram_mem[118521] = 16'b0000000000000000;
	sram_mem[118522] = 16'b0000000000000000;
	sram_mem[118523] = 16'b0000000000000000;
	sram_mem[118524] = 16'b0000000000000000;
	sram_mem[118525] = 16'b0000000000000000;
	sram_mem[118526] = 16'b0000000000000000;
	sram_mem[118527] = 16'b0000000000000000;
	sram_mem[118528] = 16'b0000000000000000;
	sram_mem[118529] = 16'b0000000000000000;
	sram_mem[118530] = 16'b0000000000000000;
	sram_mem[118531] = 16'b0000000000000000;
	sram_mem[118532] = 16'b0000000000000000;
	sram_mem[118533] = 16'b0000000000000000;
	sram_mem[118534] = 16'b0000000000000000;
	sram_mem[118535] = 16'b0000000000000000;
	sram_mem[118536] = 16'b0000000000000000;
	sram_mem[118537] = 16'b0000000000000000;
	sram_mem[118538] = 16'b0000000000000000;
	sram_mem[118539] = 16'b0000000000000000;
	sram_mem[118540] = 16'b0000000000000000;
	sram_mem[118541] = 16'b0000000000000000;
	sram_mem[118542] = 16'b0000000000000000;
	sram_mem[118543] = 16'b0000000000000000;
	sram_mem[118544] = 16'b0000000000000000;
	sram_mem[118545] = 16'b0000000000000000;
	sram_mem[118546] = 16'b0000000000000000;
	sram_mem[118547] = 16'b0000000000000000;
	sram_mem[118548] = 16'b0000000000000000;
	sram_mem[118549] = 16'b0000000000000000;
	sram_mem[118550] = 16'b0000000000000000;
	sram_mem[118551] = 16'b0000000000000000;
	sram_mem[118552] = 16'b0000000000000000;
	sram_mem[118553] = 16'b0000000000000000;
	sram_mem[118554] = 16'b0000000000000000;
	sram_mem[118555] = 16'b0000000000000000;
	sram_mem[118556] = 16'b0000000000000000;
	sram_mem[118557] = 16'b0000000000000000;
	sram_mem[118558] = 16'b0000000000000000;
	sram_mem[118559] = 16'b0000000000000000;
	sram_mem[118560] = 16'b0000000000000000;
	sram_mem[118561] = 16'b0000000000000000;
	sram_mem[118562] = 16'b0000000000000000;
	sram_mem[118563] = 16'b0000000000000000;
	sram_mem[118564] = 16'b0000000000000000;
	sram_mem[118565] = 16'b0000000000000000;
	sram_mem[118566] = 16'b0000000000000000;
	sram_mem[118567] = 16'b0000000000000000;
	sram_mem[118568] = 16'b0000000000000000;
	sram_mem[118569] = 16'b0000000000000000;
	sram_mem[118570] = 16'b0000000000000000;
	sram_mem[118571] = 16'b0000000000000000;
	sram_mem[118572] = 16'b0000000000000000;
	sram_mem[118573] = 16'b0000000000000000;
	sram_mem[118574] = 16'b0000000000000000;
	sram_mem[118575] = 16'b0000000000000000;
	sram_mem[118576] = 16'b0000000000000000;
	sram_mem[118577] = 16'b0000000000000000;
	sram_mem[118578] = 16'b0000000000000000;
	sram_mem[118579] = 16'b0000000000000000;
	sram_mem[118580] = 16'b0000000000000000;
	sram_mem[118581] = 16'b0000000000000000;
	sram_mem[118582] = 16'b0000000000000000;
	sram_mem[118583] = 16'b0000000000000000;
	sram_mem[118584] = 16'b0000000000000000;
	sram_mem[118585] = 16'b0000000000000000;
	sram_mem[118586] = 16'b0000000000000000;
	sram_mem[118587] = 16'b0000000000000000;
	sram_mem[118588] = 16'b0000000000000000;
	sram_mem[118589] = 16'b0000000000000000;
	sram_mem[118590] = 16'b0000000000000000;
	sram_mem[118591] = 16'b0000000000000000;
	sram_mem[118592] = 16'b0000000000000000;
	sram_mem[118593] = 16'b0000000000000000;
	sram_mem[118594] = 16'b0000000000000000;
	sram_mem[118595] = 16'b0000000000000000;
	sram_mem[118596] = 16'b0000000000000000;
	sram_mem[118597] = 16'b0000000000000000;
	sram_mem[118598] = 16'b0000000000000000;
	sram_mem[118599] = 16'b0000000000000000;
	sram_mem[118600] = 16'b0000000000000000;
	sram_mem[118601] = 16'b0000000000000000;
	sram_mem[118602] = 16'b0000000000000000;
	sram_mem[118603] = 16'b0000000000000000;
	sram_mem[118604] = 16'b0000000000000000;
	sram_mem[118605] = 16'b0000000000000000;
	sram_mem[118606] = 16'b0000000000000000;
	sram_mem[118607] = 16'b0000000000000000;
	sram_mem[118608] = 16'b0000000000000000;
	sram_mem[118609] = 16'b0000000000000000;
	sram_mem[118610] = 16'b0000000000000000;
	sram_mem[118611] = 16'b0000000000000000;
	sram_mem[118612] = 16'b0000000000000000;
	sram_mem[118613] = 16'b0000000000000000;
	sram_mem[118614] = 16'b0000000000000000;
	sram_mem[118615] = 16'b0000000000000000;
	sram_mem[118616] = 16'b0000000000000000;
	sram_mem[118617] = 16'b0000000000000000;
	sram_mem[118618] = 16'b0000000000000000;
	sram_mem[118619] = 16'b0000000000000000;
	sram_mem[118620] = 16'b0000000000000000;
	sram_mem[118621] = 16'b0000000000000000;
	sram_mem[118622] = 16'b0000000000000000;
	sram_mem[118623] = 16'b0000000000000000;
	sram_mem[118624] = 16'b0000000000000000;
	sram_mem[118625] = 16'b0000000000000000;
	sram_mem[118626] = 16'b0000000000000000;
	sram_mem[118627] = 16'b0000000000000000;
	sram_mem[118628] = 16'b0000000000000000;
	sram_mem[118629] = 16'b0000000000000000;
	sram_mem[118630] = 16'b0000000000000000;
	sram_mem[118631] = 16'b0000000000000000;
	sram_mem[118632] = 16'b0000000000000000;
	sram_mem[118633] = 16'b0000000000000000;
	sram_mem[118634] = 16'b0000000000000000;
	sram_mem[118635] = 16'b0000000000000000;
	sram_mem[118636] = 16'b0000000000000000;
	sram_mem[118637] = 16'b0000000000000000;
	sram_mem[118638] = 16'b0000000000000000;
	sram_mem[118639] = 16'b0000000000000000;
	sram_mem[118640] = 16'b0000000000000000;
	sram_mem[118641] = 16'b0000000000000000;
	sram_mem[118642] = 16'b0000000000000000;
	sram_mem[118643] = 16'b0000000000000000;
	sram_mem[118644] = 16'b0000000000000000;
	sram_mem[118645] = 16'b0000000000000000;
	sram_mem[118646] = 16'b0000000000000000;
	sram_mem[118647] = 16'b0000000000000000;
	sram_mem[118648] = 16'b0000000000000000;
	sram_mem[118649] = 16'b0000000000000000;
	sram_mem[118650] = 16'b0000000000000000;
	sram_mem[118651] = 16'b0000000000000000;
	sram_mem[118652] = 16'b0000000000000000;
	sram_mem[118653] = 16'b0000000000000000;
	sram_mem[118654] = 16'b0000000000000000;
	sram_mem[118655] = 16'b0000000000000000;
	sram_mem[118656] = 16'b0000000000000000;
	sram_mem[118657] = 16'b0000000000000000;
	sram_mem[118658] = 16'b0000000000000000;
	sram_mem[118659] = 16'b0000000000000000;
	sram_mem[118660] = 16'b0000000000000000;
	sram_mem[118661] = 16'b0000000000000000;
	sram_mem[118662] = 16'b0000000000000000;
	sram_mem[118663] = 16'b0000000000000000;
	sram_mem[118664] = 16'b0000000000000000;
	sram_mem[118665] = 16'b0000000000000000;
	sram_mem[118666] = 16'b0000000000000000;
	sram_mem[118667] = 16'b0000000000000000;
	sram_mem[118668] = 16'b0000000000000000;
	sram_mem[118669] = 16'b0000000000000000;
	sram_mem[118670] = 16'b0000000000000000;
	sram_mem[118671] = 16'b0000000000000000;
	sram_mem[118672] = 16'b0000000000000000;
	sram_mem[118673] = 16'b0000000000000000;
	sram_mem[118674] = 16'b0000000000000000;
	sram_mem[118675] = 16'b0000000000000000;
	sram_mem[118676] = 16'b0000000000000000;
	sram_mem[118677] = 16'b0000000000000000;
	sram_mem[118678] = 16'b0000000000000000;
	sram_mem[118679] = 16'b0000000000000000;
	sram_mem[118680] = 16'b0000000000000000;
	sram_mem[118681] = 16'b0000000000000000;
	sram_mem[118682] = 16'b0000000000000000;
	sram_mem[118683] = 16'b0000000000000000;
	sram_mem[118684] = 16'b0000000000000000;
	sram_mem[118685] = 16'b0000000000000000;
	sram_mem[118686] = 16'b0000000000000000;
	sram_mem[118687] = 16'b0000000000000000;
	sram_mem[118688] = 16'b0000000000000000;
	sram_mem[118689] = 16'b0000000000000000;
	sram_mem[118690] = 16'b0000000000000000;
	sram_mem[118691] = 16'b0000000000000000;
	sram_mem[118692] = 16'b0000000000000000;
	sram_mem[118693] = 16'b0000000000000000;
	sram_mem[118694] = 16'b0000000000000000;
	sram_mem[118695] = 16'b0000000000000000;
	sram_mem[118696] = 16'b0000000000000000;
	sram_mem[118697] = 16'b0000000000000000;
	sram_mem[118698] = 16'b0000000000000000;
	sram_mem[118699] = 16'b0000000000000000;
	sram_mem[118700] = 16'b0000000000000000;
	sram_mem[118701] = 16'b0000000000000000;
	sram_mem[118702] = 16'b0000000000000000;
	sram_mem[118703] = 16'b0000000000000000;
	sram_mem[118704] = 16'b0000000000000000;
	sram_mem[118705] = 16'b0000000000000000;
	sram_mem[118706] = 16'b0000000000000000;
	sram_mem[118707] = 16'b0000000000000000;
	sram_mem[118708] = 16'b0000000000000000;
	sram_mem[118709] = 16'b0000000000000000;
	sram_mem[118710] = 16'b0000000000000000;
	sram_mem[118711] = 16'b0000000000000000;
	sram_mem[118712] = 16'b0000000000000000;
	sram_mem[118713] = 16'b0000000000000000;
	sram_mem[118714] = 16'b0000000000000000;
	sram_mem[118715] = 16'b0000000000000000;
	sram_mem[118716] = 16'b0000000000000000;
	sram_mem[118717] = 16'b0000000000000000;
	sram_mem[118718] = 16'b0000000000000000;
	sram_mem[118719] = 16'b0000000000000000;
	sram_mem[118720] = 16'b0000000000000000;
	sram_mem[118721] = 16'b0000000000000000;
	sram_mem[118722] = 16'b0000000000000000;
	sram_mem[118723] = 16'b0000000000000000;
	sram_mem[118724] = 16'b0000000000000000;
	sram_mem[118725] = 16'b0000000000000000;
	sram_mem[118726] = 16'b0000000000000000;
	sram_mem[118727] = 16'b0000000000000000;
	sram_mem[118728] = 16'b0000000000000000;
	sram_mem[118729] = 16'b0000000000000000;
	sram_mem[118730] = 16'b0000000000000000;
	sram_mem[118731] = 16'b0000000000000000;
	sram_mem[118732] = 16'b0000000000000000;
	sram_mem[118733] = 16'b0000000000000000;
	sram_mem[118734] = 16'b0000000000000000;
	sram_mem[118735] = 16'b0000000000000000;
	sram_mem[118736] = 16'b0000000000000000;
	sram_mem[118737] = 16'b0000000000000000;
	sram_mem[118738] = 16'b0000000000000000;
	sram_mem[118739] = 16'b0000000000000000;
	sram_mem[118740] = 16'b0000000000000000;
	sram_mem[118741] = 16'b0000000000000000;
	sram_mem[118742] = 16'b0000000000000000;
	sram_mem[118743] = 16'b0000000000000000;
	sram_mem[118744] = 16'b0000000000000000;
	sram_mem[118745] = 16'b0000000000000000;
	sram_mem[118746] = 16'b0000000000000000;
	sram_mem[118747] = 16'b0000000000000000;
	sram_mem[118748] = 16'b0000000000000000;
	sram_mem[118749] = 16'b0000000000000000;
	sram_mem[118750] = 16'b0000000000000000;
	sram_mem[118751] = 16'b0000000000000000;
	sram_mem[118752] = 16'b0000000000000000;
	sram_mem[118753] = 16'b0000000000000000;
	sram_mem[118754] = 16'b0000000000000000;
	sram_mem[118755] = 16'b0000000000000000;
	sram_mem[118756] = 16'b0000000000000000;
	sram_mem[118757] = 16'b0000000000000000;
	sram_mem[118758] = 16'b0000000000000000;
	sram_mem[118759] = 16'b0000000000000000;
	sram_mem[118760] = 16'b0000000000000000;
	sram_mem[118761] = 16'b0000000000000000;
	sram_mem[118762] = 16'b0000000000000000;
	sram_mem[118763] = 16'b0000000000000000;
	sram_mem[118764] = 16'b0000000000000000;
	sram_mem[118765] = 16'b0000000000000000;
	sram_mem[118766] = 16'b0000000000000000;
	sram_mem[118767] = 16'b0000000000000000;
	sram_mem[118768] = 16'b0000000000000000;
	sram_mem[118769] = 16'b0000000000000000;
	sram_mem[118770] = 16'b0000000000000000;
	sram_mem[118771] = 16'b0000000000000000;
	sram_mem[118772] = 16'b0000000000000000;
	sram_mem[118773] = 16'b0000000000000000;
	sram_mem[118774] = 16'b0000000000000000;
	sram_mem[118775] = 16'b0000000000000000;
	sram_mem[118776] = 16'b0000000000000000;
	sram_mem[118777] = 16'b0000000000000000;
	sram_mem[118778] = 16'b0000000000000000;
	sram_mem[118779] = 16'b0000000000000000;
	sram_mem[118780] = 16'b0000000000000000;
	sram_mem[118781] = 16'b0000000000000000;
	sram_mem[118782] = 16'b0000000000000000;
	sram_mem[118783] = 16'b0000000000000000;
	sram_mem[118784] = 16'b0000000000000000;
	sram_mem[118785] = 16'b0000000000000000;
	sram_mem[118786] = 16'b0000000000000000;
	sram_mem[118787] = 16'b0000000000000000;
	sram_mem[118788] = 16'b0000000000000000;
	sram_mem[118789] = 16'b0000000000000000;
	sram_mem[118790] = 16'b0000000000000000;
	sram_mem[118791] = 16'b0000000000000000;
	sram_mem[118792] = 16'b0000000000000000;
	sram_mem[118793] = 16'b0000000000000000;
	sram_mem[118794] = 16'b0000000000000000;
	sram_mem[118795] = 16'b0000000000000000;
	sram_mem[118796] = 16'b0000000000000000;
	sram_mem[118797] = 16'b0000000000000000;
	sram_mem[118798] = 16'b0000000000000000;
	sram_mem[118799] = 16'b0000000000000000;
	sram_mem[118800] = 16'b0000000000000000;
	sram_mem[118801] = 16'b0000000000000000;
	sram_mem[118802] = 16'b0000000000000000;
	sram_mem[118803] = 16'b0000000000000000;
	sram_mem[118804] = 16'b0000000000000000;
	sram_mem[118805] = 16'b0000000000000000;
	sram_mem[118806] = 16'b0000000000000000;
	sram_mem[118807] = 16'b0000000000000000;
	sram_mem[118808] = 16'b0000000000000000;
	sram_mem[118809] = 16'b0000000000000000;
	sram_mem[118810] = 16'b0000000000000000;
	sram_mem[118811] = 16'b0000000000000000;
	sram_mem[118812] = 16'b0000000000000000;
	sram_mem[118813] = 16'b0000000000000000;
	sram_mem[118814] = 16'b0000000000000000;
	sram_mem[118815] = 16'b0000000000000000;
	sram_mem[118816] = 16'b0000000000000000;
	sram_mem[118817] = 16'b0000000000000000;
	sram_mem[118818] = 16'b0000000000000000;
	sram_mem[118819] = 16'b0000000000000000;
	sram_mem[118820] = 16'b0000000000000000;
	sram_mem[118821] = 16'b0000000000000000;
	sram_mem[118822] = 16'b0000000000000000;
	sram_mem[118823] = 16'b0000000000000000;
	sram_mem[118824] = 16'b0000000000000000;
	sram_mem[118825] = 16'b0000000000000000;
	sram_mem[118826] = 16'b0000000000000000;
	sram_mem[118827] = 16'b0000000000000000;
	sram_mem[118828] = 16'b0000000000000000;
	sram_mem[118829] = 16'b0000000000000000;
	sram_mem[118830] = 16'b0000000000000000;
	sram_mem[118831] = 16'b0000000000000000;
	sram_mem[118832] = 16'b0000000000000000;
	sram_mem[118833] = 16'b0000000000000000;
	sram_mem[118834] = 16'b0000000000000000;
	sram_mem[118835] = 16'b0000000000000000;
	sram_mem[118836] = 16'b0000000000000000;
	sram_mem[118837] = 16'b0000000000000000;
	sram_mem[118838] = 16'b0000000000000000;
	sram_mem[118839] = 16'b0000000000000000;
	sram_mem[118840] = 16'b0000000000000000;
	sram_mem[118841] = 16'b0000000000000000;
	sram_mem[118842] = 16'b0000000000000000;
	sram_mem[118843] = 16'b0000000000000000;
	sram_mem[118844] = 16'b0000000000000000;
	sram_mem[118845] = 16'b0000000000000000;
	sram_mem[118846] = 16'b0000000000000000;
	sram_mem[118847] = 16'b0000000000000000;
	sram_mem[118848] = 16'b0000000000000000;
	sram_mem[118849] = 16'b0000000000000000;
	sram_mem[118850] = 16'b0000000000000000;
	sram_mem[118851] = 16'b0000000000000000;
	sram_mem[118852] = 16'b0000000000000000;
	sram_mem[118853] = 16'b0000000000000000;
	sram_mem[118854] = 16'b0000000000000000;
	sram_mem[118855] = 16'b0000000000000000;
	sram_mem[118856] = 16'b0000000000000000;
	sram_mem[118857] = 16'b0000000000000000;
	sram_mem[118858] = 16'b0000000000000000;
	sram_mem[118859] = 16'b0000000000000000;
	sram_mem[118860] = 16'b0000000000000000;
	sram_mem[118861] = 16'b0000000000000000;
	sram_mem[118862] = 16'b0000000000000000;
	sram_mem[118863] = 16'b0000000000000000;
	sram_mem[118864] = 16'b0000000000000000;
	sram_mem[118865] = 16'b0000000000000000;
	sram_mem[118866] = 16'b0000000000000000;
	sram_mem[118867] = 16'b0000000000000000;
	sram_mem[118868] = 16'b0000000000000000;
	sram_mem[118869] = 16'b0000000000000000;
	sram_mem[118870] = 16'b0000000000000000;
	sram_mem[118871] = 16'b0000000000000000;
	sram_mem[118872] = 16'b0000000000000000;
	sram_mem[118873] = 16'b0000000000000000;
	sram_mem[118874] = 16'b0000000000000000;
	sram_mem[118875] = 16'b0000000000000000;
	sram_mem[118876] = 16'b0000000000000000;
	sram_mem[118877] = 16'b0000000000000000;
	sram_mem[118878] = 16'b0000000000000000;
	sram_mem[118879] = 16'b0000000000000000;
	sram_mem[118880] = 16'b0000000000000000;
	sram_mem[118881] = 16'b0000000000000000;
	sram_mem[118882] = 16'b0000000000000000;
	sram_mem[118883] = 16'b0000000000000000;
	sram_mem[118884] = 16'b0000000000000000;
	sram_mem[118885] = 16'b0000000000000000;
	sram_mem[118886] = 16'b0000000000000000;
	sram_mem[118887] = 16'b0000000000000000;
	sram_mem[118888] = 16'b0000000000000000;
	sram_mem[118889] = 16'b0000000000000000;
	sram_mem[118890] = 16'b0000000000000000;
	sram_mem[118891] = 16'b0000000000000000;
	sram_mem[118892] = 16'b0000000000000000;
	sram_mem[118893] = 16'b0000000000000000;
	sram_mem[118894] = 16'b0000000000000000;
	sram_mem[118895] = 16'b0000000000000000;
	sram_mem[118896] = 16'b0000000000000000;
	sram_mem[118897] = 16'b0000000000000000;
	sram_mem[118898] = 16'b0000000000000000;
	sram_mem[118899] = 16'b0000000000000000;
	sram_mem[118900] = 16'b0000000000000000;
	sram_mem[118901] = 16'b0000000000000000;
	sram_mem[118902] = 16'b0000000000000000;
	sram_mem[118903] = 16'b0000000000000000;
	sram_mem[118904] = 16'b0000000000000000;
	sram_mem[118905] = 16'b0000000000000000;
	sram_mem[118906] = 16'b0000000000000000;
	sram_mem[118907] = 16'b0000000000000000;
	sram_mem[118908] = 16'b0000000000000000;
	sram_mem[118909] = 16'b0000000000000000;
	sram_mem[118910] = 16'b0000000000000000;
	sram_mem[118911] = 16'b0000000000000000;
	sram_mem[118912] = 16'b0000000000000000;
	sram_mem[118913] = 16'b0000000000000000;
	sram_mem[118914] = 16'b0000000000000000;
	sram_mem[118915] = 16'b0000000000000000;
	sram_mem[118916] = 16'b0000000000000000;
	sram_mem[118917] = 16'b0000000000000000;
	sram_mem[118918] = 16'b0000000000000000;
	sram_mem[118919] = 16'b0000000000000000;
	sram_mem[118920] = 16'b0000000000000000;
	sram_mem[118921] = 16'b0000000000000000;
	sram_mem[118922] = 16'b0000000000000000;
	sram_mem[118923] = 16'b0000000000000000;
	sram_mem[118924] = 16'b0000000000000000;
	sram_mem[118925] = 16'b0000000000000000;
	sram_mem[118926] = 16'b0000000000000000;
	sram_mem[118927] = 16'b0000000000000000;
	sram_mem[118928] = 16'b0000000000000000;
	sram_mem[118929] = 16'b0000000000000000;
	sram_mem[118930] = 16'b0000000000000000;
	sram_mem[118931] = 16'b0000000000000000;
	sram_mem[118932] = 16'b0000000000000000;
	sram_mem[118933] = 16'b0000000000000000;
	sram_mem[118934] = 16'b0000000000000000;
	sram_mem[118935] = 16'b0000000000000000;
	sram_mem[118936] = 16'b0000000000000000;
	sram_mem[118937] = 16'b0000000000000000;
	sram_mem[118938] = 16'b0000000000000000;
	sram_mem[118939] = 16'b0000000000000000;
	sram_mem[118940] = 16'b0000000000000000;
	sram_mem[118941] = 16'b0000000000000000;
	sram_mem[118942] = 16'b0000000000000000;
	sram_mem[118943] = 16'b0000000000000000;
	sram_mem[118944] = 16'b0000000000000000;
	sram_mem[118945] = 16'b0000000000000000;
	sram_mem[118946] = 16'b0000000000000000;
	sram_mem[118947] = 16'b0000000000000000;
	sram_mem[118948] = 16'b0000000000000000;
	sram_mem[118949] = 16'b0000000000000000;
	sram_mem[118950] = 16'b0000000000000000;
	sram_mem[118951] = 16'b0000000000000000;
	sram_mem[118952] = 16'b0000000000000000;
	sram_mem[118953] = 16'b0000000000000000;
	sram_mem[118954] = 16'b0000000000000000;
	sram_mem[118955] = 16'b0000000000000000;
	sram_mem[118956] = 16'b0000000000000000;
	sram_mem[118957] = 16'b0000000000000000;
	sram_mem[118958] = 16'b0000000000000000;
	sram_mem[118959] = 16'b0000000000000000;
	sram_mem[118960] = 16'b0000000000000000;
	sram_mem[118961] = 16'b0000000000000000;
	sram_mem[118962] = 16'b0000000000000000;
	sram_mem[118963] = 16'b0000000000000000;
	sram_mem[118964] = 16'b0000000000000000;
	sram_mem[118965] = 16'b0000000000000000;
	sram_mem[118966] = 16'b0000000000000000;
	sram_mem[118967] = 16'b0000000000000000;
	sram_mem[118968] = 16'b0000000000000000;
	sram_mem[118969] = 16'b0000000000000000;
	sram_mem[118970] = 16'b0000000000000000;
	sram_mem[118971] = 16'b0000000000000000;
	sram_mem[118972] = 16'b0000000000000000;
	sram_mem[118973] = 16'b0000000000000000;
	sram_mem[118974] = 16'b0000000000000000;
	sram_mem[118975] = 16'b0000000000000000;
	sram_mem[118976] = 16'b0000000000000000;
	sram_mem[118977] = 16'b0000000000000000;
	sram_mem[118978] = 16'b0000000000000000;
	sram_mem[118979] = 16'b0000000000000000;
	sram_mem[118980] = 16'b0000000000000000;
	sram_mem[118981] = 16'b0000000000000000;
	sram_mem[118982] = 16'b0000000000000000;
	sram_mem[118983] = 16'b0000000000000000;
	sram_mem[118984] = 16'b0000000000000000;
	sram_mem[118985] = 16'b0000000000000000;
	sram_mem[118986] = 16'b0000000000000000;
	sram_mem[118987] = 16'b0000000000000000;
	sram_mem[118988] = 16'b0000000000000000;
	sram_mem[118989] = 16'b0000000000000000;
	sram_mem[118990] = 16'b0000000000000000;
	sram_mem[118991] = 16'b0000000000000000;
	sram_mem[118992] = 16'b0000000000000000;
	sram_mem[118993] = 16'b0000000000000000;
	sram_mem[118994] = 16'b0000000000000000;
	sram_mem[118995] = 16'b0000000000000000;
	sram_mem[118996] = 16'b0000000000000000;
	sram_mem[118997] = 16'b0000000000000000;
	sram_mem[118998] = 16'b0000000000000000;
	sram_mem[118999] = 16'b0000000000000000;
	sram_mem[119000] = 16'b0000000000000000;
	sram_mem[119001] = 16'b0000000000000000;
	sram_mem[119002] = 16'b0000000000000000;
	sram_mem[119003] = 16'b0000000000000000;
	sram_mem[119004] = 16'b0000000000000000;
	sram_mem[119005] = 16'b0000000000000000;
	sram_mem[119006] = 16'b0000000000000000;
	sram_mem[119007] = 16'b0000000000000000;
	sram_mem[119008] = 16'b0000000000000000;
	sram_mem[119009] = 16'b0000000000000000;
	sram_mem[119010] = 16'b0000000000000000;
	sram_mem[119011] = 16'b0000000000000000;
	sram_mem[119012] = 16'b0000000000000000;
	sram_mem[119013] = 16'b0000000000000000;
	sram_mem[119014] = 16'b0000000000000000;
	sram_mem[119015] = 16'b0000000000000000;
	sram_mem[119016] = 16'b0000000000000000;
	sram_mem[119017] = 16'b0000000000000000;
	sram_mem[119018] = 16'b0000000000000000;
	sram_mem[119019] = 16'b0000000000000000;
	sram_mem[119020] = 16'b0000000000000000;
	sram_mem[119021] = 16'b0000000000000000;
	sram_mem[119022] = 16'b0000000000000000;
	sram_mem[119023] = 16'b0000000000000000;
	sram_mem[119024] = 16'b0000000000000000;
	sram_mem[119025] = 16'b0000000000000000;
	sram_mem[119026] = 16'b0000000000000000;
	sram_mem[119027] = 16'b0000000000000000;
	sram_mem[119028] = 16'b0000000000000000;
	sram_mem[119029] = 16'b0000000000000000;
	sram_mem[119030] = 16'b0000000000000000;
	sram_mem[119031] = 16'b0000000000000000;
	sram_mem[119032] = 16'b0000000000000000;
	sram_mem[119033] = 16'b0000000000000000;
	sram_mem[119034] = 16'b0000000000000000;
	sram_mem[119035] = 16'b0000000000000000;
	sram_mem[119036] = 16'b0000000000000000;
	sram_mem[119037] = 16'b0000000000000000;
	sram_mem[119038] = 16'b0000000000000000;
	sram_mem[119039] = 16'b0000000000000000;
	sram_mem[119040] = 16'b0000000000000000;
	sram_mem[119041] = 16'b0000000000000000;
	sram_mem[119042] = 16'b0000000000000000;
	sram_mem[119043] = 16'b0000000000000000;
	sram_mem[119044] = 16'b0000000000000000;
	sram_mem[119045] = 16'b0000000000000000;
	sram_mem[119046] = 16'b0000000000000000;
	sram_mem[119047] = 16'b0000000000000000;
	sram_mem[119048] = 16'b0000000000000000;
	sram_mem[119049] = 16'b0000000000000000;
	sram_mem[119050] = 16'b0000000000000000;
	sram_mem[119051] = 16'b0000000000000000;
	sram_mem[119052] = 16'b0000000000000000;
	sram_mem[119053] = 16'b0000000000000000;
	sram_mem[119054] = 16'b0000000000000000;
	sram_mem[119055] = 16'b0000000000000000;
	sram_mem[119056] = 16'b0000000000000000;
	sram_mem[119057] = 16'b0000000000000000;
	sram_mem[119058] = 16'b0000000000000000;
	sram_mem[119059] = 16'b0000000000000000;
	sram_mem[119060] = 16'b0000000000000000;
	sram_mem[119061] = 16'b0000000000000000;
	sram_mem[119062] = 16'b0000000000000000;
	sram_mem[119063] = 16'b0000000000000000;
	sram_mem[119064] = 16'b0000000000000000;
	sram_mem[119065] = 16'b0000000000000000;
	sram_mem[119066] = 16'b0000000000000000;
	sram_mem[119067] = 16'b0000000000000000;
	sram_mem[119068] = 16'b0000000000000000;
	sram_mem[119069] = 16'b0000000000000000;
	sram_mem[119070] = 16'b0000000000000000;
	sram_mem[119071] = 16'b0000000000000000;
	sram_mem[119072] = 16'b0000000000000000;
	sram_mem[119073] = 16'b0000000000000000;
	sram_mem[119074] = 16'b0000000000000000;
	sram_mem[119075] = 16'b0000000000000000;
	sram_mem[119076] = 16'b0000000000000000;
	sram_mem[119077] = 16'b0000000000000000;
	sram_mem[119078] = 16'b0000000000000000;
	sram_mem[119079] = 16'b0000000000000000;
	sram_mem[119080] = 16'b0000000000000000;
	sram_mem[119081] = 16'b0000000000000000;
	sram_mem[119082] = 16'b0000000000000000;
	sram_mem[119083] = 16'b0000000000000000;
	sram_mem[119084] = 16'b0000000000000000;
	sram_mem[119085] = 16'b0000000000000000;
	sram_mem[119086] = 16'b0000000000000000;
	sram_mem[119087] = 16'b0000000000000000;
	sram_mem[119088] = 16'b0000000000000000;
	sram_mem[119089] = 16'b0000000000000000;
	sram_mem[119090] = 16'b0000000000000000;
	sram_mem[119091] = 16'b0000000000000000;
	sram_mem[119092] = 16'b0000000000000000;
	sram_mem[119093] = 16'b0000000000000000;
	sram_mem[119094] = 16'b0000000000000000;
	sram_mem[119095] = 16'b0000000000000000;
	sram_mem[119096] = 16'b0000000000000000;
	sram_mem[119097] = 16'b0000000000000000;
	sram_mem[119098] = 16'b0000000000000000;
	sram_mem[119099] = 16'b0000000000000000;
	sram_mem[119100] = 16'b0000000000000000;
	sram_mem[119101] = 16'b0000000000000000;
	sram_mem[119102] = 16'b0000000000000000;
	sram_mem[119103] = 16'b0000000000000000;
	sram_mem[119104] = 16'b0000000000000000;
	sram_mem[119105] = 16'b0000000000000000;
	sram_mem[119106] = 16'b0000000000000000;
	sram_mem[119107] = 16'b0000000000000000;
	sram_mem[119108] = 16'b0000000000000000;
	sram_mem[119109] = 16'b0000000000000000;
	sram_mem[119110] = 16'b0000000000000000;
	sram_mem[119111] = 16'b0000000000000000;
	sram_mem[119112] = 16'b0000000000000000;
	sram_mem[119113] = 16'b0000000000000000;
	sram_mem[119114] = 16'b0000000000000000;
	sram_mem[119115] = 16'b0000000000000000;
	sram_mem[119116] = 16'b0000000000000000;
	sram_mem[119117] = 16'b0000000000000000;
	sram_mem[119118] = 16'b0000000000000000;
	sram_mem[119119] = 16'b0000000000000000;
	sram_mem[119120] = 16'b0000000000000000;
	sram_mem[119121] = 16'b0000000000000000;
	sram_mem[119122] = 16'b0000000000000000;
	sram_mem[119123] = 16'b0000000000000000;
	sram_mem[119124] = 16'b0000000000000000;
	sram_mem[119125] = 16'b0000000000000000;
	sram_mem[119126] = 16'b0000000000000000;
	sram_mem[119127] = 16'b0000000000000000;
	sram_mem[119128] = 16'b0000000000000000;
	sram_mem[119129] = 16'b0000000000000000;
	sram_mem[119130] = 16'b0000000000000000;
	sram_mem[119131] = 16'b0000000000000000;
	sram_mem[119132] = 16'b0000000000000000;
	sram_mem[119133] = 16'b0000000000000000;
	sram_mem[119134] = 16'b0000000000000000;
	sram_mem[119135] = 16'b0000000000000000;
	sram_mem[119136] = 16'b0000000000000000;
	sram_mem[119137] = 16'b0000000000000000;
	sram_mem[119138] = 16'b0000000000000000;
	sram_mem[119139] = 16'b0000000000000000;
	sram_mem[119140] = 16'b0000000000000000;
	sram_mem[119141] = 16'b0000000000000000;
	sram_mem[119142] = 16'b0000000000000000;
	sram_mem[119143] = 16'b0000000000000000;
	sram_mem[119144] = 16'b0000000000000000;
	sram_mem[119145] = 16'b0000000000000000;
	sram_mem[119146] = 16'b0000000000000000;
	sram_mem[119147] = 16'b0000000000000000;
	sram_mem[119148] = 16'b0000000000000000;
	sram_mem[119149] = 16'b0000000000000000;
	sram_mem[119150] = 16'b0000000000000000;
	sram_mem[119151] = 16'b0000000000000000;
	sram_mem[119152] = 16'b0000000000000000;
	sram_mem[119153] = 16'b0000000000000000;
	sram_mem[119154] = 16'b0000000000000000;
	sram_mem[119155] = 16'b0000000000000000;
	sram_mem[119156] = 16'b0000000000000000;
	sram_mem[119157] = 16'b0000000000000000;
	sram_mem[119158] = 16'b0000000000000000;
	sram_mem[119159] = 16'b0000000000000000;
	sram_mem[119160] = 16'b0000000000000000;
	sram_mem[119161] = 16'b0000000000000000;
	sram_mem[119162] = 16'b0000000000000000;
	sram_mem[119163] = 16'b0000000000000000;
	sram_mem[119164] = 16'b0000000000000000;
	sram_mem[119165] = 16'b0000000000000000;
	sram_mem[119166] = 16'b0000000000000000;
	sram_mem[119167] = 16'b0000000000000000;
	sram_mem[119168] = 16'b0000000000000000;
	sram_mem[119169] = 16'b0000000000000000;
	sram_mem[119170] = 16'b0000000000000000;
	sram_mem[119171] = 16'b0000000000000000;
	sram_mem[119172] = 16'b0000000000000000;
	sram_mem[119173] = 16'b0000000000000000;
	sram_mem[119174] = 16'b0000000000000000;
	sram_mem[119175] = 16'b0000000000000000;
	sram_mem[119176] = 16'b0000000000000000;
	sram_mem[119177] = 16'b0000000000000000;
	sram_mem[119178] = 16'b0000000000000000;
	sram_mem[119179] = 16'b0000000000000000;
	sram_mem[119180] = 16'b0000000000000000;
	sram_mem[119181] = 16'b0000000000000000;
	sram_mem[119182] = 16'b0000000000000000;
	sram_mem[119183] = 16'b0000000000000000;
	sram_mem[119184] = 16'b0000000000000000;
	sram_mem[119185] = 16'b0000000000000000;
	sram_mem[119186] = 16'b0000000000000000;
	sram_mem[119187] = 16'b0000000000000000;
	sram_mem[119188] = 16'b0000000000000000;
	sram_mem[119189] = 16'b0000000000000000;
	sram_mem[119190] = 16'b0000000000000000;
	sram_mem[119191] = 16'b0000000000000000;
	sram_mem[119192] = 16'b0000000000000000;
	sram_mem[119193] = 16'b0000000000000000;
	sram_mem[119194] = 16'b0000000000000000;
	sram_mem[119195] = 16'b0000000000000000;
	sram_mem[119196] = 16'b0000000000000000;
	sram_mem[119197] = 16'b0000000000000000;
	sram_mem[119198] = 16'b0000000000000000;
	sram_mem[119199] = 16'b0000000000000000;
	sram_mem[119200] = 16'b0000000000000000;
	sram_mem[119201] = 16'b0000000000000000;
	sram_mem[119202] = 16'b0000000000000000;
	sram_mem[119203] = 16'b0000000000000000;
	sram_mem[119204] = 16'b0000000000000000;
	sram_mem[119205] = 16'b0000000000000000;
	sram_mem[119206] = 16'b0000000000000000;
	sram_mem[119207] = 16'b0000000000000000;
	sram_mem[119208] = 16'b0000000000000000;
	sram_mem[119209] = 16'b0000000000000000;
	sram_mem[119210] = 16'b0000000000000000;
	sram_mem[119211] = 16'b0000000000000000;
	sram_mem[119212] = 16'b0000000000000000;
	sram_mem[119213] = 16'b0000000000000000;
	sram_mem[119214] = 16'b0000000000000000;
	sram_mem[119215] = 16'b0000000000000000;
	sram_mem[119216] = 16'b0000000000000000;
	sram_mem[119217] = 16'b0000000000000000;
	sram_mem[119218] = 16'b0000000000000000;
	sram_mem[119219] = 16'b0000000000000000;
	sram_mem[119220] = 16'b0000000000000000;
	sram_mem[119221] = 16'b0000000000000000;
	sram_mem[119222] = 16'b0000000000000000;
	sram_mem[119223] = 16'b0000000000000000;
	sram_mem[119224] = 16'b0000000000000000;
	sram_mem[119225] = 16'b0000000000000000;
	sram_mem[119226] = 16'b0000000000000000;
	sram_mem[119227] = 16'b0000000000000000;
	sram_mem[119228] = 16'b0000000000000000;
	sram_mem[119229] = 16'b0000000000000000;
	sram_mem[119230] = 16'b0000000000000000;
	sram_mem[119231] = 16'b0000000000000000;
	sram_mem[119232] = 16'b0000000000000000;
	sram_mem[119233] = 16'b0000000000000000;
	sram_mem[119234] = 16'b0000000000000000;
	sram_mem[119235] = 16'b0000000000000000;
	sram_mem[119236] = 16'b0000000000000000;
	sram_mem[119237] = 16'b0000000000000000;
	sram_mem[119238] = 16'b0000000000000000;
	sram_mem[119239] = 16'b0000000000000000;
	sram_mem[119240] = 16'b0000000000000000;
	sram_mem[119241] = 16'b0000000000000000;
	sram_mem[119242] = 16'b0000000000000000;
	sram_mem[119243] = 16'b0000000000000000;
	sram_mem[119244] = 16'b0000000000000000;
	sram_mem[119245] = 16'b0000000000000000;
	sram_mem[119246] = 16'b0000000000000000;
	sram_mem[119247] = 16'b0000000000000000;
	sram_mem[119248] = 16'b0000000000000000;
	sram_mem[119249] = 16'b0000000000000000;
	sram_mem[119250] = 16'b0000000000000000;
	sram_mem[119251] = 16'b0000000000000000;
	sram_mem[119252] = 16'b0000000000000000;
	sram_mem[119253] = 16'b0000000000000000;
	sram_mem[119254] = 16'b0000000000000000;
	sram_mem[119255] = 16'b0000000000000000;
	sram_mem[119256] = 16'b0000000000000000;
	sram_mem[119257] = 16'b0000000000000000;
	sram_mem[119258] = 16'b0000000000000000;
	sram_mem[119259] = 16'b0000000000000000;
	sram_mem[119260] = 16'b0000000000000000;
	sram_mem[119261] = 16'b0000000000000000;
	sram_mem[119262] = 16'b0000000000000000;
	sram_mem[119263] = 16'b0000000000000000;
	sram_mem[119264] = 16'b0000000000000000;
	sram_mem[119265] = 16'b0000000000000000;
	sram_mem[119266] = 16'b0000000000000000;
	sram_mem[119267] = 16'b0000000000000000;
	sram_mem[119268] = 16'b0000000000000000;
	sram_mem[119269] = 16'b0000000000000000;
	sram_mem[119270] = 16'b0000000000000000;
	sram_mem[119271] = 16'b0000000000000000;
	sram_mem[119272] = 16'b0000000000000000;
	sram_mem[119273] = 16'b0000000000000000;
	sram_mem[119274] = 16'b0000000000000000;
	sram_mem[119275] = 16'b0000000000000000;
	sram_mem[119276] = 16'b0000000000000000;
	sram_mem[119277] = 16'b0000000000000000;
	sram_mem[119278] = 16'b0000000000000000;
	sram_mem[119279] = 16'b0000000000000000;
	sram_mem[119280] = 16'b0000000000000000;
	sram_mem[119281] = 16'b0000000000000000;
	sram_mem[119282] = 16'b0000000000000000;
	sram_mem[119283] = 16'b0000000000000000;
	sram_mem[119284] = 16'b0000000000000000;
	sram_mem[119285] = 16'b0000000000000000;
	sram_mem[119286] = 16'b0000000000000000;
	sram_mem[119287] = 16'b0000000000000000;
	sram_mem[119288] = 16'b0000000000000000;
	sram_mem[119289] = 16'b0000000000000000;
	sram_mem[119290] = 16'b0000000000000000;
	sram_mem[119291] = 16'b0000000000000000;
	sram_mem[119292] = 16'b0000000000000000;
	sram_mem[119293] = 16'b0000000000000000;
	sram_mem[119294] = 16'b0000000000000000;
	sram_mem[119295] = 16'b0000000000000000;
	sram_mem[119296] = 16'b0000000000000000;
	sram_mem[119297] = 16'b0000000000000000;
	sram_mem[119298] = 16'b0000000000000000;
	sram_mem[119299] = 16'b0000000000000000;
	sram_mem[119300] = 16'b0000000000000000;
	sram_mem[119301] = 16'b0000000000000000;
	sram_mem[119302] = 16'b0000000000000000;
	sram_mem[119303] = 16'b0000000000000000;
	sram_mem[119304] = 16'b0000000000000000;
	sram_mem[119305] = 16'b0000000000000000;
	sram_mem[119306] = 16'b0000000000000000;
	sram_mem[119307] = 16'b0000000000000000;
	sram_mem[119308] = 16'b0000000000000000;
	sram_mem[119309] = 16'b0000000000000000;
	sram_mem[119310] = 16'b0000000000000000;
	sram_mem[119311] = 16'b0000000000000000;
	sram_mem[119312] = 16'b0000000000000000;
	sram_mem[119313] = 16'b0000000000000000;
	sram_mem[119314] = 16'b0000000000000000;
	sram_mem[119315] = 16'b0000000000000000;
	sram_mem[119316] = 16'b0000000000000000;
	sram_mem[119317] = 16'b0000000000000000;
	sram_mem[119318] = 16'b0000000000000000;
	sram_mem[119319] = 16'b0000000000000000;
	sram_mem[119320] = 16'b0000000000000000;
	sram_mem[119321] = 16'b0000000000000000;
	sram_mem[119322] = 16'b0000000000000000;
	sram_mem[119323] = 16'b0000000000000000;
	sram_mem[119324] = 16'b0000000000000000;
	sram_mem[119325] = 16'b0000000000000000;
	sram_mem[119326] = 16'b0000000000000000;
	sram_mem[119327] = 16'b0000000000000000;
	sram_mem[119328] = 16'b0000000000000000;
	sram_mem[119329] = 16'b0000000000000000;
	sram_mem[119330] = 16'b0000000000000000;
	sram_mem[119331] = 16'b0000000000000000;
	sram_mem[119332] = 16'b0000000000000000;
	sram_mem[119333] = 16'b0000000000000000;
	sram_mem[119334] = 16'b0000000000000000;
	sram_mem[119335] = 16'b0000000000000000;
	sram_mem[119336] = 16'b0000000000000000;
	sram_mem[119337] = 16'b0000000000000000;
	sram_mem[119338] = 16'b0000000000000000;
	sram_mem[119339] = 16'b0000000000000000;
	sram_mem[119340] = 16'b0000000000000000;
	sram_mem[119341] = 16'b0000000000000000;
	sram_mem[119342] = 16'b0000000000000000;
	sram_mem[119343] = 16'b0000000000000000;
	sram_mem[119344] = 16'b0000000000000000;
	sram_mem[119345] = 16'b0000000000000000;
	sram_mem[119346] = 16'b0000000000000000;
	sram_mem[119347] = 16'b0000000000000000;
	sram_mem[119348] = 16'b0000000000000000;
	sram_mem[119349] = 16'b0000000000000000;
	sram_mem[119350] = 16'b0000000000000000;
	sram_mem[119351] = 16'b0000000000000000;
	sram_mem[119352] = 16'b0000000000000000;
	sram_mem[119353] = 16'b0000000000000000;
	sram_mem[119354] = 16'b0000000000000000;
	sram_mem[119355] = 16'b0000000000000000;
	sram_mem[119356] = 16'b0000000000000000;
	sram_mem[119357] = 16'b0000000000000000;
	sram_mem[119358] = 16'b0000000000000000;
	sram_mem[119359] = 16'b0000000000000000;
	sram_mem[119360] = 16'b0000000000000000;
	sram_mem[119361] = 16'b0000000000000000;
	sram_mem[119362] = 16'b0000000000000000;
	sram_mem[119363] = 16'b0000000000000000;
	sram_mem[119364] = 16'b0000000000000000;
	sram_mem[119365] = 16'b0000000000000000;
	sram_mem[119366] = 16'b0000000000000000;
	sram_mem[119367] = 16'b0000000000000000;
	sram_mem[119368] = 16'b0000000000000000;
	sram_mem[119369] = 16'b0000000000000000;
	sram_mem[119370] = 16'b0000000000000000;
	sram_mem[119371] = 16'b0000000000000000;
	sram_mem[119372] = 16'b0000000000000000;
	sram_mem[119373] = 16'b0000000000000000;
	sram_mem[119374] = 16'b0000000000000000;
	sram_mem[119375] = 16'b0000000000000000;
	sram_mem[119376] = 16'b0000000000000000;
	sram_mem[119377] = 16'b0000000000000000;
	sram_mem[119378] = 16'b0000000000000000;
	sram_mem[119379] = 16'b0000000000000000;
	sram_mem[119380] = 16'b0000000000000000;
	sram_mem[119381] = 16'b0000000000000000;
	sram_mem[119382] = 16'b0000000000000000;
	sram_mem[119383] = 16'b0000000000000000;
	sram_mem[119384] = 16'b0000000000000000;
	sram_mem[119385] = 16'b0000000000000000;
	sram_mem[119386] = 16'b0000000000000000;
	sram_mem[119387] = 16'b0000000000000000;
	sram_mem[119388] = 16'b0000000000000000;
	sram_mem[119389] = 16'b0000000000000000;
	sram_mem[119390] = 16'b0000000000000000;
	sram_mem[119391] = 16'b0000000000000000;
	sram_mem[119392] = 16'b0000000000000000;
	sram_mem[119393] = 16'b0000000000000000;
	sram_mem[119394] = 16'b0000000000000000;
	sram_mem[119395] = 16'b0000000000000000;
	sram_mem[119396] = 16'b0000000000000000;
	sram_mem[119397] = 16'b0000000000000000;
	sram_mem[119398] = 16'b0000000000000000;
	sram_mem[119399] = 16'b0000000000000000;
	sram_mem[119400] = 16'b0000000000000000;
	sram_mem[119401] = 16'b0000000000000000;
	sram_mem[119402] = 16'b0000000000000000;
	sram_mem[119403] = 16'b0000000000000000;
	sram_mem[119404] = 16'b0000000000000000;
	sram_mem[119405] = 16'b0000000000000000;
	sram_mem[119406] = 16'b0000000000000000;
	sram_mem[119407] = 16'b0000000000000000;
	sram_mem[119408] = 16'b0000000000000000;
	sram_mem[119409] = 16'b0000000000000000;
	sram_mem[119410] = 16'b0000000000000000;
	sram_mem[119411] = 16'b0000000000000000;
	sram_mem[119412] = 16'b0000000000000000;
	sram_mem[119413] = 16'b0000000000000000;
	sram_mem[119414] = 16'b0000000000000000;
	sram_mem[119415] = 16'b0000000000000000;
	sram_mem[119416] = 16'b0000000000000000;
	sram_mem[119417] = 16'b0000000000000000;
	sram_mem[119418] = 16'b0000000000000000;
	sram_mem[119419] = 16'b0000000000000000;
	sram_mem[119420] = 16'b0000000000000000;
	sram_mem[119421] = 16'b0000000000000000;
	sram_mem[119422] = 16'b0000000000000000;
	sram_mem[119423] = 16'b0000000000000000;
	sram_mem[119424] = 16'b0000000000000000;
	sram_mem[119425] = 16'b0000000000000000;
	sram_mem[119426] = 16'b0000000000000000;
	sram_mem[119427] = 16'b0000000000000000;
	sram_mem[119428] = 16'b0000000000000000;
	sram_mem[119429] = 16'b0000000000000000;
	sram_mem[119430] = 16'b0000000000000000;
	sram_mem[119431] = 16'b0000000000000000;
	sram_mem[119432] = 16'b0000000000000000;
	sram_mem[119433] = 16'b0000000000000000;
	sram_mem[119434] = 16'b0000000000000000;
	sram_mem[119435] = 16'b0000000000000000;
	sram_mem[119436] = 16'b0000000000000000;
	sram_mem[119437] = 16'b0000000000000000;
	sram_mem[119438] = 16'b0000000000000000;
	sram_mem[119439] = 16'b0000000000000000;
	sram_mem[119440] = 16'b0000000000000000;
	sram_mem[119441] = 16'b0000000000000000;
	sram_mem[119442] = 16'b0000000000000000;
	sram_mem[119443] = 16'b0000000000000000;
	sram_mem[119444] = 16'b0000000000000000;
	sram_mem[119445] = 16'b0000000000000000;
	sram_mem[119446] = 16'b0000000000000000;
	sram_mem[119447] = 16'b0000000000000000;
	sram_mem[119448] = 16'b0000000000000000;
	sram_mem[119449] = 16'b0000000000000000;
	sram_mem[119450] = 16'b0000000000000000;
	sram_mem[119451] = 16'b0000000000000000;
	sram_mem[119452] = 16'b0000000000000000;
	sram_mem[119453] = 16'b0000000000000000;
	sram_mem[119454] = 16'b0000000000000000;
	sram_mem[119455] = 16'b0000000000000000;
	sram_mem[119456] = 16'b0000000000000000;
	sram_mem[119457] = 16'b0000000000000000;
	sram_mem[119458] = 16'b0000000000000000;
	sram_mem[119459] = 16'b0000000000000000;
	sram_mem[119460] = 16'b0000000000000000;
	sram_mem[119461] = 16'b0000000000000000;
	sram_mem[119462] = 16'b0000000000000000;
	sram_mem[119463] = 16'b0000000000000000;
	sram_mem[119464] = 16'b0000000000000000;
	sram_mem[119465] = 16'b0000000000000000;
	sram_mem[119466] = 16'b0000000000000000;
	sram_mem[119467] = 16'b0000000000000000;
	sram_mem[119468] = 16'b0000000000000000;
	sram_mem[119469] = 16'b0000000000000000;
	sram_mem[119470] = 16'b0000000000000000;
	sram_mem[119471] = 16'b0000000000000000;
	sram_mem[119472] = 16'b0000000000000000;
	sram_mem[119473] = 16'b0000000000000000;
	sram_mem[119474] = 16'b0000000000000000;
	sram_mem[119475] = 16'b0000000000000000;
	sram_mem[119476] = 16'b0000000000000000;
	sram_mem[119477] = 16'b0000000000000000;
	sram_mem[119478] = 16'b0000000000000000;
	sram_mem[119479] = 16'b0000000000000000;
	sram_mem[119480] = 16'b0000000000000000;
	sram_mem[119481] = 16'b0000000000000000;
	sram_mem[119482] = 16'b0000000000000000;
	sram_mem[119483] = 16'b0000000000000000;
	sram_mem[119484] = 16'b0000000000000000;
	sram_mem[119485] = 16'b0000000000000000;
	sram_mem[119486] = 16'b0000000000000000;
	sram_mem[119487] = 16'b0000000000000000;
	sram_mem[119488] = 16'b0000000000000000;
	sram_mem[119489] = 16'b0000000000000000;
	sram_mem[119490] = 16'b0000000000000000;
	sram_mem[119491] = 16'b0000000000000000;
	sram_mem[119492] = 16'b0000000000000000;
	sram_mem[119493] = 16'b0000000000000000;
	sram_mem[119494] = 16'b0000000000000000;
	sram_mem[119495] = 16'b0000000000000000;
	sram_mem[119496] = 16'b0000000000000000;
	sram_mem[119497] = 16'b0000000000000000;
	sram_mem[119498] = 16'b0000000000000000;
	sram_mem[119499] = 16'b0000000000000000;
	sram_mem[119500] = 16'b0000000000000000;
	sram_mem[119501] = 16'b0000000000000000;
	sram_mem[119502] = 16'b0000000000000000;
	sram_mem[119503] = 16'b0000000000000000;
	sram_mem[119504] = 16'b0000000000000000;
	sram_mem[119505] = 16'b0000000000000000;
	sram_mem[119506] = 16'b0000000000000000;
	sram_mem[119507] = 16'b0000000000000000;
	sram_mem[119508] = 16'b0000000000000000;
	sram_mem[119509] = 16'b0000000000000000;
	sram_mem[119510] = 16'b0000000000000000;
	sram_mem[119511] = 16'b0000000000000000;
	sram_mem[119512] = 16'b0000000000000000;
	sram_mem[119513] = 16'b0000000000000000;
	sram_mem[119514] = 16'b0000000000000000;
	sram_mem[119515] = 16'b0000000000000000;
	sram_mem[119516] = 16'b0000000000000000;
	sram_mem[119517] = 16'b0000000000000000;
	sram_mem[119518] = 16'b0000000000000000;
	sram_mem[119519] = 16'b0000000000000000;
	sram_mem[119520] = 16'b0000000000000000;
	sram_mem[119521] = 16'b0000000000000000;
	sram_mem[119522] = 16'b0000000000000000;
	sram_mem[119523] = 16'b0000000000000000;
	sram_mem[119524] = 16'b0000000000000000;
	sram_mem[119525] = 16'b0000000000000000;
	sram_mem[119526] = 16'b0000000000000000;
	sram_mem[119527] = 16'b0000000000000000;
	sram_mem[119528] = 16'b0000000000000000;
	sram_mem[119529] = 16'b0000000000000000;
	sram_mem[119530] = 16'b0000000000000000;
	sram_mem[119531] = 16'b0000000000000000;
	sram_mem[119532] = 16'b0000000000000000;
	sram_mem[119533] = 16'b0000000000000000;
	sram_mem[119534] = 16'b0000000000000000;
	sram_mem[119535] = 16'b0000000000000000;
	sram_mem[119536] = 16'b0000000000000000;
	sram_mem[119537] = 16'b0000000000000000;
	sram_mem[119538] = 16'b0000000000000000;
	sram_mem[119539] = 16'b0000000000000000;
	sram_mem[119540] = 16'b0000000000000000;
	sram_mem[119541] = 16'b0000000000000000;
	sram_mem[119542] = 16'b0000000000000000;
	sram_mem[119543] = 16'b0000000000000000;
	sram_mem[119544] = 16'b0000000000000000;
	sram_mem[119545] = 16'b0000000000000000;
	sram_mem[119546] = 16'b0000000000000000;
	sram_mem[119547] = 16'b0000000000000000;
	sram_mem[119548] = 16'b0000000000000000;
	sram_mem[119549] = 16'b0000000000000000;
	sram_mem[119550] = 16'b0000000000000000;
	sram_mem[119551] = 16'b0000000000000000;
	sram_mem[119552] = 16'b0000000000000000;
	sram_mem[119553] = 16'b0000000000000000;
	sram_mem[119554] = 16'b0000000000000000;
	sram_mem[119555] = 16'b0000000000000000;
	sram_mem[119556] = 16'b0000000000000000;
	sram_mem[119557] = 16'b0000000000000000;
	sram_mem[119558] = 16'b0000000000000000;
	sram_mem[119559] = 16'b0000000000000000;
	sram_mem[119560] = 16'b0000000000000000;
	sram_mem[119561] = 16'b0000000000000000;
	sram_mem[119562] = 16'b0000000000000000;
	sram_mem[119563] = 16'b0000000000000000;
	sram_mem[119564] = 16'b0000000000000000;
	sram_mem[119565] = 16'b0000000000000000;
	sram_mem[119566] = 16'b0000000000000000;
	sram_mem[119567] = 16'b0000000000000000;
	sram_mem[119568] = 16'b0000000000000000;
	sram_mem[119569] = 16'b0000000000000000;
	sram_mem[119570] = 16'b0000000000000000;
	sram_mem[119571] = 16'b0000000000000000;
	sram_mem[119572] = 16'b0000000000000000;
	sram_mem[119573] = 16'b0000000000000000;
	sram_mem[119574] = 16'b0000000000000000;
	sram_mem[119575] = 16'b0000000000000000;
	sram_mem[119576] = 16'b0000000000000000;
	sram_mem[119577] = 16'b0000000000000000;
	sram_mem[119578] = 16'b0000000000000000;
	sram_mem[119579] = 16'b0000000000000000;
	sram_mem[119580] = 16'b0000000000000000;
	sram_mem[119581] = 16'b0000000000000000;
	sram_mem[119582] = 16'b0000000000000000;
	sram_mem[119583] = 16'b0000000000000000;
	sram_mem[119584] = 16'b0000000000000000;
	sram_mem[119585] = 16'b0000000000000000;
	sram_mem[119586] = 16'b0000000000000000;
	sram_mem[119587] = 16'b0000000000000000;
	sram_mem[119588] = 16'b0000000000000000;
	sram_mem[119589] = 16'b0000000000000000;
	sram_mem[119590] = 16'b0000000000000000;
	sram_mem[119591] = 16'b0000000000000000;
	sram_mem[119592] = 16'b0000000000000000;
	sram_mem[119593] = 16'b0000000000000000;
	sram_mem[119594] = 16'b0000000000000000;
	sram_mem[119595] = 16'b0000000000000000;
	sram_mem[119596] = 16'b0000000000000000;
	sram_mem[119597] = 16'b0000000000000000;
	sram_mem[119598] = 16'b0000000000000000;
	sram_mem[119599] = 16'b0000000000000000;
	sram_mem[119600] = 16'b0000000000000000;
	sram_mem[119601] = 16'b0000000000000000;
	sram_mem[119602] = 16'b0000000000000000;
	sram_mem[119603] = 16'b0000000000000000;
	sram_mem[119604] = 16'b0000000000000000;
	sram_mem[119605] = 16'b0000000000000000;
	sram_mem[119606] = 16'b0000000000000000;
	sram_mem[119607] = 16'b0000000000000000;
	sram_mem[119608] = 16'b0000000000000000;
	sram_mem[119609] = 16'b0000000000000000;
	sram_mem[119610] = 16'b0000000000000000;
	sram_mem[119611] = 16'b0000000000000000;
	sram_mem[119612] = 16'b0000000000000000;
	sram_mem[119613] = 16'b0000000000000000;
	sram_mem[119614] = 16'b0000000000000000;
	sram_mem[119615] = 16'b0000000000000000;
	sram_mem[119616] = 16'b0000000000000000;
	sram_mem[119617] = 16'b0000000000000000;
	sram_mem[119618] = 16'b0000000000000000;
	sram_mem[119619] = 16'b0000000000000000;
	sram_mem[119620] = 16'b0000000000000000;
	sram_mem[119621] = 16'b0000000000000000;
	sram_mem[119622] = 16'b0000000000000000;
	sram_mem[119623] = 16'b0000000000000000;
	sram_mem[119624] = 16'b0000000000000000;
	sram_mem[119625] = 16'b0000000000000000;
	sram_mem[119626] = 16'b0000000000000000;
	sram_mem[119627] = 16'b0000000000000000;
	sram_mem[119628] = 16'b0000000000000000;
	sram_mem[119629] = 16'b0000000000000000;
	sram_mem[119630] = 16'b0000000000000000;
	sram_mem[119631] = 16'b0000000000000000;
	sram_mem[119632] = 16'b0000000000000000;
	sram_mem[119633] = 16'b0000000000000000;
	sram_mem[119634] = 16'b0000000000000000;
	sram_mem[119635] = 16'b0000000000000000;
	sram_mem[119636] = 16'b0000000000000000;
	sram_mem[119637] = 16'b0000000000000000;
	sram_mem[119638] = 16'b0000000000000000;
	sram_mem[119639] = 16'b0000000000000000;
	sram_mem[119640] = 16'b0000000000000000;
	sram_mem[119641] = 16'b0000000000000000;
	sram_mem[119642] = 16'b0000000000000000;
	sram_mem[119643] = 16'b0000000000000000;
	sram_mem[119644] = 16'b0000000000000000;
	sram_mem[119645] = 16'b0000000000000000;
	sram_mem[119646] = 16'b0000000000000000;
	sram_mem[119647] = 16'b0000000000000000;
	sram_mem[119648] = 16'b0000000000000000;
	sram_mem[119649] = 16'b0000000000000000;
	sram_mem[119650] = 16'b0000000000000000;
	sram_mem[119651] = 16'b0000000000000000;
	sram_mem[119652] = 16'b0000000000000000;
	sram_mem[119653] = 16'b0000000000000000;
	sram_mem[119654] = 16'b0000000000000000;
	sram_mem[119655] = 16'b0000000000000000;
	sram_mem[119656] = 16'b0000000000000000;
	sram_mem[119657] = 16'b0000000000000000;
	sram_mem[119658] = 16'b0000000000000000;
	sram_mem[119659] = 16'b0000000000000000;
	sram_mem[119660] = 16'b0000000000000000;
	sram_mem[119661] = 16'b0000000000000000;
	sram_mem[119662] = 16'b0000000000000000;
	sram_mem[119663] = 16'b0000000000000000;
	sram_mem[119664] = 16'b0000000000000000;
	sram_mem[119665] = 16'b0000000000000000;
	sram_mem[119666] = 16'b0000000000000000;
	sram_mem[119667] = 16'b0000000000000000;
	sram_mem[119668] = 16'b0000000000000000;
	sram_mem[119669] = 16'b0000000000000000;
	sram_mem[119670] = 16'b0000000000000000;
	sram_mem[119671] = 16'b0000000000000000;
	sram_mem[119672] = 16'b0000000000000000;
	sram_mem[119673] = 16'b0000000000000000;
	sram_mem[119674] = 16'b0000000000000000;
	sram_mem[119675] = 16'b0000000000000000;
	sram_mem[119676] = 16'b0000000000000000;
	sram_mem[119677] = 16'b0000000000000000;
	sram_mem[119678] = 16'b0000000000000000;
	sram_mem[119679] = 16'b0000000000000000;
	sram_mem[119680] = 16'b0000000000000000;
	sram_mem[119681] = 16'b0000000000000000;
	sram_mem[119682] = 16'b0000000000000000;
	sram_mem[119683] = 16'b0000000000000000;
	sram_mem[119684] = 16'b0000000000000000;
	sram_mem[119685] = 16'b0000000000000000;
	sram_mem[119686] = 16'b0000000000000000;
	sram_mem[119687] = 16'b0000000000000000;
	sram_mem[119688] = 16'b0000000000000000;
	sram_mem[119689] = 16'b0000000000000000;
	sram_mem[119690] = 16'b0000000000000000;
	sram_mem[119691] = 16'b0000000000000000;
	sram_mem[119692] = 16'b0000000000000000;
	sram_mem[119693] = 16'b0000000000000000;
	sram_mem[119694] = 16'b0000000000000000;
	sram_mem[119695] = 16'b0000000000000000;
	sram_mem[119696] = 16'b0000000000000000;
	sram_mem[119697] = 16'b0000000000000000;
	sram_mem[119698] = 16'b0000000000000000;
	sram_mem[119699] = 16'b0000000000000000;
	sram_mem[119700] = 16'b0000000000000000;
	sram_mem[119701] = 16'b0000000000000000;
	sram_mem[119702] = 16'b0000000000000000;
	sram_mem[119703] = 16'b0000000000000000;
	sram_mem[119704] = 16'b0000000000000000;
	sram_mem[119705] = 16'b0000000000000000;
	sram_mem[119706] = 16'b0000000000000000;
	sram_mem[119707] = 16'b0000000000000000;
	sram_mem[119708] = 16'b0000000000000000;
	sram_mem[119709] = 16'b0000000000000000;
	sram_mem[119710] = 16'b0000000000000000;
	sram_mem[119711] = 16'b0000000000000000;
	sram_mem[119712] = 16'b0000000000000000;
	sram_mem[119713] = 16'b0000000000000000;
	sram_mem[119714] = 16'b0000000000000000;
	sram_mem[119715] = 16'b0000000000000000;
	sram_mem[119716] = 16'b0000000000000000;
	sram_mem[119717] = 16'b0000000000000000;
	sram_mem[119718] = 16'b0000000000000000;
	sram_mem[119719] = 16'b0000000000000000;
	sram_mem[119720] = 16'b0000000000000000;
	sram_mem[119721] = 16'b0000000000000000;
	sram_mem[119722] = 16'b0000000000000000;
	sram_mem[119723] = 16'b0000000000000000;
	sram_mem[119724] = 16'b0000000000000000;
	sram_mem[119725] = 16'b0000000000000000;
	sram_mem[119726] = 16'b0000000000000000;
	sram_mem[119727] = 16'b0000000000000000;
	sram_mem[119728] = 16'b0000000000000000;
	sram_mem[119729] = 16'b0000000000000000;
	sram_mem[119730] = 16'b0000000000000000;
	sram_mem[119731] = 16'b0000000000000000;
	sram_mem[119732] = 16'b0000000000000000;
	sram_mem[119733] = 16'b0000000000000000;
	sram_mem[119734] = 16'b0000000000000000;
	sram_mem[119735] = 16'b0000000000000000;
	sram_mem[119736] = 16'b0000000000000000;
	sram_mem[119737] = 16'b0000000000000000;
	sram_mem[119738] = 16'b0000000000000000;
	sram_mem[119739] = 16'b0000000000000000;
	sram_mem[119740] = 16'b0000000000000000;
	sram_mem[119741] = 16'b0000000000000000;
	sram_mem[119742] = 16'b0000000000000000;
	sram_mem[119743] = 16'b0000000000000000;
	sram_mem[119744] = 16'b0000000000000000;
	sram_mem[119745] = 16'b0000000000000000;
	sram_mem[119746] = 16'b0000000000000000;
	sram_mem[119747] = 16'b0000000000000000;
	sram_mem[119748] = 16'b0000000000000000;
	sram_mem[119749] = 16'b0000000000000000;
	sram_mem[119750] = 16'b0000000000000000;
	sram_mem[119751] = 16'b0000000000000000;
	sram_mem[119752] = 16'b0000000000000000;
	sram_mem[119753] = 16'b0000000000000000;
	sram_mem[119754] = 16'b0000000000000000;
	sram_mem[119755] = 16'b0000000000000000;
	sram_mem[119756] = 16'b0000000000000000;
	sram_mem[119757] = 16'b0000000000000000;
	sram_mem[119758] = 16'b0000000000000000;
	sram_mem[119759] = 16'b0000000000000000;
	sram_mem[119760] = 16'b0000000000000000;
	sram_mem[119761] = 16'b0000000000000000;
	sram_mem[119762] = 16'b0000000000000000;
	sram_mem[119763] = 16'b0000000000000000;
	sram_mem[119764] = 16'b0000000000000000;
	sram_mem[119765] = 16'b0000000000000000;
	sram_mem[119766] = 16'b0000000000000000;
	sram_mem[119767] = 16'b0000000000000000;
	sram_mem[119768] = 16'b0000000000000000;
	sram_mem[119769] = 16'b0000000000000000;
	sram_mem[119770] = 16'b0000000000000000;
	sram_mem[119771] = 16'b0000000000000000;
	sram_mem[119772] = 16'b0000000000000000;
	sram_mem[119773] = 16'b0000000000000000;
	sram_mem[119774] = 16'b0000000000000000;
	sram_mem[119775] = 16'b0000000000000000;
	sram_mem[119776] = 16'b0000000000000000;
	sram_mem[119777] = 16'b0000000000000000;
	sram_mem[119778] = 16'b0000000000000000;
	sram_mem[119779] = 16'b0000000000000000;
	sram_mem[119780] = 16'b0000000000000000;
	sram_mem[119781] = 16'b0000000000000000;
	sram_mem[119782] = 16'b0000000000000000;
	sram_mem[119783] = 16'b0000000000000000;
	sram_mem[119784] = 16'b0000000000000000;
	sram_mem[119785] = 16'b0000000000000000;
	sram_mem[119786] = 16'b0000000000000000;
	sram_mem[119787] = 16'b0000000000000000;
	sram_mem[119788] = 16'b0000000000000000;
	sram_mem[119789] = 16'b0000000000000000;
	sram_mem[119790] = 16'b0000000000000000;
	sram_mem[119791] = 16'b0000000000000000;
	sram_mem[119792] = 16'b0000000000000000;
	sram_mem[119793] = 16'b0000000000000000;
	sram_mem[119794] = 16'b0000000000000000;
	sram_mem[119795] = 16'b0000000000000000;
	sram_mem[119796] = 16'b0000000000000000;
	sram_mem[119797] = 16'b0000000000000000;
	sram_mem[119798] = 16'b0000000000000000;
	sram_mem[119799] = 16'b0000000000000000;
	sram_mem[119800] = 16'b0000000000000000;
	sram_mem[119801] = 16'b0000000000000000;
	sram_mem[119802] = 16'b0000000000000000;
	sram_mem[119803] = 16'b0000000000000000;
	sram_mem[119804] = 16'b0000000000000000;
	sram_mem[119805] = 16'b0000000000000000;
	sram_mem[119806] = 16'b0000000000000000;
	sram_mem[119807] = 16'b0000000000000000;
	sram_mem[119808] = 16'b0000000000000000;
	sram_mem[119809] = 16'b0000000000000000;
	sram_mem[119810] = 16'b0000000000000000;
	sram_mem[119811] = 16'b0000000000000000;
	sram_mem[119812] = 16'b0000000000000000;
	sram_mem[119813] = 16'b0000000000000000;
	sram_mem[119814] = 16'b0000000000000000;
	sram_mem[119815] = 16'b0000000000000000;
	sram_mem[119816] = 16'b0000000000000000;
	sram_mem[119817] = 16'b0000000000000000;
	sram_mem[119818] = 16'b0000000000000000;
	sram_mem[119819] = 16'b0000000000000000;
	sram_mem[119820] = 16'b0000000000000000;
	sram_mem[119821] = 16'b0000000000000000;
	sram_mem[119822] = 16'b0000000000000000;
	sram_mem[119823] = 16'b0000000000000000;
	sram_mem[119824] = 16'b0000000000000000;
	sram_mem[119825] = 16'b0000000000000000;
	sram_mem[119826] = 16'b0000000000000000;
	sram_mem[119827] = 16'b0000000000000000;
	sram_mem[119828] = 16'b0000000000000000;
	sram_mem[119829] = 16'b0000000000000000;
	sram_mem[119830] = 16'b0000000000000000;
	sram_mem[119831] = 16'b0000000000000000;
	sram_mem[119832] = 16'b0000000000000000;
	sram_mem[119833] = 16'b0000000000000000;
	sram_mem[119834] = 16'b0000000000000000;
	sram_mem[119835] = 16'b0000000000000000;
	sram_mem[119836] = 16'b0000000000000000;
	sram_mem[119837] = 16'b0000000000000000;
	sram_mem[119838] = 16'b0000000000000000;
	sram_mem[119839] = 16'b0000000000000000;
	sram_mem[119840] = 16'b0000000000000000;
	sram_mem[119841] = 16'b0000000000000000;
	sram_mem[119842] = 16'b0000000000000000;
	sram_mem[119843] = 16'b0000000000000000;
	sram_mem[119844] = 16'b0000000000000000;
	sram_mem[119845] = 16'b0000000000000000;
	sram_mem[119846] = 16'b0000000000000000;
	sram_mem[119847] = 16'b0000000000000000;
	sram_mem[119848] = 16'b0000000000000000;
	sram_mem[119849] = 16'b0000000000000000;
	sram_mem[119850] = 16'b0000000000000000;
	sram_mem[119851] = 16'b0000000000000000;
	sram_mem[119852] = 16'b0000000000000000;
	sram_mem[119853] = 16'b0000000000000000;
	sram_mem[119854] = 16'b0000000000000000;
	sram_mem[119855] = 16'b0000000000000000;
	sram_mem[119856] = 16'b0000000000000000;
	sram_mem[119857] = 16'b0000000000000000;
	sram_mem[119858] = 16'b0000000000000000;
	sram_mem[119859] = 16'b0000000000000000;
	sram_mem[119860] = 16'b0000000000000000;
	sram_mem[119861] = 16'b0000000000000000;
	sram_mem[119862] = 16'b0000000000000000;
	sram_mem[119863] = 16'b0000000000000000;
	sram_mem[119864] = 16'b0000000000000000;
	sram_mem[119865] = 16'b0000000000000000;
	sram_mem[119866] = 16'b0000000000000000;
	sram_mem[119867] = 16'b0000000000000000;
	sram_mem[119868] = 16'b0000000000000000;
	sram_mem[119869] = 16'b0000000000000000;
	sram_mem[119870] = 16'b0000000000000000;
	sram_mem[119871] = 16'b0000000000000000;
	sram_mem[119872] = 16'b0000000000000000;
	sram_mem[119873] = 16'b0000000000000000;
	sram_mem[119874] = 16'b0000000000000000;
	sram_mem[119875] = 16'b0000000000000000;
	sram_mem[119876] = 16'b0000000000000000;
	sram_mem[119877] = 16'b0000000000000000;
	sram_mem[119878] = 16'b0000000000000000;
	sram_mem[119879] = 16'b0000000000000000;
	sram_mem[119880] = 16'b0000000000000000;
	sram_mem[119881] = 16'b0000000000000000;
	sram_mem[119882] = 16'b0000000000000000;
	sram_mem[119883] = 16'b0000000000000000;
	sram_mem[119884] = 16'b0000000000000000;
	sram_mem[119885] = 16'b0000000000000000;
	sram_mem[119886] = 16'b0000000000000000;
	sram_mem[119887] = 16'b0000000000000000;
	sram_mem[119888] = 16'b0000000000000000;
	sram_mem[119889] = 16'b0000000000000000;
	sram_mem[119890] = 16'b0000000000000000;
	sram_mem[119891] = 16'b0000000000000000;
	sram_mem[119892] = 16'b0000000000000000;
	sram_mem[119893] = 16'b0000000000000000;
	sram_mem[119894] = 16'b0000000000000000;
	sram_mem[119895] = 16'b0000000000000000;
	sram_mem[119896] = 16'b0000000000000000;
	sram_mem[119897] = 16'b0000000000000000;
	sram_mem[119898] = 16'b0000000000000000;
	sram_mem[119899] = 16'b0000000000000000;
	sram_mem[119900] = 16'b0000000000000000;
	sram_mem[119901] = 16'b0000000000000000;
	sram_mem[119902] = 16'b0000000000000000;
	sram_mem[119903] = 16'b0000000000000000;
	sram_mem[119904] = 16'b0000000000000000;
	sram_mem[119905] = 16'b0000000000000000;
	sram_mem[119906] = 16'b0000000000000000;
	sram_mem[119907] = 16'b0000000000000000;
	sram_mem[119908] = 16'b0000000000000000;
	sram_mem[119909] = 16'b0000000000000000;
	sram_mem[119910] = 16'b0000000000000000;
	sram_mem[119911] = 16'b0000000000000000;
	sram_mem[119912] = 16'b0000000000000000;
	sram_mem[119913] = 16'b0000000000000000;
	sram_mem[119914] = 16'b0000000000000000;
	sram_mem[119915] = 16'b0000000000000000;
	sram_mem[119916] = 16'b0000000000000000;
	sram_mem[119917] = 16'b0000000000000000;
	sram_mem[119918] = 16'b0000000000000000;
	sram_mem[119919] = 16'b0000000000000000;
	sram_mem[119920] = 16'b0000000000000000;
	sram_mem[119921] = 16'b0000000000000000;
	sram_mem[119922] = 16'b0000000000000000;
	sram_mem[119923] = 16'b0000000000000000;
	sram_mem[119924] = 16'b0000000000000000;
	sram_mem[119925] = 16'b0000000000000000;
	sram_mem[119926] = 16'b0000000000000000;
	sram_mem[119927] = 16'b0000000000000000;
	sram_mem[119928] = 16'b0000000000000000;
	sram_mem[119929] = 16'b0000000000000000;
	sram_mem[119930] = 16'b0000000000000000;
	sram_mem[119931] = 16'b0000000000000000;
	sram_mem[119932] = 16'b0000000000000000;
	sram_mem[119933] = 16'b0000000000000000;
	sram_mem[119934] = 16'b0000000000000000;
	sram_mem[119935] = 16'b0000000000000000;
	sram_mem[119936] = 16'b0000000000000000;
	sram_mem[119937] = 16'b0000000000000000;
	sram_mem[119938] = 16'b0000000000000000;
	sram_mem[119939] = 16'b0000000000000000;
	sram_mem[119940] = 16'b0000000000000000;
	sram_mem[119941] = 16'b0000000000000000;
	sram_mem[119942] = 16'b0000000000000000;
	sram_mem[119943] = 16'b0000000000000000;
	sram_mem[119944] = 16'b0000000000000000;
	sram_mem[119945] = 16'b0000000000000000;
	sram_mem[119946] = 16'b0000000000000000;
	sram_mem[119947] = 16'b0000000000000000;
	sram_mem[119948] = 16'b0000000000000000;
	sram_mem[119949] = 16'b0000000000000000;
	sram_mem[119950] = 16'b0000000000000000;
	sram_mem[119951] = 16'b0000000000000000;
	sram_mem[119952] = 16'b0000000000000000;
	sram_mem[119953] = 16'b0000000000000000;
	sram_mem[119954] = 16'b0000000000000000;
	sram_mem[119955] = 16'b0000000000000000;
	sram_mem[119956] = 16'b0000000000000000;
	sram_mem[119957] = 16'b0000000000000000;
	sram_mem[119958] = 16'b0000000000000000;
	sram_mem[119959] = 16'b0000000000000000;
	sram_mem[119960] = 16'b0000000000000000;
	sram_mem[119961] = 16'b0000000000000000;
	sram_mem[119962] = 16'b0000000000000000;
	sram_mem[119963] = 16'b0000000000000000;
	sram_mem[119964] = 16'b0000000000000000;
	sram_mem[119965] = 16'b0000000000000000;
	sram_mem[119966] = 16'b0000000000000000;
	sram_mem[119967] = 16'b0000000000000000;
	sram_mem[119968] = 16'b0000000000000000;
	sram_mem[119969] = 16'b0000000000000000;
	sram_mem[119970] = 16'b0000000000000000;
	sram_mem[119971] = 16'b0000000000000000;
	sram_mem[119972] = 16'b0000000000000000;
	sram_mem[119973] = 16'b0000000000000000;
	sram_mem[119974] = 16'b0000000000000000;
	sram_mem[119975] = 16'b0000000000000000;
	sram_mem[119976] = 16'b0000000000000000;
	sram_mem[119977] = 16'b0000000000000000;
	sram_mem[119978] = 16'b0000000000000000;
	sram_mem[119979] = 16'b0000000000000000;
	sram_mem[119980] = 16'b0000000000000000;
	sram_mem[119981] = 16'b0000000000000000;
	sram_mem[119982] = 16'b0000000000000000;
	sram_mem[119983] = 16'b0000000000000000;
	sram_mem[119984] = 16'b0000000000000000;
	sram_mem[119985] = 16'b0000000000000000;
	sram_mem[119986] = 16'b0000000000000000;
	sram_mem[119987] = 16'b0000000000000000;
	sram_mem[119988] = 16'b0000000000000000;
	sram_mem[119989] = 16'b0000000000000000;
	sram_mem[119990] = 16'b0000000000000000;
	sram_mem[119991] = 16'b0000000000000000;
	sram_mem[119992] = 16'b0000000000000000;
	sram_mem[119993] = 16'b0000000000000000;
	sram_mem[119994] = 16'b0000000000000000;
	sram_mem[119995] = 16'b0000000000000000;
	sram_mem[119996] = 16'b0000000000000000;
	sram_mem[119997] = 16'b0000000000000000;
	sram_mem[119998] = 16'b0000000000000000;
	sram_mem[119999] = 16'b0000000000000000;
	sram_mem[120000] = 16'b0000000000000000;
	sram_mem[120001] = 16'b0000000000000000;
	sram_mem[120002] = 16'b0000000000000000;
	sram_mem[120003] = 16'b0000000000000000;
	sram_mem[120004] = 16'b0000000000000000;
	sram_mem[120005] = 16'b0000000000000000;
	sram_mem[120006] = 16'b0000000000000000;
	sram_mem[120007] = 16'b0000000000000000;
	sram_mem[120008] = 16'b0000000000000000;
	sram_mem[120009] = 16'b0000000000000000;
	sram_mem[120010] = 16'b0000000000000000;
	sram_mem[120011] = 16'b0000000000000000;
	sram_mem[120012] = 16'b0000000000000000;
	sram_mem[120013] = 16'b0000000000000000;
	sram_mem[120014] = 16'b0000000000000000;
	sram_mem[120015] = 16'b0000000000000000;
	sram_mem[120016] = 16'b0000000000000000;
	sram_mem[120017] = 16'b0000000000000000;
	sram_mem[120018] = 16'b0000000000000000;
	sram_mem[120019] = 16'b0000000000000000;
	sram_mem[120020] = 16'b0000000000000000;
	sram_mem[120021] = 16'b0000000000000000;
	sram_mem[120022] = 16'b0000000000000000;
	sram_mem[120023] = 16'b0000000000000000;
	sram_mem[120024] = 16'b0000000000000000;
	sram_mem[120025] = 16'b0000000000000000;
	sram_mem[120026] = 16'b0000000000000000;
	sram_mem[120027] = 16'b0000000000000000;
	sram_mem[120028] = 16'b0000000000000000;
	sram_mem[120029] = 16'b0000000000000000;
	sram_mem[120030] = 16'b0000000000000000;
	sram_mem[120031] = 16'b0000000000000000;
	sram_mem[120032] = 16'b0000000000000000;
	sram_mem[120033] = 16'b0000000000000000;
	sram_mem[120034] = 16'b0000000000000000;
	sram_mem[120035] = 16'b0000000000000000;
	sram_mem[120036] = 16'b0000000000000000;
	sram_mem[120037] = 16'b0000000000000000;
	sram_mem[120038] = 16'b0000000000000000;
	sram_mem[120039] = 16'b0000000000000000;
	sram_mem[120040] = 16'b0000000000000000;
	sram_mem[120041] = 16'b0000000000000000;
	sram_mem[120042] = 16'b0000000000000000;
	sram_mem[120043] = 16'b0000000000000000;
	sram_mem[120044] = 16'b0000000000000000;
	sram_mem[120045] = 16'b0000000000000000;
	sram_mem[120046] = 16'b0000000000000000;
	sram_mem[120047] = 16'b0000000000000000;
	sram_mem[120048] = 16'b0000000000000000;
	sram_mem[120049] = 16'b0000000000000000;
	sram_mem[120050] = 16'b0000000000000000;
	sram_mem[120051] = 16'b0000000000000000;
	sram_mem[120052] = 16'b0000000000000000;
	sram_mem[120053] = 16'b0000000000000000;
	sram_mem[120054] = 16'b0000000000000000;
	sram_mem[120055] = 16'b0000000000000000;
	sram_mem[120056] = 16'b0000000000000000;
	sram_mem[120057] = 16'b0000000000000000;
	sram_mem[120058] = 16'b0000000000000000;
	sram_mem[120059] = 16'b0000000000000000;
	sram_mem[120060] = 16'b0000000000000000;
	sram_mem[120061] = 16'b0000000000000000;
	sram_mem[120062] = 16'b0000000000000000;
	sram_mem[120063] = 16'b0000000000000000;
	sram_mem[120064] = 16'b0000000000000000;
	sram_mem[120065] = 16'b0000000000000000;
	sram_mem[120066] = 16'b0000000000000000;
	sram_mem[120067] = 16'b0000000000000000;
	sram_mem[120068] = 16'b0000000000000000;
	sram_mem[120069] = 16'b0000000000000000;
	sram_mem[120070] = 16'b0000000000000000;
	sram_mem[120071] = 16'b0000000000000000;
	sram_mem[120072] = 16'b0000000000000000;
	sram_mem[120073] = 16'b0000000000000000;
	sram_mem[120074] = 16'b0000000000000000;
	sram_mem[120075] = 16'b0000000000000000;
	sram_mem[120076] = 16'b0000000000000000;
	sram_mem[120077] = 16'b0000000000000000;
	sram_mem[120078] = 16'b0000000000000000;
	sram_mem[120079] = 16'b0000000000000000;
	sram_mem[120080] = 16'b0000000000000000;
	sram_mem[120081] = 16'b0000000000000000;
	sram_mem[120082] = 16'b0000000000000000;
	sram_mem[120083] = 16'b0000000000000000;
	sram_mem[120084] = 16'b0000000000000000;
	sram_mem[120085] = 16'b0000000000000000;
	sram_mem[120086] = 16'b0000000000000000;
	sram_mem[120087] = 16'b0000000000000000;
	sram_mem[120088] = 16'b0000000000000000;
	sram_mem[120089] = 16'b0000000000000000;
	sram_mem[120090] = 16'b0000000000000000;
	sram_mem[120091] = 16'b0000000000000000;
	sram_mem[120092] = 16'b0000000000000000;
	sram_mem[120093] = 16'b0000000000000000;
	sram_mem[120094] = 16'b0000000000000000;
	sram_mem[120095] = 16'b0000000000000000;
	sram_mem[120096] = 16'b0000000000000000;
	sram_mem[120097] = 16'b0000000000000000;
	sram_mem[120098] = 16'b0000000000000000;
	sram_mem[120099] = 16'b0000000000000000;
	sram_mem[120100] = 16'b0000000000000000;
	sram_mem[120101] = 16'b0000000000000000;
	sram_mem[120102] = 16'b0000000000000000;
	sram_mem[120103] = 16'b0000000000000000;
	sram_mem[120104] = 16'b0000000000000000;
	sram_mem[120105] = 16'b0000000000000000;
	sram_mem[120106] = 16'b0000000000000000;
	sram_mem[120107] = 16'b0000000000000000;
	sram_mem[120108] = 16'b0000000000000000;
	sram_mem[120109] = 16'b0000000000000000;
	sram_mem[120110] = 16'b0000000000000000;
	sram_mem[120111] = 16'b0000000000000000;
	sram_mem[120112] = 16'b0000000000000000;
	sram_mem[120113] = 16'b0000000000000000;
	sram_mem[120114] = 16'b0000000000000000;
	sram_mem[120115] = 16'b0000000000000000;
	sram_mem[120116] = 16'b0000000000000000;
	sram_mem[120117] = 16'b0000000000000000;
	sram_mem[120118] = 16'b0000000000000000;
	sram_mem[120119] = 16'b0000000000000000;
	sram_mem[120120] = 16'b0000000000000000;
	sram_mem[120121] = 16'b0000000000000000;
	sram_mem[120122] = 16'b0000000000000000;
	sram_mem[120123] = 16'b0000000000000000;
	sram_mem[120124] = 16'b0000000000000000;
	sram_mem[120125] = 16'b0000000000000000;
	sram_mem[120126] = 16'b0000000000000000;
	sram_mem[120127] = 16'b0000000000000000;
	sram_mem[120128] = 16'b0000000000000000;
	sram_mem[120129] = 16'b0000000000000000;
	sram_mem[120130] = 16'b0000000000000000;
	sram_mem[120131] = 16'b0000000000000000;
	sram_mem[120132] = 16'b0000000000000000;
	sram_mem[120133] = 16'b0000000000000000;
	sram_mem[120134] = 16'b0000000000000000;
	sram_mem[120135] = 16'b0000000000000000;
	sram_mem[120136] = 16'b0000000000000000;
	sram_mem[120137] = 16'b0000000000000000;
	sram_mem[120138] = 16'b0000000000000000;
	sram_mem[120139] = 16'b0000000000000000;
	sram_mem[120140] = 16'b0000000000000000;
	sram_mem[120141] = 16'b0000000000000000;
	sram_mem[120142] = 16'b0000000000000000;
	sram_mem[120143] = 16'b0000000000000000;
	sram_mem[120144] = 16'b0000000000000000;
	sram_mem[120145] = 16'b0000000000000000;
	sram_mem[120146] = 16'b0000000000000000;
	sram_mem[120147] = 16'b0000000000000000;
	sram_mem[120148] = 16'b0000000000000000;
	sram_mem[120149] = 16'b0000000000000000;
	sram_mem[120150] = 16'b0000000000000000;
	sram_mem[120151] = 16'b0000000000000000;
	sram_mem[120152] = 16'b0000000000000000;
	sram_mem[120153] = 16'b0000000000000000;
	sram_mem[120154] = 16'b0000000000000000;
	sram_mem[120155] = 16'b0000000000000000;
	sram_mem[120156] = 16'b0000000000000000;
	sram_mem[120157] = 16'b0000000000000000;
	sram_mem[120158] = 16'b0000000000000000;
	sram_mem[120159] = 16'b0000000000000000;
	sram_mem[120160] = 16'b0000000000000000;
	sram_mem[120161] = 16'b0000000000000000;
	sram_mem[120162] = 16'b0000000000000000;
	sram_mem[120163] = 16'b0000000000000000;
	sram_mem[120164] = 16'b0000000000000000;
	sram_mem[120165] = 16'b0000000000000000;
	sram_mem[120166] = 16'b0000000000000000;
	sram_mem[120167] = 16'b0000000000000000;
	sram_mem[120168] = 16'b0000000000000000;
	sram_mem[120169] = 16'b0000000000000000;
	sram_mem[120170] = 16'b0000000000000000;
	sram_mem[120171] = 16'b0000000000000000;
	sram_mem[120172] = 16'b0000000000000000;
	sram_mem[120173] = 16'b0000000000000000;
	sram_mem[120174] = 16'b0000000000000000;
	sram_mem[120175] = 16'b0000000000000000;
	sram_mem[120176] = 16'b0000000000000000;
	sram_mem[120177] = 16'b0000000000000000;
	sram_mem[120178] = 16'b0000000000000000;
	sram_mem[120179] = 16'b0000000000000000;
	sram_mem[120180] = 16'b0000000000000000;
	sram_mem[120181] = 16'b0000000000000000;
	sram_mem[120182] = 16'b0000000000000000;
	sram_mem[120183] = 16'b0000000000000000;
	sram_mem[120184] = 16'b0000000000000000;
	sram_mem[120185] = 16'b0000000000000000;
	sram_mem[120186] = 16'b0000000000000000;
	sram_mem[120187] = 16'b0000000000000000;
	sram_mem[120188] = 16'b0000000000000000;
	sram_mem[120189] = 16'b0000000000000000;
	sram_mem[120190] = 16'b0000000000000000;
	sram_mem[120191] = 16'b0000000000000000;
	sram_mem[120192] = 16'b0000000000000000;
	sram_mem[120193] = 16'b0000000000000000;
	sram_mem[120194] = 16'b0000000000000000;
	sram_mem[120195] = 16'b0000000000000000;
	sram_mem[120196] = 16'b0000000000000000;
	sram_mem[120197] = 16'b0000000000000000;
	sram_mem[120198] = 16'b0000000000000000;
	sram_mem[120199] = 16'b0000000000000000;
	sram_mem[120200] = 16'b0000000000000000;
	sram_mem[120201] = 16'b0000000000000000;
	sram_mem[120202] = 16'b0000000000000000;
	sram_mem[120203] = 16'b0000000000000000;
	sram_mem[120204] = 16'b0000000000000000;
	sram_mem[120205] = 16'b0000000000000000;
	sram_mem[120206] = 16'b0000000000000000;
	sram_mem[120207] = 16'b0000000000000000;
	sram_mem[120208] = 16'b0000000000000000;
	sram_mem[120209] = 16'b0000000000000000;
	sram_mem[120210] = 16'b0000000000000000;
	sram_mem[120211] = 16'b0000000000000000;
	sram_mem[120212] = 16'b0000000000000000;
	sram_mem[120213] = 16'b0000000000000000;
	sram_mem[120214] = 16'b0000000000000000;
	sram_mem[120215] = 16'b0000000000000000;
	sram_mem[120216] = 16'b0000000000000000;
	sram_mem[120217] = 16'b0000000000000000;
	sram_mem[120218] = 16'b0000000000000000;
	sram_mem[120219] = 16'b0000000000000000;
	sram_mem[120220] = 16'b0000000000000000;
	sram_mem[120221] = 16'b0000000000000000;
	sram_mem[120222] = 16'b0000000000000000;
	sram_mem[120223] = 16'b0000000000000000;
	sram_mem[120224] = 16'b0000000000000000;
	sram_mem[120225] = 16'b0000000000000000;
	sram_mem[120226] = 16'b0000000000000000;
	sram_mem[120227] = 16'b0000000000000000;
	sram_mem[120228] = 16'b0000000000000000;
	sram_mem[120229] = 16'b0000000000000000;
	sram_mem[120230] = 16'b0000000000000000;
	sram_mem[120231] = 16'b0000000000000000;
	sram_mem[120232] = 16'b0000000000000000;
	sram_mem[120233] = 16'b0000000000000000;
	sram_mem[120234] = 16'b0000000000000000;
	sram_mem[120235] = 16'b0000000000000000;
	sram_mem[120236] = 16'b0000000000000000;
	sram_mem[120237] = 16'b0000000000000000;
	sram_mem[120238] = 16'b0000000000000000;
	sram_mem[120239] = 16'b0000000000000000;
	sram_mem[120240] = 16'b0000000000000000;
	sram_mem[120241] = 16'b0000000000000000;
	sram_mem[120242] = 16'b0000000000000000;
	sram_mem[120243] = 16'b0000000000000000;
	sram_mem[120244] = 16'b0000000000000000;
	sram_mem[120245] = 16'b0000000000000000;
	sram_mem[120246] = 16'b0000000000000000;
	sram_mem[120247] = 16'b0000000000000000;
	sram_mem[120248] = 16'b0000000000000000;
	sram_mem[120249] = 16'b0000000000000000;
	sram_mem[120250] = 16'b0000000000000000;
	sram_mem[120251] = 16'b0000000000000000;
	sram_mem[120252] = 16'b0000000000000000;
	sram_mem[120253] = 16'b0000000000000000;
	sram_mem[120254] = 16'b0000000000000000;
	sram_mem[120255] = 16'b0000000000000000;
	sram_mem[120256] = 16'b0000000000000000;
	sram_mem[120257] = 16'b0000000000000000;
	sram_mem[120258] = 16'b0000000000000000;
	sram_mem[120259] = 16'b0000000000000000;
	sram_mem[120260] = 16'b0000000000000000;
	sram_mem[120261] = 16'b0000000000000000;
	sram_mem[120262] = 16'b0000000000000000;
	sram_mem[120263] = 16'b0000000000000000;
	sram_mem[120264] = 16'b0000000000000000;
	sram_mem[120265] = 16'b0000000000000000;
	sram_mem[120266] = 16'b0000000000000000;
	sram_mem[120267] = 16'b0000000000000000;
	sram_mem[120268] = 16'b0000000000000000;
	sram_mem[120269] = 16'b0000000000000000;
	sram_mem[120270] = 16'b0000000000000000;
	sram_mem[120271] = 16'b0000000000000000;
	sram_mem[120272] = 16'b0000000000000000;
	sram_mem[120273] = 16'b0000000000000000;
	sram_mem[120274] = 16'b0000000000000000;
	sram_mem[120275] = 16'b0000000000000000;
	sram_mem[120276] = 16'b0000000000000000;
	sram_mem[120277] = 16'b0000000000000000;
	sram_mem[120278] = 16'b0000000000000000;
	sram_mem[120279] = 16'b0000000000000000;
	sram_mem[120280] = 16'b0000000000000000;
	sram_mem[120281] = 16'b0000000000000000;
	sram_mem[120282] = 16'b0000000000000000;
	sram_mem[120283] = 16'b0000000000000000;
	sram_mem[120284] = 16'b0000000000000000;
	sram_mem[120285] = 16'b0000000000000000;
	sram_mem[120286] = 16'b0000000000000000;
	sram_mem[120287] = 16'b0000000000000000;
	sram_mem[120288] = 16'b0000000000000000;
	sram_mem[120289] = 16'b0000000000000000;
	sram_mem[120290] = 16'b0000000000000000;
	sram_mem[120291] = 16'b0000000000000000;
	sram_mem[120292] = 16'b0000000000000000;
	sram_mem[120293] = 16'b0000000000000000;
	sram_mem[120294] = 16'b0000000000000000;
	sram_mem[120295] = 16'b0000000000000000;
	sram_mem[120296] = 16'b0000000000000000;
	sram_mem[120297] = 16'b0000000000000000;
	sram_mem[120298] = 16'b0000000000000000;
	sram_mem[120299] = 16'b0000000000000000;
	sram_mem[120300] = 16'b0000000000000000;
	sram_mem[120301] = 16'b0000000000000000;
	sram_mem[120302] = 16'b0000000000000000;
	sram_mem[120303] = 16'b0000000000000000;
	sram_mem[120304] = 16'b0000000000000000;
	sram_mem[120305] = 16'b0000000000000000;
	sram_mem[120306] = 16'b0000000000000000;
	sram_mem[120307] = 16'b0000000000000000;
	sram_mem[120308] = 16'b0000000000000000;
	sram_mem[120309] = 16'b0000000000000000;
	sram_mem[120310] = 16'b0000000000000000;
	sram_mem[120311] = 16'b0000000000000000;
	sram_mem[120312] = 16'b0000000000000000;
	sram_mem[120313] = 16'b0000000000000000;
	sram_mem[120314] = 16'b0000000000000000;
	sram_mem[120315] = 16'b0000000000000000;
	sram_mem[120316] = 16'b0000000000000000;
	sram_mem[120317] = 16'b0000000000000000;
	sram_mem[120318] = 16'b0000000000000000;
	sram_mem[120319] = 16'b0000000000000000;
	sram_mem[120320] = 16'b0000000000000000;
	sram_mem[120321] = 16'b0000000000000000;
	sram_mem[120322] = 16'b0000000000000000;
	sram_mem[120323] = 16'b0000000000000000;
	sram_mem[120324] = 16'b0000000000000000;
	sram_mem[120325] = 16'b0000000000000000;
	sram_mem[120326] = 16'b0000000000000000;
	sram_mem[120327] = 16'b0000000000000000;
	sram_mem[120328] = 16'b0000000000000000;
	sram_mem[120329] = 16'b0000000000000000;
	sram_mem[120330] = 16'b0000000000000000;
	sram_mem[120331] = 16'b0000000000000000;
	sram_mem[120332] = 16'b0000000000000000;
	sram_mem[120333] = 16'b0000000000000000;
	sram_mem[120334] = 16'b0000000000000000;
	sram_mem[120335] = 16'b0000000000000000;
	sram_mem[120336] = 16'b0000000000000000;
	sram_mem[120337] = 16'b0000000000000000;
	sram_mem[120338] = 16'b0000000000000000;
	sram_mem[120339] = 16'b0000000000000000;
	sram_mem[120340] = 16'b0000000000000000;
	sram_mem[120341] = 16'b0000000000000000;
	sram_mem[120342] = 16'b0000000000000000;
	sram_mem[120343] = 16'b0000000000000000;
	sram_mem[120344] = 16'b0000000000000000;
	sram_mem[120345] = 16'b0000000000000000;
	sram_mem[120346] = 16'b0000000000000000;
	sram_mem[120347] = 16'b0000000000000000;
	sram_mem[120348] = 16'b0000000000000000;
	sram_mem[120349] = 16'b0000000000000000;
	sram_mem[120350] = 16'b0000000000000000;
	sram_mem[120351] = 16'b0000000000000000;
	sram_mem[120352] = 16'b0000000000000000;
	sram_mem[120353] = 16'b0000000000000000;
	sram_mem[120354] = 16'b0000000000000000;
	sram_mem[120355] = 16'b0000000000000000;
	sram_mem[120356] = 16'b0000000000000000;
	sram_mem[120357] = 16'b0000000000000000;
	sram_mem[120358] = 16'b0000000000000000;
	sram_mem[120359] = 16'b0000000000000000;
	sram_mem[120360] = 16'b0000000000000000;
	sram_mem[120361] = 16'b0000000000000000;
	sram_mem[120362] = 16'b0000000000000000;
	sram_mem[120363] = 16'b0000000000000000;
	sram_mem[120364] = 16'b0000000000000000;
	sram_mem[120365] = 16'b0000000000000000;
	sram_mem[120366] = 16'b0000000000000000;
	sram_mem[120367] = 16'b0000000000000000;
	sram_mem[120368] = 16'b0000000000000000;
	sram_mem[120369] = 16'b0000000000000000;
	sram_mem[120370] = 16'b0000000000000000;
	sram_mem[120371] = 16'b0000000000000000;
	sram_mem[120372] = 16'b0000000000000000;
	sram_mem[120373] = 16'b0000000000000000;
	sram_mem[120374] = 16'b0000000000000000;
	sram_mem[120375] = 16'b0000000000000000;
	sram_mem[120376] = 16'b0000000000000000;
	sram_mem[120377] = 16'b0000000000000000;
	sram_mem[120378] = 16'b0000000000000000;
	sram_mem[120379] = 16'b0000000000000000;
	sram_mem[120380] = 16'b0000000000000000;
	sram_mem[120381] = 16'b0000000000000000;
	sram_mem[120382] = 16'b0000000000000000;
	sram_mem[120383] = 16'b0000000000000000;
	sram_mem[120384] = 16'b0000000000000000;
	sram_mem[120385] = 16'b0000000000000000;
	sram_mem[120386] = 16'b0000000000000000;
	sram_mem[120387] = 16'b0000000000000000;
	sram_mem[120388] = 16'b0000000000000000;
	sram_mem[120389] = 16'b0000000000000000;
	sram_mem[120390] = 16'b0000000000000000;
	sram_mem[120391] = 16'b0000000000000000;
	sram_mem[120392] = 16'b0000000000000000;
	sram_mem[120393] = 16'b0000000000000000;
	sram_mem[120394] = 16'b0000000000000000;
	sram_mem[120395] = 16'b0000000000000000;
	sram_mem[120396] = 16'b0000000000000000;
	sram_mem[120397] = 16'b0000000000000000;
	sram_mem[120398] = 16'b0000000000000000;
	sram_mem[120399] = 16'b0000000000000000;
	sram_mem[120400] = 16'b0000000000000000;
	sram_mem[120401] = 16'b0000000000000000;
	sram_mem[120402] = 16'b0000000000000000;
	sram_mem[120403] = 16'b0000000000000000;
	sram_mem[120404] = 16'b0000000000000000;
	sram_mem[120405] = 16'b0000000000000000;
	sram_mem[120406] = 16'b0000000000000000;
	sram_mem[120407] = 16'b0000000000000000;
	sram_mem[120408] = 16'b0000000000000000;
	sram_mem[120409] = 16'b0000000000000000;
	sram_mem[120410] = 16'b0000000000000000;
	sram_mem[120411] = 16'b0000000000000000;
	sram_mem[120412] = 16'b0000000000000000;
	sram_mem[120413] = 16'b0000000000000000;
	sram_mem[120414] = 16'b0000000000000000;
	sram_mem[120415] = 16'b0000000000000000;
	sram_mem[120416] = 16'b0000000000000000;
	sram_mem[120417] = 16'b0000000000000000;
	sram_mem[120418] = 16'b0000000000000000;
	sram_mem[120419] = 16'b0000000000000000;
	sram_mem[120420] = 16'b0000000000000000;
	sram_mem[120421] = 16'b0000000000000000;
	sram_mem[120422] = 16'b0000000000000000;
	sram_mem[120423] = 16'b0000000000000000;
	sram_mem[120424] = 16'b0000000000000000;
	sram_mem[120425] = 16'b0000000000000000;
	sram_mem[120426] = 16'b0000000000000000;
	sram_mem[120427] = 16'b0000000000000000;
	sram_mem[120428] = 16'b0000000000000000;
	sram_mem[120429] = 16'b0000000000000000;
	sram_mem[120430] = 16'b0000000000000000;
	sram_mem[120431] = 16'b0000000000000000;
	sram_mem[120432] = 16'b0000000000000000;
	sram_mem[120433] = 16'b0000000000000000;
	sram_mem[120434] = 16'b0000000000000000;
	sram_mem[120435] = 16'b0000000000000000;
	sram_mem[120436] = 16'b0000000000000000;
	sram_mem[120437] = 16'b0000000000000000;
	sram_mem[120438] = 16'b0000000000000000;
	sram_mem[120439] = 16'b0000000000000000;
	sram_mem[120440] = 16'b0000000000000000;
	sram_mem[120441] = 16'b0000000000000000;
	sram_mem[120442] = 16'b0000000000000000;
	sram_mem[120443] = 16'b0000000000000000;
	sram_mem[120444] = 16'b0000000000000000;
	sram_mem[120445] = 16'b0000000000000000;
	sram_mem[120446] = 16'b0000000000000000;
	sram_mem[120447] = 16'b0000000000000000;
	sram_mem[120448] = 16'b0000000000000000;
	sram_mem[120449] = 16'b0000000000000000;
	sram_mem[120450] = 16'b0000000000000000;
	sram_mem[120451] = 16'b0000000000000000;
	sram_mem[120452] = 16'b0000000000000000;
	sram_mem[120453] = 16'b0000000000000000;
	sram_mem[120454] = 16'b0000000000000000;
	sram_mem[120455] = 16'b0000000000000000;
	sram_mem[120456] = 16'b0000000000000000;
	sram_mem[120457] = 16'b0000000000000000;
	sram_mem[120458] = 16'b0000000000000000;
	sram_mem[120459] = 16'b0000000000000000;
	sram_mem[120460] = 16'b0000000000000000;
	sram_mem[120461] = 16'b0000000000000000;
	sram_mem[120462] = 16'b0000000000000000;
	sram_mem[120463] = 16'b0000000000000000;
	sram_mem[120464] = 16'b0000000000000000;
	sram_mem[120465] = 16'b0000000000000000;
	sram_mem[120466] = 16'b0000000000000000;
	sram_mem[120467] = 16'b0000000000000000;
	sram_mem[120468] = 16'b0000000000000000;
	sram_mem[120469] = 16'b0000000000000000;
	sram_mem[120470] = 16'b0000000000000000;
	sram_mem[120471] = 16'b0000000000000000;
	sram_mem[120472] = 16'b0000000000000000;
	sram_mem[120473] = 16'b0000000000000000;
	sram_mem[120474] = 16'b0000000000000000;
	sram_mem[120475] = 16'b0000000000000000;
	sram_mem[120476] = 16'b0000000000000000;
	sram_mem[120477] = 16'b0000000000000000;
	sram_mem[120478] = 16'b0000000000000000;
	sram_mem[120479] = 16'b0000000000000000;
	sram_mem[120480] = 16'b0000000000000000;
	sram_mem[120481] = 16'b0000000000000000;
	sram_mem[120482] = 16'b0000000000000000;
	sram_mem[120483] = 16'b0000000000000000;
	sram_mem[120484] = 16'b0000000000000000;
	sram_mem[120485] = 16'b0000000000000000;
	sram_mem[120486] = 16'b0000000000000000;
	sram_mem[120487] = 16'b0000000000000000;
	sram_mem[120488] = 16'b0000000000000000;
	sram_mem[120489] = 16'b0000000000000000;
	sram_mem[120490] = 16'b0000000000000000;
	sram_mem[120491] = 16'b0000000000000000;
	sram_mem[120492] = 16'b0000000000000000;
	sram_mem[120493] = 16'b0000000000000000;
	sram_mem[120494] = 16'b0000000000000000;
	sram_mem[120495] = 16'b0000000000000000;
	sram_mem[120496] = 16'b0000000000000000;
	sram_mem[120497] = 16'b0000000000000000;
	sram_mem[120498] = 16'b0000000000000000;
	sram_mem[120499] = 16'b0000000000000000;
	sram_mem[120500] = 16'b0000000000000000;
	sram_mem[120501] = 16'b0000000000000000;
	sram_mem[120502] = 16'b0000000000000000;
	sram_mem[120503] = 16'b0000000000000000;
	sram_mem[120504] = 16'b0000000000000000;
	sram_mem[120505] = 16'b0000000000000000;
	sram_mem[120506] = 16'b0000000000000000;
	sram_mem[120507] = 16'b0000000000000000;
	sram_mem[120508] = 16'b0000000000000000;
	sram_mem[120509] = 16'b0000000000000000;
	sram_mem[120510] = 16'b0000000000000000;
	sram_mem[120511] = 16'b0000000000000000;
	sram_mem[120512] = 16'b0000000000000000;
	sram_mem[120513] = 16'b0000000000000000;
	sram_mem[120514] = 16'b0000000000000000;
	sram_mem[120515] = 16'b0000000000000000;
	sram_mem[120516] = 16'b0000000000000000;
	sram_mem[120517] = 16'b0000000000000000;
	sram_mem[120518] = 16'b0000000000000000;
	sram_mem[120519] = 16'b0000000000000000;
	sram_mem[120520] = 16'b0000000000000000;
	sram_mem[120521] = 16'b0000000000000000;
	sram_mem[120522] = 16'b0000000000000000;
	sram_mem[120523] = 16'b0000000000000000;
	sram_mem[120524] = 16'b0000000000000000;
	sram_mem[120525] = 16'b0000000000000000;
	sram_mem[120526] = 16'b0000000000000000;
	sram_mem[120527] = 16'b0000000000000000;
	sram_mem[120528] = 16'b0000000000000000;
	sram_mem[120529] = 16'b0000000000000000;
	sram_mem[120530] = 16'b0000000000000000;
	sram_mem[120531] = 16'b0000000000000000;
	sram_mem[120532] = 16'b0000000000000000;
	sram_mem[120533] = 16'b0000000000000000;
	sram_mem[120534] = 16'b0000000000000000;
	sram_mem[120535] = 16'b0000000000000000;
	sram_mem[120536] = 16'b0000000000000000;
	sram_mem[120537] = 16'b0000000000000000;
	sram_mem[120538] = 16'b0000000000000000;
	sram_mem[120539] = 16'b0000000000000000;
	sram_mem[120540] = 16'b0000000000000000;
	sram_mem[120541] = 16'b0000000000000000;
	sram_mem[120542] = 16'b0000000000000000;
	sram_mem[120543] = 16'b0000000000000000;
	sram_mem[120544] = 16'b0000000000000000;
	sram_mem[120545] = 16'b0000000000000000;
	sram_mem[120546] = 16'b0000000000000000;
	sram_mem[120547] = 16'b0000000000000000;
	sram_mem[120548] = 16'b0000000000000000;
	sram_mem[120549] = 16'b0000000000000000;
	sram_mem[120550] = 16'b0000000000000000;
	sram_mem[120551] = 16'b0000000000000000;
	sram_mem[120552] = 16'b0000000000000000;
	sram_mem[120553] = 16'b0000000000000000;
	sram_mem[120554] = 16'b0000000000000000;
	sram_mem[120555] = 16'b0000000000000000;
	sram_mem[120556] = 16'b0000000000000000;
	sram_mem[120557] = 16'b0000000000000000;
	sram_mem[120558] = 16'b0000000000000000;
	sram_mem[120559] = 16'b0000000000000000;
	sram_mem[120560] = 16'b0000000000000000;
	sram_mem[120561] = 16'b0000000000000000;
	sram_mem[120562] = 16'b0000000000000000;
	sram_mem[120563] = 16'b0000000000000000;
	sram_mem[120564] = 16'b0000000000000000;
	sram_mem[120565] = 16'b0000000000000000;
	sram_mem[120566] = 16'b0000000000000000;
	sram_mem[120567] = 16'b0000000000000000;
	sram_mem[120568] = 16'b0000000000000000;
	sram_mem[120569] = 16'b0000000000000000;
	sram_mem[120570] = 16'b0000000000000000;
	sram_mem[120571] = 16'b0000000000000000;
	sram_mem[120572] = 16'b0000000000000000;
	sram_mem[120573] = 16'b0000000000000000;
	sram_mem[120574] = 16'b0000000000000000;
	sram_mem[120575] = 16'b0000000000000000;
	sram_mem[120576] = 16'b0000000000000000;
	sram_mem[120577] = 16'b0000000000000000;
	sram_mem[120578] = 16'b0000000000000000;
	sram_mem[120579] = 16'b0000000000000000;
	sram_mem[120580] = 16'b0000000000000000;
	sram_mem[120581] = 16'b0000000000000000;
	sram_mem[120582] = 16'b0000000000000000;
	sram_mem[120583] = 16'b0000000000000000;
	sram_mem[120584] = 16'b0000000000000000;
	sram_mem[120585] = 16'b0000000000000000;
	sram_mem[120586] = 16'b0000000000000000;
	sram_mem[120587] = 16'b0000000000000000;
	sram_mem[120588] = 16'b0000000000000000;
	sram_mem[120589] = 16'b0000000000000000;
	sram_mem[120590] = 16'b0000000000000000;
	sram_mem[120591] = 16'b0000000000000000;
	sram_mem[120592] = 16'b0000000000000000;
	sram_mem[120593] = 16'b0000000000000000;
	sram_mem[120594] = 16'b0000000000000000;
	sram_mem[120595] = 16'b0000000000000000;
	sram_mem[120596] = 16'b0000000000000000;
	sram_mem[120597] = 16'b0000000000000000;
	sram_mem[120598] = 16'b0000000000000000;
	sram_mem[120599] = 16'b0000000000000000;
	sram_mem[120600] = 16'b0000000000000000;
	sram_mem[120601] = 16'b0000000000000000;
	sram_mem[120602] = 16'b0000000000000000;
	sram_mem[120603] = 16'b0000000000000000;
	sram_mem[120604] = 16'b0000000000000000;
	sram_mem[120605] = 16'b0000000000000000;
	sram_mem[120606] = 16'b0000000000000000;
	sram_mem[120607] = 16'b0000000000000000;
	sram_mem[120608] = 16'b0000000000000000;
	sram_mem[120609] = 16'b0000000000000000;
	sram_mem[120610] = 16'b0000000000000000;
	sram_mem[120611] = 16'b0000000000000000;
	sram_mem[120612] = 16'b0000000000000000;
	sram_mem[120613] = 16'b0000000000000000;
	sram_mem[120614] = 16'b0000000000000000;
	sram_mem[120615] = 16'b0000000000000000;
	sram_mem[120616] = 16'b0000000000000000;
	sram_mem[120617] = 16'b0000000000000000;
	sram_mem[120618] = 16'b0000000000000000;
	sram_mem[120619] = 16'b0000000000000000;
	sram_mem[120620] = 16'b0000000000000000;
	sram_mem[120621] = 16'b0000000000000000;
	sram_mem[120622] = 16'b0000000000000000;
	sram_mem[120623] = 16'b0000000000000000;
	sram_mem[120624] = 16'b0000000000000000;
	sram_mem[120625] = 16'b0000000000000000;
	sram_mem[120626] = 16'b0000000000000000;
	sram_mem[120627] = 16'b0000000000000000;
	sram_mem[120628] = 16'b0000000000000000;
	sram_mem[120629] = 16'b0000000000000000;
	sram_mem[120630] = 16'b0000000000000000;
	sram_mem[120631] = 16'b0000000000000000;
	sram_mem[120632] = 16'b0000000000000000;
	sram_mem[120633] = 16'b0000000000000000;
	sram_mem[120634] = 16'b0000000000000000;
	sram_mem[120635] = 16'b0000000000000000;
	sram_mem[120636] = 16'b0000000000000000;
	sram_mem[120637] = 16'b0000000000000000;
	sram_mem[120638] = 16'b0000000000000000;
	sram_mem[120639] = 16'b0000000000000000;
	sram_mem[120640] = 16'b0000000000000000;
	sram_mem[120641] = 16'b0000000000000000;
	sram_mem[120642] = 16'b0000000000000000;
	sram_mem[120643] = 16'b0000000000000000;
	sram_mem[120644] = 16'b0000000000000000;
	sram_mem[120645] = 16'b0000000000000000;
	sram_mem[120646] = 16'b0000000000000000;
	sram_mem[120647] = 16'b0000000000000000;
	sram_mem[120648] = 16'b0000000000000000;
	sram_mem[120649] = 16'b0000000000000000;
	sram_mem[120650] = 16'b0000000000000000;
	sram_mem[120651] = 16'b0000000000000000;
	sram_mem[120652] = 16'b0000000000000000;
	sram_mem[120653] = 16'b0000000000000000;
	sram_mem[120654] = 16'b0000000000000000;
	sram_mem[120655] = 16'b0000000000000000;
	sram_mem[120656] = 16'b0000000000000000;
	sram_mem[120657] = 16'b0000000000000000;
	sram_mem[120658] = 16'b0000000000000000;
	sram_mem[120659] = 16'b0000000000000000;
	sram_mem[120660] = 16'b0000000000000000;
	sram_mem[120661] = 16'b0000000000000000;
	sram_mem[120662] = 16'b0000000000000000;
	sram_mem[120663] = 16'b0000000000000000;
	sram_mem[120664] = 16'b0000000000000000;
	sram_mem[120665] = 16'b0000000000000000;
	sram_mem[120666] = 16'b0000000000000000;
	sram_mem[120667] = 16'b0000000000000000;
	sram_mem[120668] = 16'b0000000000000000;
	sram_mem[120669] = 16'b0000000000000000;
	sram_mem[120670] = 16'b0000000000000000;
	sram_mem[120671] = 16'b0000000000000000;
	sram_mem[120672] = 16'b0000000000000000;
	sram_mem[120673] = 16'b0000000000000000;
	sram_mem[120674] = 16'b0000000000000000;
	sram_mem[120675] = 16'b0000000000000000;
	sram_mem[120676] = 16'b0000000000000000;
	sram_mem[120677] = 16'b0000000000000000;
	sram_mem[120678] = 16'b0000000000000000;
	sram_mem[120679] = 16'b0000000000000000;
	sram_mem[120680] = 16'b0000000000000000;
	sram_mem[120681] = 16'b0000000000000000;
	sram_mem[120682] = 16'b0000000000000000;
	sram_mem[120683] = 16'b0000000000000000;
	sram_mem[120684] = 16'b0000000000000000;
	sram_mem[120685] = 16'b0000000000000000;
	sram_mem[120686] = 16'b0000000000000000;
	sram_mem[120687] = 16'b0000000000000000;
	sram_mem[120688] = 16'b0000000000000000;
	sram_mem[120689] = 16'b0000000000000000;
	sram_mem[120690] = 16'b0000000000000000;
	sram_mem[120691] = 16'b0000000000000000;
	sram_mem[120692] = 16'b0000000000000000;
	sram_mem[120693] = 16'b0000000000000000;
	sram_mem[120694] = 16'b0000000000000000;
	sram_mem[120695] = 16'b0000000000000000;
	sram_mem[120696] = 16'b0000000000000000;
	sram_mem[120697] = 16'b0000000000000000;
	sram_mem[120698] = 16'b0000000000000000;
	sram_mem[120699] = 16'b0000000000000000;
	sram_mem[120700] = 16'b0000000000000000;
	sram_mem[120701] = 16'b0000000000000000;
	sram_mem[120702] = 16'b0000000000000000;
	sram_mem[120703] = 16'b0000000000000000;
	sram_mem[120704] = 16'b0000000000000000;
	sram_mem[120705] = 16'b0000000000000000;
	sram_mem[120706] = 16'b0000000000000000;
	sram_mem[120707] = 16'b0000000000000000;
	sram_mem[120708] = 16'b0000000000000000;
	sram_mem[120709] = 16'b0000000000000000;
	sram_mem[120710] = 16'b0000000000000000;
	sram_mem[120711] = 16'b0000000000000000;
	sram_mem[120712] = 16'b0000000000000000;
	sram_mem[120713] = 16'b0000000000000000;
	sram_mem[120714] = 16'b0000000000000000;
	sram_mem[120715] = 16'b0000000000000000;
	sram_mem[120716] = 16'b0000000000000000;
	sram_mem[120717] = 16'b0000000000000000;
	sram_mem[120718] = 16'b0000000000000000;
	sram_mem[120719] = 16'b0000000000000000;
	sram_mem[120720] = 16'b0000000000000000;
	sram_mem[120721] = 16'b0000000000000000;
	sram_mem[120722] = 16'b0000000000000000;
	sram_mem[120723] = 16'b0000000000000000;
	sram_mem[120724] = 16'b0000000000000000;
	sram_mem[120725] = 16'b0000000000000000;
	sram_mem[120726] = 16'b0000000000000000;
	sram_mem[120727] = 16'b0000000000000000;
	sram_mem[120728] = 16'b0000000000000000;
	sram_mem[120729] = 16'b0000000000000000;
	sram_mem[120730] = 16'b0000000000000000;
	sram_mem[120731] = 16'b0000000000000000;
	sram_mem[120732] = 16'b0000000000000000;
	sram_mem[120733] = 16'b0000000000000000;
	sram_mem[120734] = 16'b0000000000000000;
	sram_mem[120735] = 16'b0000000000000000;
	sram_mem[120736] = 16'b0000000000000000;
	sram_mem[120737] = 16'b0000000000000000;
	sram_mem[120738] = 16'b0000000000000000;
	sram_mem[120739] = 16'b0000000000000000;
	sram_mem[120740] = 16'b0000000000000000;
	sram_mem[120741] = 16'b0000000000000000;
	sram_mem[120742] = 16'b0000000000000000;
	sram_mem[120743] = 16'b0000000000000000;
	sram_mem[120744] = 16'b0000000000000000;
	sram_mem[120745] = 16'b0000000000000000;
	sram_mem[120746] = 16'b0000000000000000;
	sram_mem[120747] = 16'b0000000000000000;
	sram_mem[120748] = 16'b0000000000000000;
	sram_mem[120749] = 16'b0000000000000000;
	sram_mem[120750] = 16'b0000000000000000;
	sram_mem[120751] = 16'b0000000000000000;
	sram_mem[120752] = 16'b0000000000000000;
	sram_mem[120753] = 16'b0000000000000000;
	sram_mem[120754] = 16'b0000000000000000;
	sram_mem[120755] = 16'b0000000000000000;
	sram_mem[120756] = 16'b0000000000000000;
	sram_mem[120757] = 16'b0000000000000000;
	sram_mem[120758] = 16'b0000000000000000;
	sram_mem[120759] = 16'b0000000000000000;
	sram_mem[120760] = 16'b0000000000000000;
	sram_mem[120761] = 16'b0000000000000000;
	sram_mem[120762] = 16'b0000000000000000;
	sram_mem[120763] = 16'b0000000000000000;
	sram_mem[120764] = 16'b0000000000000000;
	sram_mem[120765] = 16'b0000000000000000;
	sram_mem[120766] = 16'b0000000000000000;
	sram_mem[120767] = 16'b0000000000000000;
	sram_mem[120768] = 16'b0000000000000000;
	sram_mem[120769] = 16'b0000000000000000;
	sram_mem[120770] = 16'b0000000000000000;
	sram_mem[120771] = 16'b0000000000000000;
	sram_mem[120772] = 16'b0000000000000000;
	sram_mem[120773] = 16'b0000000000000000;
	sram_mem[120774] = 16'b0000000000000000;
	sram_mem[120775] = 16'b0000000000000000;
	sram_mem[120776] = 16'b0000000000000000;
	sram_mem[120777] = 16'b0000000000000000;
	sram_mem[120778] = 16'b0000000000000000;
	sram_mem[120779] = 16'b0000000000000000;
	sram_mem[120780] = 16'b0000000000000000;
	sram_mem[120781] = 16'b0000000000000000;
	sram_mem[120782] = 16'b0000000000000000;
	sram_mem[120783] = 16'b0000000000000000;
	sram_mem[120784] = 16'b0000000000000000;
	sram_mem[120785] = 16'b0000000000000000;
	sram_mem[120786] = 16'b0000000000000000;
	sram_mem[120787] = 16'b0000000000000000;
	sram_mem[120788] = 16'b0000000000000000;
	sram_mem[120789] = 16'b0000000000000000;
	sram_mem[120790] = 16'b0000000000000000;
	sram_mem[120791] = 16'b0000000000000000;
	sram_mem[120792] = 16'b0000000000000000;
	sram_mem[120793] = 16'b0000000000000000;
	sram_mem[120794] = 16'b0000000000000000;
	sram_mem[120795] = 16'b0000000000000000;
	sram_mem[120796] = 16'b0000000000000000;
	sram_mem[120797] = 16'b0000000000000000;
	sram_mem[120798] = 16'b0000000000000000;
	sram_mem[120799] = 16'b0000000000000000;
	sram_mem[120800] = 16'b0000000000000000;
	sram_mem[120801] = 16'b0000000000000000;
	sram_mem[120802] = 16'b0000000000000000;
	sram_mem[120803] = 16'b0000000000000000;
	sram_mem[120804] = 16'b0000000000000000;
	sram_mem[120805] = 16'b0000000000000000;
	sram_mem[120806] = 16'b0000000000000000;
	sram_mem[120807] = 16'b0000000000000000;
	sram_mem[120808] = 16'b0000000000000000;
	sram_mem[120809] = 16'b0000000000000000;
	sram_mem[120810] = 16'b0000000000000000;
	sram_mem[120811] = 16'b0000000000000000;
	sram_mem[120812] = 16'b0000000000000000;
	sram_mem[120813] = 16'b0000000000000000;
	sram_mem[120814] = 16'b0000000000000000;
	sram_mem[120815] = 16'b0000000000000000;
	sram_mem[120816] = 16'b0000000000000000;
	sram_mem[120817] = 16'b0000000000000000;
	sram_mem[120818] = 16'b0000000000000000;
	sram_mem[120819] = 16'b0000000000000000;
	sram_mem[120820] = 16'b0000000000000000;
	sram_mem[120821] = 16'b0000000000000000;
	sram_mem[120822] = 16'b0000000000000000;
	sram_mem[120823] = 16'b0000000000000000;
	sram_mem[120824] = 16'b0000000000000000;
	sram_mem[120825] = 16'b0000000000000000;
	sram_mem[120826] = 16'b0000000000000000;
	sram_mem[120827] = 16'b0000000000000000;
	sram_mem[120828] = 16'b0000000000000000;
	sram_mem[120829] = 16'b0000000000000000;
	sram_mem[120830] = 16'b0000000000000000;
	sram_mem[120831] = 16'b0000000000000000;
	sram_mem[120832] = 16'b0000000000000000;
	sram_mem[120833] = 16'b0000000000000000;
	sram_mem[120834] = 16'b0000000000000000;
	sram_mem[120835] = 16'b0000000000000000;
	sram_mem[120836] = 16'b0000000000000000;
	sram_mem[120837] = 16'b0000000000000000;
	sram_mem[120838] = 16'b0000000000000000;
	sram_mem[120839] = 16'b0000000000000000;
	sram_mem[120840] = 16'b0000000000000000;
	sram_mem[120841] = 16'b0000000000000000;
	sram_mem[120842] = 16'b0000000000000000;
	sram_mem[120843] = 16'b0000000000000000;
	sram_mem[120844] = 16'b0000000000000000;
	sram_mem[120845] = 16'b0000000000000000;
	sram_mem[120846] = 16'b0000000000000000;
	sram_mem[120847] = 16'b0000000000000000;
	sram_mem[120848] = 16'b0000000000000000;
	sram_mem[120849] = 16'b0000000000000000;
	sram_mem[120850] = 16'b0000000000000000;
	sram_mem[120851] = 16'b0000000000000000;
	sram_mem[120852] = 16'b0000000000000000;
	sram_mem[120853] = 16'b0000000000000000;
	sram_mem[120854] = 16'b0000000000000000;
	sram_mem[120855] = 16'b0000000000000000;
	sram_mem[120856] = 16'b0000000000000000;
	sram_mem[120857] = 16'b0000000000000000;
	sram_mem[120858] = 16'b0000000000000000;
	sram_mem[120859] = 16'b0000000000000000;
	sram_mem[120860] = 16'b0000000000000000;
	sram_mem[120861] = 16'b0000000000000000;
	sram_mem[120862] = 16'b0000000000000000;
	sram_mem[120863] = 16'b0000000000000000;
	sram_mem[120864] = 16'b0000000000000000;
	sram_mem[120865] = 16'b0000000000000000;
	sram_mem[120866] = 16'b0000000000000000;
	sram_mem[120867] = 16'b0000000000000000;
	sram_mem[120868] = 16'b0000000000000000;
	sram_mem[120869] = 16'b0000000000000000;
	sram_mem[120870] = 16'b0000000000000000;
	sram_mem[120871] = 16'b0000000000000000;
	sram_mem[120872] = 16'b0000000000000000;
	sram_mem[120873] = 16'b0000000000000000;
	sram_mem[120874] = 16'b0000000000000000;
	sram_mem[120875] = 16'b0000000000000000;
	sram_mem[120876] = 16'b0000000000000000;
	sram_mem[120877] = 16'b0000000000000000;
	sram_mem[120878] = 16'b0000000000000000;
	sram_mem[120879] = 16'b0000000000000000;
	sram_mem[120880] = 16'b0000000000000000;
	sram_mem[120881] = 16'b0000000000000000;
	sram_mem[120882] = 16'b0000000000000000;
	sram_mem[120883] = 16'b0000000000000000;
	sram_mem[120884] = 16'b0000000000000000;
	sram_mem[120885] = 16'b0000000000000000;
	sram_mem[120886] = 16'b0000000000000000;
	sram_mem[120887] = 16'b0000000000000000;
	sram_mem[120888] = 16'b0000000000000000;
	sram_mem[120889] = 16'b0000000000000000;
	sram_mem[120890] = 16'b0000000000000000;
	sram_mem[120891] = 16'b0000000000000000;
	sram_mem[120892] = 16'b0000000000000000;
	sram_mem[120893] = 16'b0000000000000000;
	sram_mem[120894] = 16'b0000000000000000;
	sram_mem[120895] = 16'b0000000000000000;
	sram_mem[120896] = 16'b0000000000000000;
	sram_mem[120897] = 16'b0000000000000000;
	sram_mem[120898] = 16'b0000000000000000;
	sram_mem[120899] = 16'b0000000000000000;
	sram_mem[120900] = 16'b0000000000000000;
	sram_mem[120901] = 16'b0000000000000000;
	sram_mem[120902] = 16'b0000000000000000;
	sram_mem[120903] = 16'b0000000000000000;
	sram_mem[120904] = 16'b0000000000000000;
	sram_mem[120905] = 16'b0000000000000000;
	sram_mem[120906] = 16'b0000000000000000;
	sram_mem[120907] = 16'b0000000000000000;
	sram_mem[120908] = 16'b0000000000000000;
	sram_mem[120909] = 16'b0000000000000000;
	sram_mem[120910] = 16'b0000000000000000;
	sram_mem[120911] = 16'b0000000000000000;
	sram_mem[120912] = 16'b0000000000000000;
	sram_mem[120913] = 16'b0000000000000000;
	sram_mem[120914] = 16'b0000000000000000;
	sram_mem[120915] = 16'b0000000000000000;
	sram_mem[120916] = 16'b0000000000000000;
	sram_mem[120917] = 16'b0000000000000000;
	sram_mem[120918] = 16'b0000000000000000;
	sram_mem[120919] = 16'b0000000000000000;
	sram_mem[120920] = 16'b0000000000000000;
	sram_mem[120921] = 16'b0000000000000000;
	sram_mem[120922] = 16'b0000000000000000;
	sram_mem[120923] = 16'b0000000000000000;
	sram_mem[120924] = 16'b0000000000000000;
	sram_mem[120925] = 16'b0000000000000000;
	sram_mem[120926] = 16'b0000000000000000;
	sram_mem[120927] = 16'b0000000000000000;
	sram_mem[120928] = 16'b0000000000000000;
	sram_mem[120929] = 16'b0000000000000000;
	sram_mem[120930] = 16'b0000000000000000;
	sram_mem[120931] = 16'b0000000000000000;
	sram_mem[120932] = 16'b0000000000000000;
	sram_mem[120933] = 16'b0000000000000000;
	sram_mem[120934] = 16'b0000000000000000;
	sram_mem[120935] = 16'b0000000000000000;
	sram_mem[120936] = 16'b0000000000000000;
	sram_mem[120937] = 16'b0000000000000000;
	sram_mem[120938] = 16'b0000000000000000;
	sram_mem[120939] = 16'b0000000000000000;
	sram_mem[120940] = 16'b0000000000000000;
	sram_mem[120941] = 16'b0000000000000000;
	sram_mem[120942] = 16'b0000000000000000;
	sram_mem[120943] = 16'b0000000000000000;
	sram_mem[120944] = 16'b0000000000000000;
	sram_mem[120945] = 16'b0000000000000000;
	sram_mem[120946] = 16'b0000000000000000;
	sram_mem[120947] = 16'b0000000000000000;
	sram_mem[120948] = 16'b0000000000000000;
	sram_mem[120949] = 16'b0000000000000000;
	sram_mem[120950] = 16'b0000000000000000;
	sram_mem[120951] = 16'b0000000000000000;
	sram_mem[120952] = 16'b0000000000000000;
	sram_mem[120953] = 16'b0000000000000000;
	sram_mem[120954] = 16'b0000000000000000;
	sram_mem[120955] = 16'b0000000000000000;
	sram_mem[120956] = 16'b0000000000000000;
	sram_mem[120957] = 16'b0000000000000000;
	sram_mem[120958] = 16'b0000000000000000;
	sram_mem[120959] = 16'b0000000000000000;
	sram_mem[120960] = 16'b0000000000000000;
	sram_mem[120961] = 16'b0000000000000000;
	sram_mem[120962] = 16'b0000000000000000;
	sram_mem[120963] = 16'b0000000000000000;
	sram_mem[120964] = 16'b0000000000000000;
	sram_mem[120965] = 16'b0000000000000000;
	sram_mem[120966] = 16'b0000000000000000;
	sram_mem[120967] = 16'b0000000000000000;
	sram_mem[120968] = 16'b0000000000000000;
	sram_mem[120969] = 16'b0000000000000000;
	sram_mem[120970] = 16'b0000000000000000;
	sram_mem[120971] = 16'b0000000000000000;
	sram_mem[120972] = 16'b0000000000000000;
	sram_mem[120973] = 16'b0000000000000000;
	sram_mem[120974] = 16'b0000000000000000;
	sram_mem[120975] = 16'b0000000000000000;
	sram_mem[120976] = 16'b0000000000000000;
	sram_mem[120977] = 16'b0000000000000000;
	sram_mem[120978] = 16'b0000000000000000;
	sram_mem[120979] = 16'b0000000000000000;
	sram_mem[120980] = 16'b0000000000000000;
	sram_mem[120981] = 16'b0000000000000000;
	sram_mem[120982] = 16'b0000000000000000;
	sram_mem[120983] = 16'b0000000000000000;
	sram_mem[120984] = 16'b0000000000000000;
	sram_mem[120985] = 16'b0000000000000000;
	sram_mem[120986] = 16'b0000000000000000;
	sram_mem[120987] = 16'b0000000000000000;
	sram_mem[120988] = 16'b0000000000000000;
	sram_mem[120989] = 16'b0000000000000000;
	sram_mem[120990] = 16'b0000000000000000;
	sram_mem[120991] = 16'b0000000000000000;
	sram_mem[120992] = 16'b0000000000000000;
	sram_mem[120993] = 16'b0000000000000000;
	sram_mem[120994] = 16'b0000000000000000;
	sram_mem[120995] = 16'b0000000000000000;
	sram_mem[120996] = 16'b0000000000000000;
	sram_mem[120997] = 16'b0000000000000000;
	sram_mem[120998] = 16'b0000000000000000;
	sram_mem[120999] = 16'b0000000000000000;
	sram_mem[121000] = 16'b0000000000000000;
	sram_mem[121001] = 16'b0000000000000000;
	sram_mem[121002] = 16'b0000000000000000;
	sram_mem[121003] = 16'b0000000000000000;
	sram_mem[121004] = 16'b0000000000000000;
	sram_mem[121005] = 16'b0000000000000000;
	sram_mem[121006] = 16'b0000000000000000;
	sram_mem[121007] = 16'b0000000000000000;
	sram_mem[121008] = 16'b0000000000000000;
	sram_mem[121009] = 16'b0000000000000000;
	sram_mem[121010] = 16'b0000000000000000;
	sram_mem[121011] = 16'b0000000000000000;
	sram_mem[121012] = 16'b0000000000000000;
	sram_mem[121013] = 16'b0000000000000000;
	sram_mem[121014] = 16'b0000000000000000;
	sram_mem[121015] = 16'b0000000000000000;
	sram_mem[121016] = 16'b0000000000000000;
	sram_mem[121017] = 16'b0000000000000000;
	sram_mem[121018] = 16'b0000000000000000;
	sram_mem[121019] = 16'b0000000000000000;
	sram_mem[121020] = 16'b0000000000000000;
	sram_mem[121021] = 16'b0000000000000000;
	sram_mem[121022] = 16'b0000000000000000;
	sram_mem[121023] = 16'b0000000000000000;
	sram_mem[121024] = 16'b0000000000000000;
	sram_mem[121025] = 16'b0000000000000000;
	sram_mem[121026] = 16'b0000000000000000;
	sram_mem[121027] = 16'b0000000000000000;
	sram_mem[121028] = 16'b0000000000000000;
	sram_mem[121029] = 16'b0000000000000000;
	sram_mem[121030] = 16'b0000000000000000;
	sram_mem[121031] = 16'b0000000000000000;
	sram_mem[121032] = 16'b0000000000000000;
	sram_mem[121033] = 16'b0000000000000000;
	sram_mem[121034] = 16'b0000000000000000;
	sram_mem[121035] = 16'b0000000000000000;
	sram_mem[121036] = 16'b0000000000000000;
	sram_mem[121037] = 16'b0000000000000000;
	sram_mem[121038] = 16'b0000000000000000;
	sram_mem[121039] = 16'b0000000000000000;
	sram_mem[121040] = 16'b0000000000000000;
	sram_mem[121041] = 16'b0000000000000000;
	sram_mem[121042] = 16'b0000000000000000;
	sram_mem[121043] = 16'b0000000000000000;
	sram_mem[121044] = 16'b0000000000000000;
	sram_mem[121045] = 16'b0000000000000000;
	sram_mem[121046] = 16'b0000000000000000;
	sram_mem[121047] = 16'b0000000000000000;
	sram_mem[121048] = 16'b0000000000000000;
	sram_mem[121049] = 16'b0000000000000000;
	sram_mem[121050] = 16'b0000000000000000;
	sram_mem[121051] = 16'b0000000000000000;
	sram_mem[121052] = 16'b0000000000000000;
	sram_mem[121053] = 16'b0000000000000000;
	sram_mem[121054] = 16'b0000000000000000;
	sram_mem[121055] = 16'b0000000000000000;
	sram_mem[121056] = 16'b0000000000000000;
	sram_mem[121057] = 16'b0000000000000000;
	sram_mem[121058] = 16'b0000000000000000;
	sram_mem[121059] = 16'b0000000000000000;
	sram_mem[121060] = 16'b0000000000000000;
	sram_mem[121061] = 16'b0000000000000000;
	sram_mem[121062] = 16'b0000000000000000;
	sram_mem[121063] = 16'b0000000000000000;
	sram_mem[121064] = 16'b0000000000000000;
	sram_mem[121065] = 16'b0000000000000000;
	sram_mem[121066] = 16'b0000000000000000;
	sram_mem[121067] = 16'b0000000000000000;
	sram_mem[121068] = 16'b0000000000000000;
	sram_mem[121069] = 16'b0000000000000000;
	sram_mem[121070] = 16'b0000000000000000;
	sram_mem[121071] = 16'b0000000000000000;
	sram_mem[121072] = 16'b0000000000000000;
	sram_mem[121073] = 16'b0000000000000000;
	sram_mem[121074] = 16'b0000000000000000;
	sram_mem[121075] = 16'b0000000000000000;
	sram_mem[121076] = 16'b0000000000000000;
	sram_mem[121077] = 16'b0000000000000000;
	sram_mem[121078] = 16'b0000000000000000;
	sram_mem[121079] = 16'b0000000000000000;
	sram_mem[121080] = 16'b0000000000000000;
	sram_mem[121081] = 16'b0000000000000000;
	sram_mem[121082] = 16'b0000000000000000;
	sram_mem[121083] = 16'b0000000000000000;
	sram_mem[121084] = 16'b0000000000000000;
	sram_mem[121085] = 16'b0000000000000000;
	sram_mem[121086] = 16'b0000000000000000;
	sram_mem[121087] = 16'b0000000000000000;
	sram_mem[121088] = 16'b0000000000000000;
	sram_mem[121089] = 16'b0000000000000000;
	sram_mem[121090] = 16'b0000000000000000;
	sram_mem[121091] = 16'b0000000000000000;
	sram_mem[121092] = 16'b0000000000000000;
	sram_mem[121093] = 16'b0000000000000000;
	sram_mem[121094] = 16'b0000000000000000;
	sram_mem[121095] = 16'b0000000000000000;
	sram_mem[121096] = 16'b0000000000000000;
	sram_mem[121097] = 16'b0000000000000000;
	sram_mem[121098] = 16'b0000000000000000;
	sram_mem[121099] = 16'b0000000000000000;
	sram_mem[121100] = 16'b0000000000000000;
	sram_mem[121101] = 16'b0000000000000000;
	sram_mem[121102] = 16'b0000000000000000;
	sram_mem[121103] = 16'b0000000000000000;
	sram_mem[121104] = 16'b0000000000000000;
	sram_mem[121105] = 16'b0000000000000000;
	sram_mem[121106] = 16'b0000000000000000;
	sram_mem[121107] = 16'b0000000000000000;
	sram_mem[121108] = 16'b0000000000000000;
	sram_mem[121109] = 16'b0000000000000000;
	sram_mem[121110] = 16'b0000000000000000;
	sram_mem[121111] = 16'b0000000000000000;
	sram_mem[121112] = 16'b0000000000000000;
	sram_mem[121113] = 16'b0000000000000000;
	sram_mem[121114] = 16'b0000000000000000;
	sram_mem[121115] = 16'b0000000000000000;
	sram_mem[121116] = 16'b0000000000000000;
	sram_mem[121117] = 16'b0000000000000000;
	sram_mem[121118] = 16'b0000000000000000;
	sram_mem[121119] = 16'b0000000000000000;
	sram_mem[121120] = 16'b0000000000000000;
	sram_mem[121121] = 16'b0000000000000000;
	sram_mem[121122] = 16'b0000000000000000;
	sram_mem[121123] = 16'b0000000000000000;
	sram_mem[121124] = 16'b0000000000000000;
	sram_mem[121125] = 16'b0000000000000000;
	sram_mem[121126] = 16'b0000000000000000;
	sram_mem[121127] = 16'b0000000000000000;
	sram_mem[121128] = 16'b0000000000000000;
	sram_mem[121129] = 16'b0000000000000000;
	sram_mem[121130] = 16'b0000000000000000;
	sram_mem[121131] = 16'b0000000000000000;
	sram_mem[121132] = 16'b0000000000000000;
	sram_mem[121133] = 16'b0000000000000000;
	sram_mem[121134] = 16'b0000000000000000;
	sram_mem[121135] = 16'b0000000000000000;
	sram_mem[121136] = 16'b0000000000000000;
	sram_mem[121137] = 16'b0000000000000000;
	sram_mem[121138] = 16'b0000000000000000;
	sram_mem[121139] = 16'b0000000000000000;
	sram_mem[121140] = 16'b0000000000000000;
	sram_mem[121141] = 16'b0000000000000000;
	sram_mem[121142] = 16'b0000000000000000;
	sram_mem[121143] = 16'b0000000000000000;
	sram_mem[121144] = 16'b0000000000000000;
	sram_mem[121145] = 16'b0000000000000000;
	sram_mem[121146] = 16'b0000000000000000;
	sram_mem[121147] = 16'b0000000000000000;
	sram_mem[121148] = 16'b0000000000000000;
	sram_mem[121149] = 16'b0000000000000000;
	sram_mem[121150] = 16'b0000000000000000;
	sram_mem[121151] = 16'b0000000000000000;
	sram_mem[121152] = 16'b0000000000000000;
	sram_mem[121153] = 16'b0000000000000000;
	sram_mem[121154] = 16'b0000000000000000;
	sram_mem[121155] = 16'b0000000000000000;
	sram_mem[121156] = 16'b0000000000000000;
	sram_mem[121157] = 16'b0000000000000000;
	sram_mem[121158] = 16'b0000000000000000;
	sram_mem[121159] = 16'b0000000000000000;
	sram_mem[121160] = 16'b0000000000000000;
	sram_mem[121161] = 16'b0000000000000000;
	sram_mem[121162] = 16'b0000000000000000;
	sram_mem[121163] = 16'b0000000000000000;
	sram_mem[121164] = 16'b0000000000000000;
	sram_mem[121165] = 16'b0000000000000000;
	sram_mem[121166] = 16'b0000000000000000;
	sram_mem[121167] = 16'b0000000000000000;
	sram_mem[121168] = 16'b0000000000000000;
	sram_mem[121169] = 16'b0000000000000000;
	sram_mem[121170] = 16'b0000000000000000;
	sram_mem[121171] = 16'b0000000000000000;
	sram_mem[121172] = 16'b0000000000000000;
	sram_mem[121173] = 16'b0000000000000000;
	sram_mem[121174] = 16'b0000000000000000;
	sram_mem[121175] = 16'b0000000000000000;
	sram_mem[121176] = 16'b0000000000000000;
	sram_mem[121177] = 16'b0000000000000000;
	sram_mem[121178] = 16'b0000000000000000;
	sram_mem[121179] = 16'b0000000000000000;
	sram_mem[121180] = 16'b0000000000000000;
	sram_mem[121181] = 16'b0000000000000000;
	sram_mem[121182] = 16'b0000000000000000;
	sram_mem[121183] = 16'b0000000000000000;
	sram_mem[121184] = 16'b0000000000000000;
	sram_mem[121185] = 16'b0000000000000000;
	sram_mem[121186] = 16'b0000000000000000;
	sram_mem[121187] = 16'b0000000000000000;
	sram_mem[121188] = 16'b0000000000000000;
	sram_mem[121189] = 16'b0000000000000000;
	sram_mem[121190] = 16'b0000000000000000;
	sram_mem[121191] = 16'b0000000000000000;
	sram_mem[121192] = 16'b0000000000000000;
	sram_mem[121193] = 16'b0000000000000000;
	sram_mem[121194] = 16'b0000000000000000;
	sram_mem[121195] = 16'b0000000000000000;
	sram_mem[121196] = 16'b0000000000000000;
	sram_mem[121197] = 16'b0000000000000000;
	sram_mem[121198] = 16'b0000000000000000;
	sram_mem[121199] = 16'b0000000000000000;
	sram_mem[121200] = 16'b0000000000000000;
	sram_mem[121201] = 16'b0000000000000000;
	sram_mem[121202] = 16'b0000000000000000;
	sram_mem[121203] = 16'b0000000000000000;
	sram_mem[121204] = 16'b0000000000000000;
	sram_mem[121205] = 16'b0000000000000000;
	sram_mem[121206] = 16'b0000000000000000;
	sram_mem[121207] = 16'b0000000000000000;
	sram_mem[121208] = 16'b0000000000000000;
	sram_mem[121209] = 16'b0000000000000000;
	sram_mem[121210] = 16'b0000000000000000;
	sram_mem[121211] = 16'b0000000000000000;
	sram_mem[121212] = 16'b0000000000000000;
	sram_mem[121213] = 16'b0000000000000000;
	sram_mem[121214] = 16'b0000000000000000;
	sram_mem[121215] = 16'b0000000000000000;
	sram_mem[121216] = 16'b0000000000000000;
	sram_mem[121217] = 16'b0000000000000000;
	sram_mem[121218] = 16'b0000000000000000;
	sram_mem[121219] = 16'b0000000000000000;
	sram_mem[121220] = 16'b0000000000000000;
	sram_mem[121221] = 16'b0000000000000000;
	sram_mem[121222] = 16'b0000000000000000;
	sram_mem[121223] = 16'b0000000000000000;
	sram_mem[121224] = 16'b0000000000000000;
	sram_mem[121225] = 16'b0000000000000000;
	sram_mem[121226] = 16'b0000000000000000;
	sram_mem[121227] = 16'b0000000000000000;
	sram_mem[121228] = 16'b0000000000000000;
	sram_mem[121229] = 16'b0000000000000000;
	sram_mem[121230] = 16'b0000000000000000;
	sram_mem[121231] = 16'b0000000000000000;
	sram_mem[121232] = 16'b0000000000000000;
	sram_mem[121233] = 16'b0000000000000000;
	sram_mem[121234] = 16'b0000000000000000;
	sram_mem[121235] = 16'b0000000000000000;
	sram_mem[121236] = 16'b0000000000000000;
	sram_mem[121237] = 16'b0000000000000000;
	sram_mem[121238] = 16'b0000000000000000;
	sram_mem[121239] = 16'b0000000000000000;
	sram_mem[121240] = 16'b0000000000000000;
	sram_mem[121241] = 16'b0000000000000000;
	sram_mem[121242] = 16'b0000000000000000;
	sram_mem[121243] = 16'b0000000000000000;
	sram_mem[121244] = 16'b0000000000000000;
	sram_mem[121245] = 16'b0000000000000000;
	sram_mem[121246] = 16'b0000000000000000;
	sram_mem[121247] = 16'b0000000000000000;
	sram_mem[121248] = 16'b0000000000000000;
	sram_mem[121249] = 16'b0000000000000000;
	sram_mem[121250] = 16'b0000000000000000;
	sram_mem[121251] = 16'b0000000000000000;
	sram_mem[121252] = 16'b0000000000000000;
	sram_mem[121253] = 16'b0000000000000000;
	sram_mem[121254] = 16'b0000000000000000;
	sram_mem[121255] = 16'b0000000000000000;
	sram_mem[121256] = 16'b0000000000000000;
	sram_mem[121257] = 16'b0000000000000000;
	sram_mem[121258] = 16'b0000000000000000;
	sram_mem[121259] = 16'b0000000000000000;
	sram_mem[121260] = 16'b0000000000000000;
	sram_mem[121261] = 16'b0000000000000000;
	sram_mem[121262] = 16'b0000000000000000;
	sram_mem[121263] = 16'b0000000000000000;
	sram_mem[121264] = 16'b0000000000000000;
	sram_mem[121265] = 16'b0000000000000000;
	sram_mem[121266] = 16'b0000000000000000;
	sram_mem[121267] = 16'b0000000000000000;
	sram_mem[121268] = 16'b0000000000000000;
	sram_mem[121269] = 16'b0000000000000000;
	sram_mem[121270] = 16'b0000000000000000;
	sram_mem[121271] = 16'b0000000000000000;
	sram_mem[121272] = 16'b0000000000000000;
	sram_mem[121273] = 16'b0000000000000000;
	sram_mem[121274] = 16'b0000000000000000;
	sram_mem[121275] = 16'b0000000000000000;
	sram_mem[121276] = 16'b0000000000000000;
	sram_mem[121277] = 16'b0000000000000000;
	sram_mem[121278] = 16'b0000000000000000;
	sram_mem[121279] = 16'b0000000000000000;
	sram_mem[121280] = 16'b0000000000000000;
	sram_mem[121281] = 16'b0000000000000000;
	sram_mem[121282] = 16'b0000000000000000;
	sram_mem[121283] = 16'b0000000000000000;
	sram_mem[121284] = 16'b0000000000000000;
	sram_mem[121285] = 16'b0000000000000000;
	sram_mem[121286] = 16'b0000000000000000;
	sram_mem[121287] = 16'b0000000000000000;
	sram_mem[121288] = 16'b0000000000000000;
	sram_mem[121289] = 16'b0000000000000000;
	sram_mem[121290] = 16'b0000000000000000;
	sram_mem[121291] = 16'b0000000000000000;
	sram_mem[121292] = 16'b0000000000000000;
	sram_mem[121293] = 16'b0000000000000000;
	sram_mem[121294] = 16'b0000000000000000;
	sram_mem[121295] = 16'b0000000000000000;
	sram_mem[121296] = 16'b0000000000000000;
	sram_mem[121297] = 16'b0000000000000000;
	sram_mem[121298] = 16'b0000000000000000;
	sram_mem[121299] = 16'b0000000000000000;
	sram_mem[121300] = 16'b0000000000000000;
	sram_mem[121301] = 16'b0000000000000000;
	sram_mem[121302] = 16'b0000000000000000;
	sram_mem[121303] = 16'b0000000000000000;
	sram_mem[121304] = 16'b0000000000000000;
	sram_mem[121305] = 16'b0000000000000000;
	sram_mem[121306] = 16'b0000000000000000;
	sram_mem[121307] = 16'b0000000000000000;
	sram_mem[121308] = 16'b0000000000000000;
	sram_mem[121309] = 16'b0000000000000000;
	sram_mem[121310] = 16'b0000000000000000;
	sram_mem[121311] = 16'b0000000000000000;
	sram_mem[121312] = 16'b0000000000000000;
	sram_mem[121313] = 16'b0000000000000000;
	sram_mem[121314] = 16'b0000000000000000;
	sram_mem[121315] = 16'b0000000000000000;
	sram_mem[121316] = 16'b0000000000000000;
	sram_mem[121317] = 16'b0000000000000000;
	sram_mem[121318] = 16'b0000000000000000;
	sram_mem[121319] = 16'b0000000000000000;
	sram_mem[121320] = 16'b0000000000000000;
	sram_mem[121321] = 16'b0000000000000000;
	sram_mem[121322] = 16'b0000000000000000;
	sram_mem[121323] = 16'b0000000000000000;
	sram_mem[121324] = 16'b0000000000000000;
	sram_mem[121325] = 16'b0000000000000000;
	sram_mem[121326] = 16'b0000000000000000;
	sram_mem[121327] = 16'b0000000000000000;
	sram_mem[121328] = 16'b0000000000000000;
	sram_mem[121329] = 16'b0000000000000000;
	sram_mem[121330] = 16'b0000000000000000;
	sram_mem[121331] = 16'b0000000000000000;
	sram_mem[121332] = 16'b0000000000000000;
	sram_mem[121333] = 16'b0000000000000000;
	sram_mem[121334] = 16'b0000000000000000;
	sram_mem[121335] = 16'b0000000000000000;
	sram_mem[121336] = 16'b0000000000000000;
	sram_mem[121337] = 16'b0000000000000000;
	sram_mem[121338] = 16'b0000000000000000;
	sram_mem[121339] = 16'b0000000000000000;
	sram_mem[121340] = 16'b0000000000000000;
	sram_mem[121341] = 16'b0000000000000000;
	sram_mem[121342] = 16'b0000000000000000;
	sram_mem[121343] = 16'b0000000000000000;
	sram_mem[121344] = 16'b0000000000000000;
	sram_mem[121345] = 16'b0000000000000000;
	sram_mem[121346] = 16'b0000000000000000;
	sram_mem[121347] = 16'b0000000000000000;
	sram_mem[121348] = 16'b0000000000000000;
	sram_mem[121349] = 16'b0000000000000000;
	sram_mem[121350] = 16'b0000000000000000;
	sram_mem[121351] = 16'b0000000000000000;
	sram_mem[121352] = 16'b0000000000000000;
	sram_mem[121353] = 16'b0000000000000000;
	sram_mem[121354] = 16'b0000000000000000;
	sram_mem[121355] = 16'b0000000000000000;
	sram_mem[121356] = 16'b0000000000000000;
	sram_mem[121357] = 16'b0000000000000000;
	sram_mem[121358] = 16'b0000000000000000;
	sram_mem[121359] = 16'b0000000000000000;
	sram_mem[121360] = 16'b0000000000000000;
	sram_mem[121361] = 16'b0000000000000000;
	sram_mem[121362] = 16'b0000000000000000;
	sram_mem[121363] = 16'b0000000000000000;
	sram_mem[121364] = 16'b0000000000000000;
	sram_mem[121365] = 16'b0000000000000000;
	sram_mem[121366] = 16'b0000000000000000;
	sram_mem[121367] = 16'b0000000000000000;
	sram_mem[121368] = 16'b0000000000000000;
	sram_mem[121369] = 16'b0000000000000000;
	sram_mem[121370] = 16'b0000000000000000;
	sram_mem[121371] = 16'b0000000000000000;
	sram_mem[121372] = 16'b0000000000000000;
	sram_mem[121373] = 16'b0000000000000000;
	sram_mem[121374] = 16'b0000000000000000;
	sram_mem[121375] = 16'b0000000000000000;
	sram_mem[121376] = 16'b0000000000000000;
	sram_mem[121377] = 16'b0000000000000000;
	sram_mem[121378] = 16'b0000000000000000;
	sram_mem[121379] = 16'b0000000000000000;
	sram_mem[121380] = 16'b0000000000000000;
	sram_mem[121381] = 16'b0000000000000000;
	sram_mem[121382] = 16'b0000000000000000;
	sram_mem[121383] = 16'b0000000000000000;
	sram_mem[121384] = 16'b0000000000000000;
	sram_mem[121385] = 16'b0000000000000000;
	sram_mem[121386] = 16'b0000000000000000;
	sram_mem[121387] = 16'b0000000000000000;
	sram_mem[121388] = 16'b0000000000000000;
	sram_mem[121389] = 16'b0000000000000000;
	sram_mem[121390] = 16'b0000000000000000;
	sram_mem[121391] = 16'b0000000000000000;
	sram_mem[121392] = 16'b0000000000000000;
	sram_mem[121393] = 16'b0000000000000000;
	sram_mem[121394] = 16'b0000000000000000;
	sram_mem[121395] = 16'b0000000000000000;
	sram_mem[121396] = 16'b0000000000000000;
	sram_mem[121397] = 16'b0000000000000000;
	sram_mem[121398] = 16'b0000000000000000;
	sram_mem[121399] = 16'b0000000000000000;
	sram_mem[121400] = 16'b0000000000000000;
	sram_mem[121401] = 16'b0000000000000000;
	sram_mem[121402] = 16'b0000000000000000;
	sram_mem[121403] = 16'b0000000000000000;
	sram_mem[121404] = 16'b0000000000000000;
	sram_mem[121405] = 16'b0000000000000000;
	sram_mem[121406] = 16'b0000000000000000;
	sram_mem[121407] = 16'b0000000000000000;
	sram_mem[121408] = 16'b0000000000000000;
	sram_mem[121409] = 16'b0000000000000000;
	sram_mem[121410] = 16'b0000000000000000;
	sram_mem[121411] = 16'b0000000000000000;
	sram_mem[121412] = 16'b0000000000000000;
	sram_mem[121413] = 16'b0000000000000000;
	sram_mem[121414] = 16'b0000000000000000;
	sram_mem[121415] = 16'b0000000000000000;
	sram_mem[121416] = 16'b0000000000000000;
	sram_mem[121417] = 16'b0000000000000000;
	sram_mem[121418] = 16'b0000000000000000;
	sram_mem[121419] = 16'b0000000000000000;
	sram_mem[121420] = 16'b0000000000000000;
	sram_mem[121421] = 16'b0000000000000000;
	sram_mem[121422] = 16'b0000000000000000;
	sram_mem[121423] = 16'b0000000000000000;
	sram_mem[121424] = 16'b0000000000000000;
	sram_mem[121425] = 16'b0000000000000000;
	sram_mem[121426] = 16'b0000000000000000;
	sram_mem[121427] = 16'b0000000000000000;
	sram_mem[121428] = 16'b0000000000000000;
	sram_mem[121429] = 16'b0000000000000000;
	sram_mem[121430] = 16'b0000000000000000;
	sram_mem[121431] = 16'b0000000000000000;
	sram_mem[121432] = 16'b0000000000000000;
	sram_mem[121433] = 16'b0000000000000000;
	sram_mem[121434] = 16'b0000000000000000;
	sram_mem[121435] = 16'b0000000000000000;
	sram_mem[121436] = 16'b0000000000000000;
	sram_mem[121437] = 16'b0000000000000000;
	sram_mem[121438] = 16'b0000000000000000;
	sram_mem[121439] = 16'b0000000000000000;
	sram_mem[121440] = 16'b0000000000000000;
	sram_mem[121441] = 16'b0000000000000000;
	sram_mem[121442] = 16'b0000000000000000;
	sram_mem[121443] = 16'b0000000000000000;
	sram_mem[121444] = 16'b0000000000000000;
	sram_mem[121445] = 16'b0000000000000000;
	sram_mem[121446] = 16'b0000000000000000;
	sram_mem[121447] = 16'b0000000000000000;
	sram_mem[121448] = 16'b0000000000000000;
	sram_mem[121449] = 16'b0000000000000000;
	sram_mem[121450] = 16'b0000000000000000;
	sram_mem[121451] = 16'b0000000000000000;
	sram_mem[121452] = 16'b0000000000000000;
	sram_mem[121453] = 16'b0000000000000000;
	sram_mem[121454] = 16'b0000000000000000;
	sram_mem[121455] = 16'b0000000000000000;
	sram_mem[121456] = 16'b0000000000000000;
	sram_mem[121457] = 16'b0000000000000000;
	sram_mem[121458] = 16'b0000000000000000;
	sram_mem[121459] = 16'b0000000000000000;
	sram_mem[121460] = 16'b0000000000000000;
	sram_mem[121461] = 16'b0000000000000000;
	sram_mem[121462] = 16'b0000000000000000;
	sram_mem[121463] = 16'b0000000000000000;
	sram_mem[121464] = 16'b0000000000000000;
	sram_mem[121465] = 16'b0000000000000000;
	sram_mem[121466] = 16'b0000000000000000;
	sram_mem[121467] = 16'b0000000000000000;
	sram_mem[121468] = 16'b0000000000000000;
	sram_mem[121469] = 16'b0000000000000000;
	sram_mem[121470] = 16'b0000000000000000;
	sram_mem[121471] = 16'b0000000000000000;
	sram_mem[121472] = 16'b0000000000000000;
	sram_mem[121473] = 16'b0000000000000000;
	sram_mem[121474] = 16'b0000000000000000;
	sram_mem[121475] = 16'b0000000000000000;
	sram_mem[121476] = 16'b0000000000000000;
	sram_mem[121477] = 16'b0000000000000000;
	sram_mem[121478] = 16'b0000000000000000;
	sram_mem[121479] = 16'b0000000000000000;
	sram_mem[121480] = 16'b0000000000000000;
	sram_mem[121481] = 16'b0000000000000000;
	sram_mem[121482] = 16'b0000000000000000;
	sram_mem[121483] = 16'b0000000000000000;
	sram_mem[121484] = 16'b0000000000000000;
	sram_mem[121485] = 16'b0000000000000000;
	sram_mem[121486] = 16'b0000000000000000;
	sram_mem[121487] = 16'b0000000000000000;
	sram_mem[121488] = 16'b0000000000000000;
	sram_mem[121489] = 16'b0000000000000000;
	sram_mem[121490] = 16'b0000000000000000;
	sram_mem[121491] = 16'b0000000000000000;
	sram_mem[121492] = 16'b0000000000000000;
	sram_mem[121493] = 16'b0000000000000000;
	sram_mem[121494] = 16'b0000000000000000;
	sram_mem[121495] = 16'b0000000000000000;
	sram_mem[121496] = 16'b0000000000000000;
	sram_mem[121497] = 16'b0000000000000000;
	sram_mem[121498] = 16'b0000000000000000;
	sram_mem[121499] = 16'b0000000000000000;
	sram_mem[121500] = 16'b0000000000000000;
	sram_mem[121501] = 16'b0000000000000000;
	sram_mem[121502] = 16'b0000000000000000;
	sram_mem[121503] = 16'b0000000000000000;
	sram_mem[121504] = 16'b0000000000000000;
	sram_mem[121505] = 16'b0000000000000000;
	sram_mem[121506] = 16'b0000000000000000;
	sram_mem[121507] = 16'b0000000000000000;
	sram_mem[121508] = 16'b0000000000000000;
	sram_mem[121509] = 16'b0000000000000000;
	sram_mem[121510] = 16'b0000000000000000;
	sram_mem[121511] = 16'b0000000000000000;
	sram_mem[121512] = 16'b0000000000000000;
	sram_mem[121513] = 16'b0000000000000000;
	sram_mem[121514] = 16'b0000000000000000;
	sram_mem[121515] = 16'b0000000000000000;
	sram_mem[121516] = 16'b0000000000000000;
	sram_mem[121517] = 16'b0000000000000000;
	sram_mem[121518] = 16'b0000000000000000;
	sram_mem[121519] = 16'b0000000000000000;
	sram_mem[121520] = 16'b0000000000000000;
	sram_mem[121521] = 16'b0000000000000000;
	sram_mem[121522] = 16'b0000000000000000;
	sram_mem[121523] = 16'b0000000000000000;
	sram_mem[121524] = 16'b0000000000000000;
	sram_mem[121525] = 16'b0000000000000000;
	sram_mem[121526] = 16'b0000000000000000;
	sram_mem[121527] = 16'b0000000000000000;
	sram_mem[121528] = 16'b0000000000000000;
	sram_mem[121529] = 16'b0000000000000000;
	sram_mem[121530] = 16'b0000000000000000;
	sram_mem[121531] = 16'b0000000000000000;
	sram_mem[121532] = 16'b0000000000000000;
	sram_mem[121533] = 16'b0000000000000000;
	sram_mem[121534] = 16'b0000000000000000;
	sram_mem[121535] = 16'b0000000000000000;
	sram_mem[121536] = 16'b0000000000000000;
	sram_mem[121537] = 16'b0000000000000000;
	sram_mem[121538] = 16'b0000000000000000;
	sram_mem[121539] = 16'b0000000000000000;
	sram_mem[121540] = 16'b0000000000000000;
	sram_mem[121541] = 16'b0000000000000000;
	sram_mem[121542] = 16'b0000000000000000;
	sram_mem[121543] = 16'b0000000000000000;
	sram_mem[121544] = 16'b0000000000000000;
	sram_mem[121545] = 16'b0000000000000000;
	sram_mem[121546] = 16'b0000000000000000;
	sram_mem[121547] = 16'b0000000000000000;
	sram_mem[121548] = 16'b0000000000000000;
	sram_mem[121549] = 16'b0000000000000000;
	sram_mem[121550] = 16'b0000000000000000;
	sram_mem[121551] = 16'b0000000000000000;
	sram_mem[121552] = 16'b0000000000000000;
	sram_mem[121553] = 16'b0000000000000000;
	sram_mem[121554] = 16'b0000000000000000;
	sram_mem[121555] = 16'b0000000000000000;
	sram_mem[121556] = 16'b0000000000000000;
	sram_mem[121557] = 16'b0000000000000000;
	sram_mem[121558] = 16'b0000000000000000;
	sram_mem[121559] = 16'b0000000000000000;
	sram_mem[121560] = 16'b0000000000000000;
	sram_mem[121561] = 16'b0000000000000000;
	sram_mem[121562] = 16'b0000000000000000;
	sram_mem[121563] = 16'b0000000000000000;
	sram_mem[121564] = 16'b0000000000000000;
	sram_mem[121565] = 16'b0000000000000000;
	sram_mem[121566] = 16'b0000000000000000;
	sram_mem[121567] = 16'b0000000000000000;
	sram_mem[121568] = 16'b0000000000000000;
	sram_mem[121569] = 16'b0000000000000000;
	sram_mem[121570] = 16'b0000000000000000;
	sram_mem[121571] = 16'b0000000000000000;
	sram_mem[121572] = 16'b0000000000000000;
	sram_mem[121573] = 16'b0000000000000000;
	sram_mem[121574] = 16'b0000000000000000;
	sram_mem[121575] = 16'b0000000000000000;
	sram_mem[121576] = 16'b0000000000000000;
	sram_mem[121577] = 16'b0000000000000000;
	sram_mem[121578] = 16'b0000000000000000;
	sram_mem[121579] = 16'b0000000000000000;
	sram_mem[121580] = 16'b0000000000000000;
	sram_mem[121581] = 16'b0000000000000000;
	sram_mem[121582] = 16'b0000000000000000;
	sram_mem[121583] = 16'b0000000000000000;
	sram_mem[121584] = 16'b0000000000000000;
	sram_mem[121585] = 16'b0000000000000000;
	sram_mem[121586] = 16'b0000000000000000;
	sram_mem[121587] = 16'b0000000000000000;
	sram_mem[121588] = 16'b0000000000000000;
	sram_mem[121589] = 16'b0000000000000000;
	sram_mem[121590] = 16'b0000000000000000;
	sram_mem[121591] = 16'b0000000000000000;
	sram_mem[121592] = 16'b0000000000000000;
	sram_mem[121593] = 16'b0000000000000000;
	sram_mem[121594] = 16'b0000000000000000;
	sram_mem[121595] = 16'b0000000000000000;
	sram_mem[121596] = 16'b0000000000000000;
	sram_mem[121597] = 16'b0000000000000000;
	sram_mem[121598] = 16'b0000000000000000;
	sram_mem[121599] = 16'b0000000000000000;
	sram_mem[121600] = 16'b0000000000000000;
	sram_mem[121601] = 16'b0000000000000000;
	sram_mem[121602] = 16'b0000000000000000;
	sram_mem[121603] = 16'b0000000000000000;
	sram_mem[121604] = 16'b0000000000000000;
	sram_mem[121605] = 16'b0000000000000000;
	sram_mem[121606] = 16'b0000000000000000;
	sram_mem[121607] = 16'b0000000000000000;
	sram_mem[121608] = 16'b0000000000000000;
	sram_mem[121609] = 16'b0000000000000000;
	sram_mem[121610] = 16'b0000000000000000;
	sram_mem[121611] = 16'b0000000000000000;
	sram_mem[121612] = 16'b0000000000000000;
	sram_mem[121613] = 16'b0000000000000000;
	sram_mem[121614] = 16'b0000000000000000;
	sram_mem[121615] = 16'b0000000000000000;
	sram_mem[121616] = 16'b0000000000000000;
	sram_mem[121617] = 16'b0000000000000000;
	sram_mem[121618] = 16'b0000000000000000;
	sram_mem[121619] = 16'b0000000000000000;
	sram_mem[121620] = 16'b0000000000000000;
	sram_mem[121621] = 16'b0000000000000000;
	sram_mem[121622] = 16'b0000000000000000;
	sram_mem[121623] = 16'b0000000000000000;
	sram_mem[121624] = 16'b0000000000000000;
	sram_mem[121625] = 16'b0000000000000000;
	sram_mem[121626] = 16'b0000000000000000;
	sram_mem[121627] = 16'b0000000000000000;
	sram_mem[121628] = 16'b0000000000000000;
	sram_mem[121629] = 16'b0000000000000000;
	sram_mem[121630] = 16'b0000000000000000;
	sram_mem[121631] = 16'b0000000000000000;
	sram_mem[121632] = 16'b0000000000000000;
	sram_mem[121633] = 16'b0000000000000000;
	sram_mem[121634] = 16'b0000000000000000;
	sram_mem[121635] = 16'b0000000000000000;
	sram_mem[121636] = 16'b0000000000000000;
	sram_mem[121637] = 16'b0000000000000000;
	sram_mem[121638] = 16'b0000000000000000;
	sram_mem[121639] = 16'b0000000000000000;
	sram_mem[121640] = 16'b0000000000000000;
	sram_mem[121641] = 16'b0000000000000000;
	sram_mem[121642] = 16'b0000000000000000;
	sram_mem[121643] = 16'b0000000000000000;
	sram_mem[121644] = 16'b0000000000000000;
	sram_mem[121645] = 16'b0000000000000000;
	sram_mem[121646] = 16'b0000000000000000;
	sram_mem[121647] = 16'b0000000000000000;
	sram_mem[121648] = 16'b0000000000000000;
	sram_mem[121649] = 16'b0000000000000000;
	sram_mem[121650] = 16'b0000000000000000;
	sram_mem[121651] = 16'b0000000000000000;
	sram_mem[121652] = 16'b0000000000000000;
	sram_mem[121653] = 16'b0000000000000000;
	sram_mem[121654] = 16'b0000000000000000;
	sram_mem[121655] = 16'b0000000000000000;
	sram_mem[121656] = 16'b0000000000000000;
	sram_mem[121657] = 16'b0000000000000000;
	sram_mem[121658] = 16'b0000000000000000;
	sram_mem[121659] = 16'b0000000000000000;
	sram_mem[121660] = 16'b0000000000000000;
	sram_mem[121661] = 16'b0000000000000000;
	sram_mem[121662] = 16'b0000000000000000;
	sram_mem[121663] = 16'b0000000000000000;
	sram_mem[121664] = 16'b0000000000000000;
	sram_mem[121665] = 16'b0000000000000000;
	sram_mem[121666] = 16'b0000000000000000;
	sram_mem[121667] = 16'b0000000000000000;
	sram_mem[121668] = 16'b0000000000000000;
	sram_mem[121669] = 16'b0000000000000000;
	sram_mem[121670] = 16'b0000000000000000;
	sram_mem[121671] = 16'b0000000000000000;
	sram_mem[121672] = 16'b0000000000000000;
	sram_mem[121673] = 16'b0000000000000000;
	sram_mem[121674] = 16'b0000000000000000;
	sram_mem[121675] = 16'b0000000000000000;
	sram_mem[121676] = 16'b0000000000000000;
	sram_mem[121677] = 16'b0000000000000000;
	sram_mem[121678] = 16'b0000000000000000;
	sram_mem[121679] = 16'b0000000000000000;
	sram_mem[121680] = 16'b0000000000000000;
	sram_mem[121681] = 16'b0000000000000000;
	sram_mem[121682] = 16'b0000000000000000;
	sram_mem[121683] = 16'b0000000000000000;
	sram_mem[121684] = 16'b0000000000000000;
	sram_mem[121685] = 16'b0000000000000000;
	sram_mem[121686] = 16'b0000000000000000;
	sram_mem[121687] = 16'b0000000000000000;
	sram_mem[121688] = 16'b0000000000000000;
	sram_mem[121689] = 16'b0000000000000000;
	sram_mem[121690] = 16'b0000000000000000;
	sram_mem[121691] = 16'b0000000000000000;
	sram_mem[121692] = 16'b0000000000000000;
	sram_mem[121693] = 16'b0000000000000000;
	sram_mem[121694] = 16'b0000000000000000;
	sram_mem[121695] = 16'b0000000000000000;
	sram_mem[121696] = 16'b0000000000000000;
	sram_mem[121697] = 16'b0000000000000000;
	sram_mem[121698] = 16'b0000000000000000;
	sram_mem[121699] = 16'b0000000000000000;
	sram_mem[121700] = 16'b0000000000000000;
	sram_mem[121701] = 16'b0000000000000000;
	sram_mem[121702] = 16'b0000000000000000;
	sram_mem[121703] = 16'b0000000000000000;
	sram_mem[121704] = 16'b0000000000000000;
	sram_mem[121705] = 16'b0000000000000000;
	sram_mem[121706] = 16'b0000000000000000;
	sram_mem[121707] = 16'b0000000000000000;
	sram_mem[121708] = 16'b0000000000000000;
	sram_mem[121709] = 16'b0000000000000000;
	sram_mem[121710] = 16'b0000000000000000;
	sram_mem[121711] = 16'b0000000000000000;
	sram_mem[121712] = 16'b0000000000000000;
	sram_mem[121713] = 16'b0000000000000000;
	sram_mem[121714] = 16'b0000000000000000;
	sram_mem[121715] = 16'b0000000000000000;
	sram_mem[121716] = 16'b0000000000000000;
	sram_mem[121717] = 16'b0000000000000000;
	sram_mem[121718] = 16'b0000000000000000;
	sram_mem[121719] = 16'b0000000000000000;
	sram_mem[121720] = 16'b0000000000000000;
	sram_mem[121721] = 16'b0000000000000000;
	sram_mem[121722] = 16'b0000000000000000;
	sram_mem[121723] = 16'b0000000000000000;
	sram_mem[121724] = 16'b0000000000000000;
	sram_mem[121725] = 16'b0000000000000000;
	sram_mem[121726] = 16'b0000000000000000;
	sram_mem[121727] = 16'b0000000000000000;
	sram_mem[121728] = 16'b0000000000000000;
	sram_mem[121729] = 16'b0000000000000000;
	sram_mem[121730] = 16'b0000000000000000;
	sram_mem[121731] = 16'b0000000000000000;
	sram_mem[121732] = 16'b0000000000000000;
	sram_mem[121733] = 16'b0000000000000000;
	sram_mem[121734] = 16'b0000000000000000;
	sram_mem[121735] = 16'b0000000000000000;
	sram_mem[121736] = 16'b0000000000000000;
	sram_mem[121737] = 16'b0000000000000000;
	sram_mem[121738] = 16'b0000000000000000;
	sram_mem[121739] = 16'b0000000000000000;
	sram_mem[121740] = 16'b0000000000000000;
	sram_mem[121741] = 16'b0000000000000000;
	sram_mem[121742] = 16'b0000000000000000;
	sram_mem[121743] = 16'b0000000000000000;
	sram_mem[121744] = 16'b0000000000000000;
	sram_mem[121745] = 16'b0000000000000000;
	sram_mem[121746] = 16'b0000000000000000;
	sram_mem[121747] = 16'b0000000000000000;
	sram_mem[121748] = 16'b0000000000000000;
	sram_mem[121749] = 16'b0000000000000000;
	sram_mem[121750] = 16'b0000000000000000;
	sram_mem[121751] = 16'b0000000000000000;
	sram_mem[121752] = 16'b0000000000000000;
	sram_mem[121753] = 16'b0000000000000000;
	sram_mem[121754] = 16'b0000000000000000;
	sram_mem[121755] = 16'b0000000000000000;
	sram_mem[121756] = 16'b0000000000000000;
	sram_mem[121757] = 16'b0000000000000000;
	sram_mem[121758] = 16'b0000000000000000;
	sram_mem[121759] = 16'b0000000000000000;
	sram_mem[121760] = 16'b0000000000000000;
	sram_mem[121761] = 16'b0000000000000000;
	sram_mem[121762] = 16'b0000000000000000;
	sram_mem[121763] = 16'b0000000000000000;
	sram_mem[121764] = 16'b0000000000000000;
	sram_mem[121765] = 16'b0000000000000000;
	sram_mem[121766] = 16'b0000000000000000;
	sram_mem[121767] = 16'b0000000000000000;
	sram_mem[121768] = 16'b0000000000000000;
	sram_mem[121769] = 16'b0000000000000000;
	sram_mem[121770] = 16'b0000000000000000;
	sram_mem[121771] = 16'b0000000000000000;
	sram_mem[121772] = 16'b0000000000000000;
	sram_mem[121773] = 16'b0000000000000000;
	sram_mem[121774] = 16'b0000000000000000;
	sram_mem[121775] = 16'b0000000000000000;
	sram_mem[121776] = 16'b0000000000000000;
	sram_mem[121777] = 16'b0000000000000000;
	sram_mem[121778] = 16'b0000000000000000;
	sram_mem[121779] = 16'b0000000000000000;
	sram_mem[121780] = 16'b0000000000000000;
	sram_mem[121781] = 16'b0000000000000000;
	sram_mem[121782] = 16'b0000000000000000;
	sram_mem[121783] = 16'b0000000000000000;
	sram_mem[121784] = 16'b0000000000000000;
	sram_mem[121785] = 16'b0000000000000000;
	sram_mem[121786] = 16'b0000000000000000;
	sram_mem[121787] = 16'b0000000000000000;
	sram_mem[121788] = 16'b0000000000000000;
	sram_mem[121789] = 16'b0000000000000000;
	sram_mem[121790] = 16'b0000000000000000;
	sram_mem[121791] = 16'b0000000000000000;
	sram_mem[121792] = 16'b0000000000000000;
	sram_mem[121793] = 16'b0000000000000000;
	sram_mem[121794] = 16'b0000000000000000;
	sram_mem[121795] = 16'b0000000000000000;
	sram_mem[121796] = 16'b0000000000000000;
	sram_mem[121797] = 16'b0000000000000000;
	sram_mem[121798] = 16'b0000000000000000;
	sram_mem[121799] = 16'b0000000000000000;
	sram_mem[121800] = 16'b0000000000000000;
	sram_mem[121801] = 16'b0000000000000000;
	sram_mem[121802] = 16'b0000000000000000;
	sram_mem[121803] = 16'b0000000000000000;
	sram_mem[121804] = 16'b0000000000000000;
	sram_mem[121805] = 16'b0000000000000000;
	sram_mem[121806] = 16'b0000000000000000;
	sram_mem[121807] = 16'b0000000000000000;
	sram_mem[121808] = 16'b0000000000000000;
	sram_mem[121809] = 16'b0000000000000000;
	sram_mem[121810] = 16'b0000000000000000;
	sram_mem[121811] = 16'b0000000000000000;
	sram_mem[121812] = 16'b0000000000000000;
	sram_mem[121813] = 16'b0000000000000000;
	sram_mem[121814] = 16'b0000000000000000;
	sram_mem[121815] = 16'b0000000000000000;
	sram_mem[121816] = 16'b0000000000000000;
	sram_mem[121817] = 16'b0000000000000000;
	sram_mem[121818] = 16'b0000000000000000;
	sram_mem[121819] = 16'b0000000000000000;
	sram_mem[121820] = 16'b0000000000000000;
	sram_mem[121821] = 16'b0000000000000000;
	sram_mem[121822] = 16'b0000000000000000;
	sram_mem[121823] = 16'b0000000000000000;
	sram_mem[121824] = 16'b0000000000000000;
	sram_mem[121825] = 16'b0000000000000000;
	sram_mem[121826] = 16'b0000000000000000;
	sram_mem[121827] = 16'b0000000000000000;
	sram_mem[121828] = 16'b0000000000000000;
	sram_mem[121829] = 16'b0000000000000000;
	sram_mem[121830] = 16'b0000000000000000;
	sram_mem[121831] = 16'b0000000000000000;
	sram_mem[121832] = 16'b0000000000000000;
	sram_mem[121833] = 16'b0000000000000000;
	sram_mem[121834] = 16'b0000000000000000;
	sram_mem[121835] = 16'b0000000000000000;
	sram_mem[121836] = 16'b0000000000000000;
	sram_mem[121837] = 16'b0000000000000000;
	sram_mem[121838] = 16'b0000000000000000;
	sram_mem[121839] = 16'b0000000000000000;
	sram_mem[121840] = 16'b0000000000000000;
	sram_mem[121841] = 16'b0000000000000000;
	sram_mem[121842] = 16'b0000000000000000;
	sram_mem[121843] = 16'b0000000000000000;
	sram_mem[121844] = 16'b0000000000000000;
	sram_mem[121845] = 16'b0000000000000000;
	sram_mem[121846] = 16'b0000000000000000;
	sram_mem[121847] = 16'b0000000000000000;
	sram_mem[121848] = 16'b0000000000000000;
	sram_mem[121849] = 16'b0000000000000000;
	sram_mem[121850] = 16'b0000000000000000;
	sram_mem[121851] = 16'b0000000000000000;
	sram_mem[121852] = 16'b0000000000000000;
	sram_mem[121853] = 16'b0000000000000000;
	sram_mem[121854] = 16'b0000000000000000;
	sram_mem[121855] = 16'b0000000000000000;
	sram_mem[121856] = 16'b0000000000000000;
	sram_mem[121857] = 16'b0000000000000000;
	sram_mem[121858] = 16'b0000000000000000;
	sram_mem[121859] = 16'b0000000000000000;
	sram_mem[121860] = 16'b0000000000000000;
	sram_mem[121861] = 16'b0000000000000000;
	sram_mem[121862] = 16'b0000000000000000;
	sram_mem[121863] = 16'b0000000000000000;
	sram_mem[121864] = 16'b0000000000000000;
	sram_mem[121865] = 16'b0000000000000000;
	sram_mem[121866] = 16'b0000000000000000;
	sram_mem[121867] = 16'b0000000000000000;
	sram_mem[121868] = 16'b0000000000000000;
	sram_mem[121869] = 16'b0000000000000000;
	sram_mem[121870] = 16'b0000000000000000;
	sram_mem[121871] = 16'b0000000000000000;
	sram_mem[121872] = 16'b0000000000000000;
	sram_mem[121873] = 16'b0000000000000000;
	sram_mem[121874] = 16'b0000000000000000;
	sram_mem[121875] = 16'b0000000000000000;
	sram_mem[121876] = 16'b0000000000000000;
	sram_mem[121877] = 16'b0000000000000000;
	sram_mem[121878] = 16'b0000000000000000;
	sram_mem[121879] = 16'b0000000000000000;
	sram_mem[121880] = 16'b0000000000000000;
	sram_mem[121881] = 16'b0000000000000000;
	sram_mem[121882] = 16'b0000000000000000;
	sram_mem[121883] = 16'b0000000000000000;
	sram_mem[121884] = 16'b0000000000000000;
	sram_mem[121885] = 16'b0000000000000000;
	sram_mem[121886] = 16'b0000000000000000;
	sram_mem[121887] = 16'b0000000000000000;
	sram_mem[121888] = 16'b0000000000000000;
	sram_mem[121889] = 16'b0000000000000000;
	sram_mem[121890] = 16'b0000000000000000;
	sram_mem[121891] = 16'b0000000000000000;
	sram_mem[121892] = 16'b0000000000000000;
	sram_mem[121893] = 16'b0000000000000000;
	sram_mem[121894] = 16'b0000000000000000;
	sram_mem[121895] = 16'b0000000000000000;
	sram_mem[121896] = 16'b0000000000000000;
	sram_mem[121897] = 16'b0000000000000000;
	sram_mem[121898] = 16'b0000000000000000;
	sram_mem[121899] = 16'b0000000000000000;
	sram_mem[121900] = 16'b0000000000000000;
	sram_mem[121901] = 16'b0000000000000000;
	sram_mem[121902] = 16'b0000000000000000;
	sram_mem[121903] = 16'b0000000000000000;
	sram_mem[121904] = 16'b0000000000000000;
	sram_mem[121905] = 16'b0000000000000000;
	sram_mem[121906] = 16'b0000000000000000;
	sram_mem[121907] = 16'b0000000000000000;
	sram_mem[121908] = 16'b0000000000000000;
	sram_mem[121909] = 16'b0000000000000000;
	sram_mem[121910] = 16'b0000000000000000;
	sram_mem[121911] = 16'b0000000000000000;
	sram_mem[121912] = 16'b0000000000000000;
	sram_mem[121913] = 16'b0000000000000000;
	sram_mem[121914] = 16'b0000000000000000;
	sram_mem[121915] = 16'b0000000000000000;
	sram_mem[121916] = 16'b0000000000000000;
	sram_mem[121917] = 16'b0000000000000000;
	sram_mem[121918] = 16'b0000000000000000;
	sram_mem[121919] = 16'b0000000000000000;
	sram_mem[121920] = 16'b0000000000000000;
	sram_mem[121921] = 16'b0000000000000000;
	sram_mem[121922] = 16'b0000000000000000;
	sram_mem[121923] = 16'b0000000000000000;
	sram_mem[121924] = 16'b0000000000000000;
	sram_mem[121925] = 16'b0000000000000000;
	sram_mem[121926] = 16'b0000000000000000;
	sram_mem[121927] = 16'b0000000000000000;
	sram_mem[121928] = 16'b0000000000000000;
	sram_mem[121929] = 16'b0000000000000000;
	sram_mem[121930] = 16'b0000000000000000;
	sram_mem[121931] = 16'b0000000000000000;
	sram_mem[121932] = 16'b0000000000000000;
	sram_mem[121933] = 16'b0000000000000000;
	sram_mem[121934] = 16'b0000000000000000;
	sram_mem[121935] = 16'b0000000000000000;
	sram_mem[121936] = 16'b0000000000000000;
	sram_mem[121937] = 16'b0000000000000000;
	sram_mem[121938] = 16'b0000000000000000;
	sram_mem[121939] = 16'b0000000000000000;
	sram_mem[121940] = 16'b0000000000000000;
	sram_mem[121941] = 16'b0000000000000000;
	sram_mem[121942] = 16'b0000000000000000;
	sram_mem[121943] = 16'b0000000000000000;
	sram_mem[121944] = 16'b0000000000000000;
	sram_mem[121945] = 16'b0000000000000000;
	sram_mem[121946] = 16'b0000000000000000;
	sram_mem[121947] = 16'b0000000000000000;
	sram_mem[121948] = 16'b0000000000000000;
	sram_mem[121949] = 16'b0000000000000000;
	sram_mem[121950] = 16'b0000000000000000;
	sram_mem[121951] = 16'b0000000000000000;
	sram_mem[121952] = 16'b0000000000000000;
	sram_mem[121953] = 16'b0000000000000000;
	sram_mem[121954] = 16'b0000000000000000;
	sram_mem[121955] = 16'b0000000000000000;
	sram_mem[121956] = 16'b0000000000000000;
	sram_mem[121957] = 16'b0000000000000000;
	sram_mem[121958] = 16'b0000000000000000;
	sram_mem[121959] = 16'b0000000000000000;
	sram_mem[121960] = 16'b0000000000000000;
	sram_mem[121961] = 16'b0000000000000000;
	sram_mem[121962] = 16'b0000000000000000;
	sram_mem[121963] = 16'b0000000000000000;
	sram_mem[121964] = 16'b0000000000000000;
	sram_mem[121965] = 16'b0000000000000000;
	sram_mem[121966] = 16'b0000000000000000;
	sram_mem[121967] = 16'b0000000000000000;
	sram_mem[121968] = 16'b0000000000000000;
	sram_mem[121969] = 16'b0000000000000000;
	sram_mem[121970] = 16'b0000000000000000;
	sram_mem[121971] = 16'b0000000000000000;
	sram_mem[121972] = 16'b0000000000000000;
	sram_mem[121973] = 16'b0000000000000000;
	sram_mem[121974] = 16'b0000000000000000;
	sram_mem[121975] = 16'b0000000000000000;
	sram_mem[121976] = 16'b0000000000000000;
	sram_mem[121977] = 16'b0000000000000000;
	sram_mem[121978] = 16'b0000000000000000;
	sram_mem[121979] = 16'b0000000000000000;
	sram_mem[121980] = 16'b0000000000000000;
	sram_mem[121981] = 16'b0000000000000000;
	sram_mem[121982] = 16'b0000000000000000;
	sram_mem[121983] = 16'b0000000000000000;
	sram_mem[121984] = 16'b0000000000000000;
	sram_mem[121985] = 16'b0000000000000000;
	sram_mem[121986] = 16'b0000000000000000;
	sram_mem[121987] = 16'b0000000000000000;
	sram_mem[121988] = 16'b0000000000000000;
	sram_mem[121989] = 16'b0000000000000000;
	sram_mem[121990] = 16'b0000000000000000;
	sram_mem[121991] = 16'b0000000000000000;
	sram_mem[121992] = 16'b0000000000000000;
	sram_mem[121993] = 16'b0000000000000000;
	sram_mem[121994] = 16'b0000000000000000;
	sram_mem[121995] = 16'b0000000000000000;
	sram_mem[121996] = 16'b0000000000000000;
	sram_mem[121997] = 16'b0000000000000000;
	sram_mem[121998] = 16'b0000000000000000;
	sram_mem[121999] = 16'b0000000000000000;
	sram_mem[122000] = 16'b0000000000000000;
	sram_mem[122001] = 16'b0000000000000000;
	sram_mem[122002] = 16'b0000000000000000;
	sram_mem[122003] = 16'b0000000000000000;
	sram_mem[122004] = 16'b0000000000000000;
	sram_mem[122005] = 16'b0000000000000000;
	sram_mem[122006] = 16'b0000000000000000;
	sram_mem[122007] = 16'b0000000000000000;
	sram_mem[122008] = 16'b0000000000000000;
	sram_mem[122009] = 16'b0000000000000000;
	sram_mem[122010] = 16'b0000000000000000;
	sram_mem[122011] = 16'b0000000000000000;
	sram_mem[122012] = 16'b0000000000000000;
	sram_mem[122013] = 16'b0000000000000000;
	sram_mem[122014] = 16'b0000000000000000;
	sram_mem[122015] = 16'b0000000000000000;
	sram_mem[122016] = 16'b0000000000000000;
	sram_mem[122017] = 16'b0000000000000000;
	sram_mem[122018] = 16'b0000000000000000;
	sram_mem[122019] = 16'b0000000000000000;
	sram_mem[122020] = 16'b0000000000000000;
	sram_mem[122021] = 16'b0000000000000000;
	sram_mem[122022] = 16'b0000000000000000;
	sram_mem[122023] = 16'b0000000000000000;
	sram_mem[122024] = 16'b0000000000000000;
	sram_mem[122025] = 16'b0000000000000000;
	sram_mem[122026] = 16'b0000000000000000;
	sram_mem[122027] = 16'b0000000000000000;
	sram_mem[122028] = 16'b0000000000000000;
	sram_mem[122029] = 16'b0000000000000000;
	sram_mem[122030] = 16'b0000000000000000;
	sram_mem[122031] = 16'b0000000000000000;
	sram_mem[122032] = 16'b0000000000000000;
	sram_mem[122033] = 16'b0000000000000000;
	sram_mem[122034] = 16'b0000000000000000;
	sram_mem[122035] = 16'b0000000000000000;
	sram_mem[122036] = 16'b0000000000000000;
	sram_mem[122037] = 16'b0000000000000000;
	sram_mem[122038] = 16'b0000000000000000;
	sram_mem[122039] = 16'b0000000000000000;
	sram_mem[122040] = 16'b0000000000000000;
	sram_mem[122041] = 16'b0000000000000000;
	sram_mem[122042] = 16'b0000000000000000;
	sram_mem[122043] = 16'b0000000000000000;
	sram_mem[122044] = 16'b0000000000000000;
	sram_mem[122045] = 16'b0000000000000000;
	sram_mem[122046] = 16'b0000000000000000;
	sram_mem[122047] = 16'b0000000000000000;
	sram_mem[122048] = 16'b0000000000000000;
	sram_mem[122049] = 16'b0000000000000000;
	sram_mem[122050] = 16'b0000000000000000;
	sram_mem[122051] = 16'b0000000000000000;
	sram_mem[122052] = 16'b0000000000000000;
	sram_mem[122053] = 16'b0000000000000000;
	sram_mem[122054] = 16'b0000000000000000;
	sram_mem[122055] = 16'b0000000000000000;
	sram_mem[122056] = 16'b0000000000000000;
	sram_mem[122057] = 16'b0000000000000000;
	sram_mem[122058] = 16'b0000000000000000;
	sram_mem[122059] = 16'b0000000000000000;
	sram_mem[122060] = 16'b0000000000000000;
	sram_mem[122061] = 16'b0000000000000000;
	sram_mem[122062] = 16'b0000000000000000;
	sram_mem[122063] = 16'b0000000000000000;
	sram_mem[122064] = 16'b0000000000000000;
	sram_mem[122065] = 16'b0000000000000000;
	sram_mem[122066] = 16'b0000000000000000;
	sram_mem[122067] = 16'b0000000000000000;
	sram_mem[122068] = 16'b0000000000000000;
	sram_mem[122069] = 16'b0000000000000000;
	sram_mem[122070] = 16'b0000000000000000;
	sram_mem[122071] = 16'b0000000000000000;
	sram_mem[122072] = 16'b0000000000000000;
	sram_mem[122073] = 16'b0000000000000000;
	sram_mem[122074] = 16'b0000000000000000;
	sram_mem[122075] = 16'b0000000000000000;
	sram_mem[122076] = 16'b0000000000000000;
	sram_mem[122077] = 16'b0000000000000000;
	sram_mem[122078] = 16'b0000000000000000;
	sram_mem[122079] = 16'b0000000000000000;
	sram_mem[122080] = 16'b0000000000000000;
	sram_mem[122081] = 16'b0000000000000000;
	sram_mem[122082] = 16'b0000000000000000;
	sram_mem[122083] = 16'b0000000000000000;
	sram_mem[122084] = 16'b0000000000000000;
	sram_mem[122085] = 16'b0000000000000000;
	sram_mem[122086] = 16'b0000000000000000;
	sram_mem[122087] = 16'b0000000000000000;
	sram_mem[122088] = 16'b0000000000000000;
	sram_mem[122089] = 16'b0000000000000000;
	sram_mem[122090] = 16'b0000000000000000;
	sram_mem[122091] = 16'b0000000000000000;
	sram_mem[122092] = 16'b0000000000000000;
	sram_mem[122093] = 16'b0000000000000000;
	sram_mem[122094] = 16'b0000000000000000;
	sram_mem[122095] = 16'b0000000000000000;
	sram_mem[122096] = 16'b0000000000000000;
	sram_mem[122097] = 16'b0000000000000000;
	sram_mem[122098] = 16'b0000000000000000;
	sram_mem[122099] = 16'b0000000000000000;
	sram_mem[122100] = 16'b0000000000000000;
	sram_mem[122101] = 16'b0000000000000000;
	sram_mem[122102] = 16'b0000000000000000;
	sram_mem[122103] = 16'b0000000000000000;
	sram_mem[122104] = 16'b0000000000000000;
	sram_mem[122105] = 16'b0000000000000000;
	sram_mem[122106] = 16'b0000000000000000;
	sram_mem[122107] = 16'b0000000000000000;
	sram_mem[122108] = 16'b0000000000000000;
	sram_mem[122109] = 16'b0000000000000000;
	sram_mem[122110] = 16'b0000000000000000;
	sram_mem[122111] = 16'b0000000000000000;
	sram_mem[122112] = 16'b0000000000000000;
	sram_mem[122113] = 16'b0000000000000000;
	sram_mem[122114] = 16'b0000000000000000;
	sram_mem[122115] = 16'b0000000000000000;
	sram_mem[122116] = 16'b0000000000000000;
	sram_mem[122117] = 16'b0000000000000000;
	sram_mem[122118] = 16'b0000000000000000;
	sram_mem[122119] = 16'b0000000000000000;
	sram_mem[122120] = 16'b0000000000000000;
	sram_mem[122121] = 16'b0000000000000000;
	sram_mem[122122] = 16'b0000000000000000;
	sram_mem[122123] = 16'b0000000000000000;
	sram_mem[122124] = 16'b0000000000000000;
	sram_mem[122125] = 16'b0000000000000000;
	sram_mem[122126] = 16'b0000000000000000;
	sram_mem[122127] = 16'b0000000000000000;
	sram_mem[122128] = 16'b0000000000000000;
	sram_mem[122129] = 16'b0000000000000000;
	sram_mem[122130] = 16'b0000000000000000;
	sram_mem[122131] = 16'b0000000000000000;
	sram_mem[122132] = 16'b0000000000000000;
	sram_mem[122133] = 16'b0000000000000000;
	sram_mem[122134] = 16'b0000000000000000;
	sram_mem[122135] = 16'b0000000000000000;
	sram_mem[122136] = 16'b0000000000000000;
	sram_mem[122137] = 16'b0000000000000000;
	sram_mem[122138] = 16'b0000000000000000;
	sram_mem[122139] = 16'b0000000000000000;
	sram_mem[122140] = 16'b0000000000000000;
	sram_mem[122141] = 16'b0000000000000000;
	sram_mem[122142] = 16'b0000000000000000;
	sram_mem[122143] = 16'b0000000000000000;
	sram_mem[122144] = 16'b0000000000000000;
	sram_mem[122145] = 16'b0000000000000000;
	sram_mem[122146] = 16'b0000000000000000;
	sram_mem[122147] = 16'b0000000000000000;
	sram_mem[122148] = 16'b0000000000000000;
	sram_mem[122149] = 16'b0000000000000000;
	sram_mem[122150] = 16'b0000000000000000;
	sram_mem[122151] = 16'b0000000000000000;
	sram_mem[122152] = 16'b0000000000000000;
	sram_mem[122153] = 16'b0000000000000000;
	sram_mem[122154] = 16'b0000000000000000;
	sram_mem[122155] = 16'b0000000000000000;
	sram_mem[122156] = 16'b0000000000000000;
	sram_mem[122157] = 16'b0000000000000000;
	sram_mem[122158] = 16'b0000000000000000;
	sram_mem[122159] = 16'b0000000000000000;
	sram_mem[122160] = 16'b0000000000000000;
	sram_mem[122161] = 16'b0000000000000000;
	sram_mem[122162] = 16'b0000000000000000;
	sram_mem[122163] = 16'b0000000000000000;
	sram_mem[122164] = 16'b0000000000000000;
	sram_mem[122165] = 16'b0000000000000000;
	sram_mem[122166] = 16'b0000000000000000;
	sram_mem[122167] = 16'b0000000000000000;
	sram_mem[122168] = 16'b0000000000000000;
	sram_mem[122169] = 16'b0000000000000000;
	sram_mem[122170] = 16'b0000000000000000;
	sram_mem[122171] = 16'b0000000000000000;
	sram_mem[122172] = 16'b0000000000000000;
	sram_mem[122173] = 16'b0000000000000000;
	sram_mem[122174] = 16'b0000000000000000;
	sram_mem[122175] = 16'b0000000000000000;
	sram_mem[122176] = 16'b0000000000000000;
	sram_mem[122177] = 16'b0000000000000000;
	sram_mem[122178] = 16'b0000000000000000;
	sram_mem[122179] = 16'b0000000000000000;
	sram_mem[122180] = 16'b0000000000000000;
	sram_mem[122181] = 16'b0000000000000000;
	sram_mem[122182] = 16'b0000000000000000;
	sram_mem[122183] = 16'b0000000000000000;
	sram_mem[122184] = 16'b0000000000000000;
	sram_mem[122185] = 16'b0000000000000000;
	sram_mem[122186] = 16'b0000000000000000;
	sram_mem[122187] = 16'b0000000000000000;
	sram_mem[122188] = 16'b0000000000000000;
	sram_mem[122189] = 16'b0000000000000000;
	sram_mem[122190] = 16'b0000000000000000;
	sram_mem[122191] = 16'b0000000000000000;
	sram_mem[122192] = 16'b0000000000000000;
	sram_mem[122193] = 16'b0000000000000000;
	sram_mem[122194] = 16'b0000000000000000;
	sram_mem[122195] = 16'b0000000000000000;
	sram_mem[122196] = 16'b0000000000000000;
	sram_mem[122197] = 16'b0000000000000000;
	sram_mem[122198] = 16'b0000000000000000;
	sram_mem[122199] = 16'b0000000000000000;
	sram_mem[122200] = 16'b0000000000000000;
	sram_mem[122201] = 16'b0000000000000000;
	sram_mem[122202] = 16'b0000000000000000;
	sram_mem[122203] = 16'b0000000000000000;
	sram_mem[122204] = 16'b0000000000000000;
	sram_mem[122205] = 16'b0000000000000000;
	sram_mem[122206] = 16'b0000000000000000;
	sram_mem[122207] = 16'b0000000000000000;
	sram_mem[122208] = 16'b0000000000000000;
	sram_mem[122209] = 16'b0000000000000000;
	sram_mem[122210] = 16'b0000000000000000;
	sram_mem[122211] = 16'b0000000000000000;
	sram_mem[122212] = 16'b0000000000000000;
	sram_mem[122213] = 16'b0000000000000000;
	sram_mem[122214] = 16'b0000000000000000;
	sram_mem[122215] = 16'b0000000000000000;
	sram_mem[122216] = 16'b0000000000000000;
	sram_mem[122217] = 16'b0000000000000000;
	sram_mem[122218] = 16'b0000000000000000;
	sram_mem[122219] = 16'b0000000000000000;
	sram_mem[122220] = 16'b0000000000000000;
	sram_mem[122221] = 16'b0000000000000000;
	sram_mem[122222] = 16'b0000000000000000;
	sram_mem[122223] = 16'b0000000000000000;
	sram_mem[122224] = 16'b0000000000000000;
	sram_mem[122225] = 16'b0000000000000000;
	sram_mem[122226] = 16'b0000000000000000;
	sram_mem[122227] = 16'b0000000000000000;
	sram_mem[122228] = 16'b0000000000000000;
	sram_mem[122229] = 16'b0000000000000000;
	sram_mem[122230] = 16'b0000000000000000;
	sram_mem[122231] = 16'b0000000000000000;
	sram_mem[122232] = 16'b0000000000000000;
	sram_mem[122233] = 16'b0000000000000000;
	sram_mem[122234] = 16'b0000000000000000;
	sram_mem[122235] = 16'b0000000000000000;
	sram_mem[122236] = 16'b0000000000000000;
	sram_mem[122237] = 16'b0000000000000000;
	sram_mem[122238] = 16'b0000000000000000;
	sram_mem[122239] = 16'b0000000000000000;
	sram_mem[122240] = 16'b0000000000000000;
	sram_mem[122241] = 16'b0000000000000000;
	sram_mem[122242] = 16'b0000000000000000;
	sram_mem[122243] = 16'b0000000000000000;
	sram_mem[122244] = 16'b0000000000000000;
	sram_mem[122245] = 16'b0000000000000000;
	sram_mem[122246] = 16'b0000000000000000;
	sram_mem[122247] = 16'b0000000000000000;
	sram_mem[122248] = 16'b0000000000000000;
	sram_mem[122249] = 16'b0000000000000000;
	sram_mem[122250] = 16'b0000000000000000;
	sram_mem[122251] = 16'b0000000000000000;
	sram_mem[122252] = 16'b0000000000000000;
	sram_mem[122253] = 16'b0000000000000000;
	sram_mem[122254] = 16'b0000000000000000;
	sram_mem[122255] = 16'b0000000000000000;
	sram_mem[122256] = 16'b0000000000000000;
	sram_mem[122257] = 16'b0000000000000000;
	sram_mem[122258] = 16'b0000000000000000;
	sram_mem[122259] = 16'b0000000000000000;
	sram_mem[122260] = 16'b0000000000000000;
	sram_mem[122261] = 16'b0000000000000000;
	sram_mem[122262] = 16'b0000000000000000;
	sram_mem[122263] = 16'b0000000000000000;
	sram_mem[122264] = 16'b0000000000000000;
	sram_mem[122265] = 16'b0000000000000000;
	sram_mem[122266] = 16'b0000000000000000;
	sram_mem[122267] = 16'b0000000000000000;
	sram_mem[122268] = 16'b0000000000000000;
	sram_mem[122269] = 16'b0000000000000000;
	sram_mem[122270] = 16'b0000000000000000;
	sram_mem[122271] = 16'b0000000000000000;
	sram_mem[122272] = 16'b0000000000000000;
	sram_mem[122273] = 16'b0000000000000000;
	sram_mem[122274] = 16'b0000000000000000;
	sram_mem[122275] = 16'b0000000000000000;
	sram_mem[122276] = 16'b0000000000000000;
	sram_mem[122277] = 16'b0000000000000000;
	sram_mem[122278] = 16'b0000000000000000;
	sram_mem[122279] = 16'b0000000000000000;
	sram_mem[122280] = 16'b0000000000000000;
	sram_mem[122281] = 16'b0000000000000000;
	sram_mem[122282] = 16'b0000000000000000;
	sram_mem[122283] = 16'b0000000000000000;
	sram_mem[122284] = 16'b0000000000000000;
	sram_mem[122285] = 16'b0000000000000000;
	sram_mem[122286] = 16'b0000000000000000;
	sram_mem[122287] = 16'b0000000000000000;
	sram_mem[122288] = 16'b0000000000000000;
	sram_mem[122289] = 16'b0000000000000000;
	sram_mem[122290] = 16'b0000000000000000;
	sram_mem[122291] = 16'b0000000000000000;
	sram_mem[122292] = 16'b0000000000000000;
	sram_mem[122293] = 16'b0000000000000000;
	sram_mem[122294] = 16'b0000000000000000;
	sram_mem[122295] = 16'b0000000000000000;
	sram_mem[122296] = 16'b0000000000000000;
	sram_mem[122297] = 16'b0000000000000000;
	sram_mem[122298] = 16'b0000000000000000;
	sram_mem[122299] = 16'b0000000000000000;
	sram_mem[122300] = 16'b0000000000000000;
	sram_mem[122301] = 16'b0000000000000000;
	sram_mem[122302] = 16'b0000000000000000;
	sram_mem[122303] = 16'b0000000000000000;
	sram_mem[122304] = 16'b0000000000000000;
	sram_mem[122305] = 16'b0000000000000000;
	sram_mem[122306] = 16'b0000000000000000;
	sram_mem[122307] = 16'b0000000000000000;
	sram_mem[122308] = 16'b0000000000000000;
	sram_mem[122309] = 16'b0000000000000000;
	sram_mem[122310] = 16'b0000000000000000;
	sram_mem[122311] = 16'b0000000000000000;
	sram_mem[122312] = 16'b0000000000000000;
	sram_mem[122313] = 16'b0000000000000000;
	sram_mem[122314] = 16'b0000000000000000;
	sram_mem[122315] = 16'b0000000000000000;
	sram_mem[122316] = 16'b0000000000000000;
	sram_mem[122317] = 16'b0000000000000000;
	sram_mem[122318] = 16'b0000000000000000;
	sram_mem[122319] = 16'b0000000000000000;
	sram_mem[122320] = 16'b0000000000000000;
	sram_mem[122321] = 16'b0000000000000000;
	sram_mem[122322] = 16'b0000000000000000;
	sram_mem[122323] = 16'b0000000000000000;
	sram_mem[122324] = 16'b0000000000000000;
	sram_mem[122325] = 16'b0000000000000000;
	sram_mem[122326] = 16'b0000000000000000;
	sram_mem[122327] = 16'b0000000000000000;
	sram_mem[122328] = 16'b0000000000000000;
	sram_mem[122329] = 16'b0000000000000000;
	sram_mem[122330] = 16'b0000000000000000;
	sram_mem[122331] = 16'b0000000000000000;
	sram_mem[122332] = 16'b0000000000000000;
	sram_mem[122333] = 16'b0000000000000000;
	sram_mem[122334] = 16'b0000000000000000;
	sram_mem[122335] = 16'b0000000000000000;
	sram_mem[122336] = 16'b0000000000000000;
	sram_mem[122337] = 16'b0000000000000000;
	sram_mem[122338] = 16'b0000000000000000;
	sram_mem[122339] = 16'b0000000000000000;
	sram_mem[122340] = 16'b0000000000000000;
	sram_mem[122341] = 16'b0000000000000000;
	sram_mem[122342] = 16'b0000000000000000;
	sram_mem[122343] = 16'b0000000000000000;
	sram_mem[122344] = 16'b0000000000000000;
	sram_mem[122345] = 16'b0000000000000000;
	sram_mem[122346] = 16'b0000000000000000;
	sram_mem[122347] = 16'b0000000000000000;
	sram_mem[122348] = 16'b0000000000000000;
	sram_mem[122349] = 16'b0000000000000000;
	sram_mem[122350] = 16'b0000000000000000;
	sram_mem[122351] = 16'b0000000000000000;
	sram_mem[122352] = 16'b0000000000000000;
	sram_mem[122353] = 16'b0000000000000000;
	sram_mem[122354] = 16'b0000000000000000;
	sram_mem[122355] = 16'b0000000000000000;
	sram_mem[122356] = 16'b0000000000000000;
	sram_mem[122357] = 16'b0000000000000000;
	sram_mem[122358] = 16'b0000000000000000;
	sram_mem[122359] = 16'b0000000000000000;
	sram_mem[122360] = 16'b0000000000000000;
	sram_mem[122361] = 16'b0000000000000000;
	sram_mem[122362] = 16'b0000000000000000;
	sram_mem[122363] = 16'b0000000000000000;
	sram_mem[122364] = 16'b0000000000000000;
	sram_mem[122365] = 16'b0000000000000000;
	sram_mem[122366] = 16'b0000000000000000;
	sram_mem[122367] = 16'b0000000000000000;
	sram_mem[122368] = 16'b0000000000000000;
	sram_mem[122369] = 16'b0000000000000000;
	sram_mem[122370] = 16'b0000000000000000;
	sram_mem[122371] = 16'b0000000000000000;
	sram_mem[122372] = 16'b0000000000000000;
	sram_mem[122373] = 16'b0000000000000000;
	sram_mem[122374] = 16'b0000000000000000;
	sram_mem[122375] = 16'b0000000000000000;
	sram_mem[122376] = 16'b0000000000000000;
	sram_mem[122377] = 16'b0000000000000000;
	sram_mem[122378] = 16'b0000000000000000;
	sram_mem[122379] = 16'b0000000000000000;
	sram_mem[122380] = 16'b0000000000000000;
	sram_mem[122381] = 16'b0000000000000000;
	sram_mem[122382] = 16'b0000000000000000;
	sram_mem[122383] = 16'b0000000000000000;
	sram_mem[122384] = 16'b0000000000000000;
	sram_mem[122385] = 16'b0000000000000000;
	sram_mem[122386] = 16'b0000000000000000;
	sram_mem[122387] = 16'b0000000000000000;
	sram_mem[122388] = 16'b0000000000000000;
	sram_mem[122389] = 16'b0000000000000000;
	sram_mem[122390] = 16'b0000000000000000;
	sram_mem[122391] = 16'b0000000000000000;
	sram_mem[122392] = 16'b0000000000000000;
	sram_mem[122393] = 16'b0000000000000000;
	sram_mem[122394] = 16'b0000000000000000;
	sram_mem[122395] = 16'b0000000000000000;
	sram_mem[122396] = 16'b0000000000000000;
	sram_mem[122397] = 16'b0000000000000000;
	sram_mem[122398] = 16'b0000000000000000;
	sram_mem[122399] = 16'b0000000000000000;
	sram_mem[122400] = 16'b0000000000000000;
	sram_mem[122401] = 16'b0000000000000000;
	sram_mem[122402] = 16'b0000000000000000;
	sram_mem[122403] = 16'b0000000000000000;
	sram_mem[122404] = 16'b0000000000000000;
	sram_mem[122405] = 16'b0000000000000000;
	sram_mem[122406] = 16'b0000000000000000;
	sram_mem[122407] = 16'b0000000000000000;
	sram_mem[122408] = 16'b0000000000000000;
	sram_mem[122409] = 16'b0000000000000000;
	sram_mem[122410] = 16'b0000000000000000;
	sram_mem[122411] = 16'b0000000000000000;
	sram_mem[122412] = 16'b0000000000000000;
	sram_mem[122413] = 16'b0000000000000000;
	sram_mem[122414] = 16'b0000000000000000;
	sram_mem[122415] = 16'b0000000000000000;
	sram_mem[122416] = 16'b0000000000000000;
	sram_mem[122417] = 16'b0000000000000000;
	sram_mem[122418] = 16'b0000000000000000;
	sram_mem[122419] = 16'b0000000000000000;
	sram_mem[122420] = 16'b0000000000000000;
	sram_mem[122421] = 16'b0000000000000000;
	sram_mem[122422] = 16'b0000000000000000;
	sram_mem[122423] = 16'b0000000000000000;
	sram_mem[122424] = 16'b0000000000000000;
	sram_mem[122425] = 16'b0000000000000000;
	sram_mem[122426] = 16'b0000000000000000;
	sram_mem[122427] = 16'b0000000000000000;
	sram_mem[122428] = 16'b0000000000000000;
	sram_mem[122429] = 16'b0000000000000000;
	sram_mem[122430] = 16'b0000000000000000;
	sram_mem[122431] = 16'b0000000000000000;
	sram_mem[122432] = 16'b0000000000000000;
	sram_mem[122433] = 16'b0000000000000000;
	sram_mem[122434] = 16'b0000000000000000;
	sram_mem[122435] = 16'b0000000000000000;
	sram_mem[122436] = 16'b0000000000000000;
	sram_mem[122437] = 16'b0000000000000000;
	sram_mem[122438] = 16'b0000000000000000;
	sram_mem[122439] = 16'b0000000000000000;
	sram_mem[122440] = 16'b0000000000000000;
	sram_mem[122441] = 16'b0000000000000000;
	sram_mem[122442] = 16'b0000000000000000;
	sram_mem[122443] = 16'b0000000000000000;
	sram_mem[122444] = 16'b0000000000000000;
	sram_mem[122445] = 16'b0000000000000000;
	sram_mem[122446] = 16'b0000000000000000;
	sram_mem[122447] = 16'b0000000000000000;
	sram_mem[122448] = 16'b0000000000000000;
	sram_mem[122449] = 16'b0000000000000000;
	sram_mem[122450] = 16'b0000000000000000;
	sram_mem[122451] = 16'b0000000000000000;
	sram_mem[122452] = 16'b0000000000000000;
	sram_mem[122453] = 16'b0000000000000000;
	sram_mem[122454] = 16'b0000000000000000;
	sram_mem[122455] = 16'b0000000000000000;
	sram_mem[122456] = 16'b0000000000000000;
	sram_mem[122457] = 16'b0000000000000000;
	sram_mem[122458] = 16'b0000000000000000;
	sram_mem[122459] = 16'b0000000000000000;
	sram_mem[122460] = 16'b0000000000000000;
	sram_mem[122461] = 16'b0000000000000000;
	sram_mem[122462] = 16'b0000000000000000;
	sram_mem[122463] = 16'b0000000000000000;
	sram_mem[122464] = 16'b0000000000000000;
	sram_mem[122465] = 16'b0000000000000000;
	sram_mem[122466] = 16'b0000000000000000;
	sram_mem[122467] = 16'b0000000000000000;
	sram_mem[122468] = 16'b0000000000000000;
	sram_mem[122469] = 16'b0000000000000000;
	sram_mem[122470] = 16'b0000000000000000;
	sram_mem[122471] = 16'b0000000000000000;
	sram_mem[122472] = 16'b0000000000000000;
	sram_mem[122473] = 16'b0000000000000000;
	sram_mem[122474] = 16'b0000000000000000;
	sram_mem[122475] = 16'b0000000000000000;
	sram_mem[122476] = 16'b0000000000000000;
	sram_mem[122477] = 16'b0000000000000000;
	sram_mem[122478] = 16'b0000000000000000;
	sram_mem[122479] = 16'b0000000000000000;
	sram_mem[122480] = 16'b0000000000000000;
	sram_mem[122481] = 16'b0000000000000000;
	sram_mem[122482] = 16'b0000000000000000;
	sram_mem[122483] = 16'b0000000000000000;
	sram_mem[122484] = 16'b0000000000000000;
	sram_mem[122485] = 16'b0000000000000000;
	sram_mem[122486] = 16'b0000000000000000;
	sram_mem[122487] = 16'b0000000000000000;
	sram_mem[122488] = 16'b0000000000000000;
	sram_mem[122489] = 16'b0000000000000000;
	sram_mem[122490] = 16'b0000000000000000;
	sram_mem[122491] = 16'b0000000000000000;
	sram_mem[122492] = 16'b0000000000000000;
	sram_mem[122493] = 16'b0000000000000000;
	sram_mem[122494] = 16'b0000000000000000;
	sram_mem[122495] = 16'b0000000000000000;
	sram_mem[122496] = 16'b0000000000000000;
	sram_mem[122497] = 16'b0000000000000000;
	sram_mem[122498] = 16'b0000000000000000;
	sram_mem[122499] = 16'b0000000000000000;
	sram_mem[122500] = 16'b0000000000000000;
	sram_mem[122501] = 16'b0000000000000000;
	sram_mem[122502] = 16'b0000000000000000;
	sram_mem[122503] = 16'b0000000000000000;
	sram_mem[122504] = 16'b0000000000000000;
	sram_mem[122505] = 16'b0000000000000000;
	sram_mem[122506] = 16'b0000000000000000;
	sram_mem[122507] = 16'b0000000000000000;
	sram_mem[122508] = 16'b0000000000000000;
	sram_mem[122509] = 16'b0000000000000000;
	sram_mem[122510] = 16'b0000000000000000;
	sram_mem[122511] = 16'b0000000000000000;
	sram_mem[122512] = 16'b0000000000000000;
	sram_mem[122513] = 16'b0000000000000000;
	sram_mem[122514] = 16'b0000000000000000;
	sram_mem[122515] = 16'b0000000000000000;
	sram_mem[122516] = 16'b0000000000000000;
	sram_mem[122517] = 16'b0000000000000000;
	sram_mem[122518] = 16'b0000000000000000;
	sram_mem[122519] = 16'b0000000000000000;
	sram_mem[122520] = 16'b0000000000000000;
	sram_mem[122521] = 16'b0000000000000000;
	sram_mem[122522] = 16'b0000000000000000;
	sram_mem[122523] = 16'b0000000000000000;
	sram_mem[122524] = 16'b0000000000000000;
	sram_mem[122525] = 16'b0000000000000000;
	sram_mem[122526] = 16'b0000000000000000;
	sram_mem[122527] = 16'b0000000000000000;
	sram_mem[122528] = 16'b0000000000000000;
	sram_mem[122529] = 16'b0000000000000000;
	sram_mem[122530] = 16'b0000000000000000;
	sram_mem[122531] = 16'b0000000000000000;
	sram_mem[122532] = 16'b0000000000000000;
	sram_mem[122533] = 16'b0000000000000000;
	sram_mem[122534] = 16'b0000000000000000;
	sram_mem[122535] = 16'b0000000000000000;
	sram_mem[122536] = 16'b0000000000000000;
	sram_mem[122537] = 16'b0000000000000000;
	sram_mem[122538] = 16'b0000000000000000;
	sram_mem[122539] = 16'b0000000000000000;
	sram_mem[122540] = 16'b0000000000000000;
	sram_mem[122541] = 16'b0000000000000000;
	sram_mem[122542] = 16'b0000000000000000;
	sram_mem[122543] = 16'b0000000000000000;
	sram_mem[122544] = 16'b0000000000000000;
	sram_mem[122545] = 16'b0000000000000000;
	sram_mem[122546] = 16'b0000000000000000;
	sram_mem[122547] = 16'b0000000000000000;
	sram_mem[122548] = 16'b0000000000000000;
	sram_mem[122549] = 16'b0000000000000000;
	sram_mem[122550] = 16'b0000000000000000;
	sram_mem[122551] = 16'b0000000000000000;
	sram_mem[122552] = 16'b0000000000000000;
	sram_mem[122553] = 16'b0000000000000000;
	sram_mem[122554] = 16'b0000000000000000;
	sram_mem[122555] = 16'b0000000000000000;
	sram_mem[122556] = 16'b0000000000000000;
	sram_mem[122557] = 16'b0000000000000000;
	sram_mem[122558] = 16'b0000000000000000;
	sram_mem[122559] = 16'b0000000000000000;
	sram_mem[122560] = 16'b0000000000000000;
	sram_mem[122561] = 16'b0000000000000000;
	sram_mem[122562] = 16'b0000000000000000;
	sram_mem[122563] = 16'b0000000000000000;
	sram_mem[122564] = 16'b0000000000000000;
	sram_mem[122565] = 16'b0000000000000000;
	sram_mem[122566] = 16'b0000000000000000;
	sram_mem[122567] = 16'b0000000000000000;
	sram_mem[122568] = 16'b0000000000000000;
	sram_mem[122569] = 16'b0000000000000000;
	sram_mem[122570] = 16'b0000000000000000;
	sram_mem[122571] = 16'b0000000000000000;
	sram_mem[122572] = 16'b0000000000000000;
	sram_mem[122573] = 16'b0000000000000000;
	sram_mem[122574] = 16'b0000000000000000;
	sram_mem[122575] = 16'b0000000000000000;
	sram_mem[122576] = 16'b0000000000000000;
	sram_mem[122577] = 16'b0000000000000000;
	sram_mem[122578] = 16'b0000000000000000;
	sram_mem[122579] = 16'b0000000000000000;
	sram_mem[122580] = 16'b0000000000000000;
	sram_mem[122581] = 16'b0000000000000000;
	sram_mem[122582] = 16'b0000000000000000;
	sram_mem[122583] = 16'b0000000000000000;
	sram_mem[122584] = 16'b0000000000000000;
	sram_mem[122585] = 16'b0000000000000000;
	sram_mem[122586] = 16'b0000000000000000;
	sram_mem[122587] = 16'b0000000000000000;
	sram_mem[122588] = 16'b0000000000000000;
	sram_mem[122589] = 16'b0000000000000000;
	sram_mem[122590] = 16'b0000000000000000;
	sram_mem[122591] = 16'b0000000000000000;
	sram_mem[122592] = 16'b0000000000000000;
	sram_mem[122593] = 16'b0000000000000000;
	sram_mem[122594] = 16'b0000000000000000;
	sram_mem[122595] = 16'b0000000000000000;
	sram_mem[122596] = 16'b0000000000000000;
	sram_mem[122597] = 16'b0000000000000000;
	sram_mem[122598] = 16'b0000000000000000;
	sram_mem[122599] = 16'b0000000000000000;
	sram_mem[122600] = 16'b0000000000000000;
	sram_mem[122601] = 16'b0000000000000000;
	sram_mem[122602] = 16'b0000000000000000;
	sram_mem[122603] = 16'b0000000000000000;
	sram_mem[122604] = 16'b0000000000000000;
	sram_mem[122605] = 16'b0000000000000000;
	sram_mem[122606] = 16'b0000000000000000;
	sram_mem[122607] = 16'b0000000000000000;
	sram_mem[122608] = 16'b0000000000000000;
	sram_mem[122609] = 16'b0000000000000000;
	sram_mem[122610] = 16'b0000000000000000;
	sram_mem[122611] = 16'b0000000000000000;
	sram_mem[122612] = 16'b0000000000000000;
	sram_mem[122613] = 16'b0000000000000000;
	sram_mem[122614] = 16'b0000000000000000;
	sram_mem[122615] = 16'b0000000000000000;
	sram_mem[122616] = 16'b0000000000000000;
	sram_mem[122617] = 16'b0000000000000000;
	sram_mem[122618] = 16'b0000000000000000;
	sram_mem[122619] = 16'b0000000000000000;
	sram_mem[122620] = 16'b0000000000000000;
	sram_mem[122621] = 16'b0000000000000000;
	sram_mem[122622] = 16'b0000000000000000;
	sram_mem[122623] = 16'b0000000000000000;
	sram_mem[122624] = 16'b0000000000000000;
	sram_mem[122625] = 16'b0000000000000000;
	sram_mem[122626] = 16'b0000000000000000;
	sram_mem[122627] = 16'b0000000000000000;
	sram_mem[122628] = 16'b0000000000000000;
	sram_mem[122629] = 16'b0000000000000000;
	sram_mem[122630] = 16'b0000000000000000;
	sram_mem[122631] = 16'b0000000000000000;
	sram_mem[122632] = 16'b0000000000000000;
	sram_mem[122633] = 16'b0000000000000000;
	sram_mem[122634] = 16'b0000000000000000;
	sram_mem[122635] = 16'b0000000000000000;
	sram_mem[122636] = 16'b0000000000000000;
	sram_mem[122637] = 16'b0000000000000000;
	sram_mem[122638] = 16'b0000000000000000;
	sram_mem[122639] = 16'b0000000000000000;
	sram_mem[122640] = 16'b0000000000000000;
	sram_mem[122641] = 16'b0000000000000000;
	sram_mem[122642] = 16'b0000000000000000;
	sram_mem[122643] = 16'b0000000000000000;
	sram_mem[122644] = 16'b0000000000000000;
	sram_mem[122645] = 16'b0000000000000000;
	sram_mem[122646] = 16'b0000000000000000;
	sram_mem[122647] = 16'b0000000000000000;
	sram_mem[122648] = 16'b0000000000000000;
	sram_mem[122649] = 16'b0000000000000000;
	sram_mem[122650] = 16'b0000000000000000;
	sram_mem[122651] = 16'b0000000000000000;
	sram_mem[122652] = 16'b0000000000000000;
	sram_mem[122653] = 16'b0000000000000000;
	sram_mem[122654] = 16'b0000000000000000;
	sram_mem[122655] = 16'b0000000000000000;
	sram_mem[122656] = 16'b0000000000000000;
	sram_mem[122657] = 16'b0000000000000000;
	sram_mem[122658] = 16'b0000000000000000;
	sram_mem[122659] = 16'b0000000000000000;
	sram_mem[122660] = 16'b0000000000000000;
	sram_mem[122661] = 16'b0000000000000000;
	sram_mem[122662] = 16'b0000000000000000;
	sram_mem[122663] = 16'b0000000000000000;
	sram_mem[122664] = 16'b0000000000000000;
	sram_mem[122665] = 16'b0000000000000000;
	sram_mem[122666] = 16'b0000000000000000;
	sram_mem[122667] = 16'b0000000000000000;
	sram_mem[122668] = 16'b0000000000000000;
	sram_mem[122669] = 16'b0000000000000000;
	sram_mem[122670] = 16'b0000000000000000;
	sram_mem[122671] = 16'b0000000000000000;
	sram_mem[122672] = 16'b0000000000000000;
	sram_mem[122673] = 16'b0000000000000000;
	sram_mem[122674] = 16'b0000000000000000;
	sram_mem[122675] = 16'b0000000000000000;
	sram_mem[122676] = 16'b0000000000000000;
	sram_mem[122677] = 16'b0000000000000000;
	sram_mem[122678] = 16'b0000000000000000;
	sram_mem[122679] = 16'b0000000000000000;
	sram_mem[122680] = 16'b0000000000000000;
	sram_mem[122681] = 16'b0000000000000000;
	sram_mem[122682] = 16'b0000000000000000;
	sram_mem[122683] = 16'b0000000000000000;
	sram_mem[122684] = 16'b0000000000000000;
	sram_mem[122685] = 16'b0000000000000000;
	sram_mem[122686] = 16'b0000000000000000;
	sram_mem[122687] = 16'b0000000000000000;
	sram_mem[122688] = 16'b0000000000000000;
	sram_mem[122689] = 16'b0000000000000000;
	sram_mem[122690] = 16'b0000000000000000;
	sram_mem[122691] = 16'b0000000000000000;
	sram_mem[122692] = 16'b0000000000000000;
	sram_mem[122693] = 16'b0000000000000000;
	sram_mem[122694] = 16'b0000000000000000;
	sram_mem[122695] = 16'b0000000000000000;
	sram_mem[122696] = 16'b0000000000000000;
	sram_mem[122697] = 16'b0000000000000000;
	sram_mem[122698] = 16'b0000000000000000;
	sram_mem[122699] = 16'b0000000000000000;
	sram_mem[122700] = 16'b0000000000000000;
	sram_mem[122701] = 16'b0000000000000000;
	sram_mem[122702] = 16'b0000000000000000;
	sram_mem[122703] = 16'b0000000000000000;
	sram_mem[122704] = 16'b0000000000000000;
	sram_mem[122705] = 16'b0000000000000000;
	sram_mem[122706] = 16'b0000000000000000;
	sram_mem[122707] = 16'b0000000000000000;
	sram_mem[122708] = 16'b0000000000000000;
	sram_mem[122709] = 16'b0000000000000000;
	sram_mem[122710] = 16'b0000000000000000;
	sram_mem[122711] = 16'b0000000000000000;
	sram_mem[122712] = 16'b0000000000000000;
	sram_mem[122713] = 16'b0000000000000000;
	sram_mem[122714] = 16'b0000000000000000;
	sram_mem[122715] = 16'b0000000000000000;
	sram_mem[122716] = 16'b0000000000000000;
	sram_mem[122717] = 16'b0000000000000000;
	sram_mem[122718] = 16'b0000000000000000;
	sram_mem[122719] = 16'b0000000000000000;
	sram_mem[122720] = 16'b0000000000000000;
	sram_mem[122721] = 16'b0000000000000000;
	sram_mem[122722] = 16'b0000000000000000;
	sram_mem[122723] = 16'b0000000000000000;
	sram_mem[122724] = 16'b0000000000000000;
	sram_mem[122725] = 16'b0000000000000000;
	sram_mem[122726] = 16'b0000000000000000;
	sram_mem[122727] = 16'b0000000000000000;
	sram_mem[122728] = 16'b0000000000000000;
	sram_mem[122729] = 16'b0000000000000000;
	sram_mem[122730] = 16'b0000000000000000;
	sram_mem[122731] = 16'b0000000000000000;
	sram_mem[122732] = 16'b0000000000000000;
	sram_mem[122733] = 16'b0000000000000000;
	sram_mem[122734] = 16'b0000000000000000;
	sram_mem[122735] = 16'b0000000000000000;
	sram_mem[122736] = 16'b0000000000000000;
	sram_mem[122737] = 16'b0000000000000000;
	sram_mem[122738] = 16'b0000000000000000;
	sram_mem[122739] = 16'b0000000000000000;
	sram_mem[122740] = 16'b0000000000000000;
	sram_mem[122741] = 16'b0000000000000000;
	sram_mem[122742] = 16'b0000000000000000;
	sram_mem[122743] = 16'b0000000000000000;
	sram_mem[122744] = 16'b0000000000000000;
	sram_mem[122745] = 16'b0000000000000000;
	sram_mem[122746] = 16'b0000000000000000;
	sram_mem[122747] = 16'b0000000000000000;
	sram_mem[122748] = 16'b0000000000000000;
	sram_mem[122749] = 16'b0000000000000000;
	sram_mem[122750] = 16'b0000000000000000;
	sram_mem[122751] = 16'b0000000000000000;
	sram_mem[122752] = 16'b0000000000000000;
	sram_mem[122753] = 16'b0000000000000000;
	sram_mem[122754] = 16'b0000000000000000;
	sram_mem[122755] = 16'b0000000000000000;
	sram_mem[122756] = 16'b0000000000000000;
	sram_mem[122757] = 16'b0000000000000000;
	sram_mem[122758] = 16'b0000000000000000;
	sram_mem[122759] = 16'b0000000000000000;
	sram_mem[122760] = 16'b0000000000000000;
	sram_mem[122761] = 16'b0000000000000000;
	sram_mem[122762] = 16'b0000000000000000;
	sram_mem[122763] = 16'b0000000000000000;
	sram_mem[122764] = 16'b0000000000000000;
	sram_mem[122765] = 16'b0000000000000000;
	sram_mem[122766] = 16'b0000000000000000;
	sram_mem[122767] = 16'b0000000000000000;
	sram_mem[122768] = 16'b0000000000000000;
	sram_mem[122769] = 16'b0000000000000000;
	sram_mem[122770] = 16'b0000000000000000;
	sram_mem[122771] = 16'b0000000000000000;
	sram_mem[122772] = 16'b0000000000000000;
	sram_mem[122773] = 16'b0000000000000000;
	sram_mem[122774] = 16'b0000000000000000;
	sram_mem[122775] = 16'b0000000000000000;
	sram_mem[122776] = 16'b0000000000000000;
	sram_mem[122777] = 16'b0000000000000000;
	sram_mem[122778] = 16'b0000000000000000;
	sram_mem[122779] = 16'b0000000000000000;
	sram_mem[122780] = 16'b0000000000000000;
	sram_mem[122781] = 16'b0000000000000000;
	sram_mem[122782] = 16'b0000000000000000;
	sram_mem[122783] = 16'b0000000000000000;
	sram_mem[122784] = 16'b0000000000000000;
	sram_mem[122785] = 16'b0000000000000000;
	sram_mem[122786] = 16'b0000000000000000;
	sram_mem[122787] = 16'b0000000000000000;
	sram_mem[122788] = 16'b0000000000000000;
	sram_mem[122789] = 16'b0000000000000000;
	sram_mem[122790] = 16'b0000000000000000;
	sram_mem[122791] = 16'b0000000000000000;
	sram_mem[122792] = 16'b0000000000000000;
	sram_mem[122793] = 16'b0000000000000000;
	sram_mem[122794] = 16'b0000000000000000;
	sram_mem[122795] = 16'b0000000000000000;
	sram_mem[122796] = 16'b0000000000000000;
	sram_mem[122797] = 16'b0000000000000000;
	sram_mem[122798] = 16'b0000000000000000;
	sram_mem[122799] = 16'b0000000000000000;
	sram_mem[122800] = 16'b0000000000000000;
	sram_mem[122801] = 16'b0000000000000000;
	sram_mem[122802] = 16'b0000000000000000;
	sram_mem[122803] = 16'b0000000000000000;
	sram_mem[122804] = 16'b0000000000000000;
	sram_mem[122805] = 16'b0000000000000000;
	sram_mem[122806] = 16'b0000000000000000;
	sram_mem[122807] = 16'b0000000000000000;
	sram_mem[122808] = 16'b0000000000000000;
	sram_mem[122809] = 16'b0000000000000000;
	sram_mem[122810] = 16'b0000000000000000;
	sram_mem[122811] = 16'b0000000000000000;
	sram_mem[122812] = 16'b0000000000000000;
	sram_mem[122813] = 16'b0000000000000000;
	sram_mem[122814] = 16'b0000000000000000;
	sram_mem[122815] = 16'b0000000000000000;
	sram_mem[122816] = 16'b0000000000000000;
	sram_mem[122817] = 16'b0000000000000000;
	sram_mem[122818] = 16'b0000000000000000;
	sram_mem[122819] = 16'b0000000000000000;
	sram_mem[122820] = 16'b0000000000000000;
	sram_mem[122821] = 16'b0000000000000000;
	sram_mem[122822] = 16'b0000000000000000;
	sram_mem[122823] = 16'b0000000000000000;
	sram_mem[122824] = 16'b0000000000000000;
	sram_mem[122825] = 16'b0000000000000000;
	sram_mem[122826] = 16'b0000000000000000;
	sram_mem[122827] = 16'b0000000000000000;
	sram_mem[122828] = 16'b0000000000000000;
	sram_mem[122829] = 16'b0000000000000000;
	sram_mem[122830] = 16'b0000000000000000;
	sram_mem[122831] = 16'b0000000000000000;
	sram_mem[122832] = 16'b0000000000000000;
	sram_mem[122833] = 16'b0000000000000000;
	sram_mem[122834] = 16'b0000000000000000;
	sram_mem[122835] = 16'b0000000000000000;
	sram_mem[122836] = 16'b0000000000000000;
	sram_mem[122837] = 16'b0000000000000000;
	sram_mem[122838] = 16'b0000000000000000;
	sram_mem[122839] = 16'b0000000000000000;
	sram_mem[122840] = 16'b0000000000000000;
	sram_mem[122841] = 16'b0000000000000000;
	sram_mem[122842] = 16'b0000000000000000;
	sram_mem[122843] = 16'b0000000000000000;
	sram_mem[122844] = 16'b0000000000000000;
	sram_mem[122845] = 16'b0000000000000000;
	sram_mem[122846] = 16'b0000000000000000;
	sram_mem[122847] = 16'b0000000000000000;
	sram_mem[122848] = 16'b0000000000000000;
	sram_mem[122849] = 16'b0000000000000000;
	sram_mem[122850] = 16'b0000000000000000;
	sram_mem[122851] = 16'b0000000000000000;
	sram_mem[122852] = 16'b0000000000000000;
	sram_mem[122853] = 16'b0000000000000000;
	sram_mem[122854] = 16'b0000000000000000;
	sram_mem[122855] = 16'b0000000000000000;
	sram_mem[122856] = 16'b0000000000000000;
	sram_mem[122857] = 16'b0000000000000000;
	sram_mem[122858] = 16'b0000000000000000;
	sram_mem[122859] = 16'b0000000000000000;
	sram_mem[122860] = 16'b0000000000000000;
	sram_mem[122861] = 16'b0000000000000000;
	sram_mem[122862] = 16'b0000000000000000;
	sram_mem[122863] = 16'b0000000000000000;
	sram_mem[122864] = 16'b0000000000000000;
	sram_mem[122865] = 16'b0000000000000000;
	sram_mem[122866] = 16'b0000000000000000;
	sram_mem[122867] = 16'b0000000000000000;
	sram_mem[122868] = 16'b0000000000000000;
	sram_mem[122869] = 16'b0000000000000000;
	sram_mem[122870] = 16'b0000000000000000;
	sram_mem[122871] = 16'b0000000000000000;
	sram_mem[122872] = 16'b0000000000000000;
	sram_mem[122873] = 16'b0000000000000000;
	sram_mem[122874] = 16'b0000000000000000;
	sram_mem[122875] = 16'b0000000000000000;
	sram_mem[122876] = 16'b0000000000000000;
	sram_mem[122877] = 16'b0000000000000000;
	sram_mem[122878] = 16'b0000000000000000;
	sram_mem[122879] = 16'b0000000000000000;
	sram_mem[122880] = 16'b0000000000000000;
	sram_mem[122881] = 16'b0000000000000000;
	sram_mem[122882] = 16'b0000000000000000;
	sram_mem[122883] = 16'b0000000000000000;
	sram_mem[122884] = 16'b0000000000000000;
	sram_mem[122885] = 16'b0000000000000000;
	sram_mem[122886] = 16'b0000000000000000;
	sram_mem[122887] = 16'b0000000000000000;
	sram_mem[122888] = 16'b0000000000000000;
	sram_mem[122889] = 16'b0000000000000000;
	sram_mem[122890] = 16'b0000000000000000;
	sram_mem[122891] = 16'b0000000000000000;
	sram_mem[122892] = 16'b0000000000000000;
	sram_mem[122893] = 16'b0000000000000000;
	sram_mem[122894] = 16'b0000000000000000;
	sram_mem[122895] = 16'b0000000000000000;
	sram_mem[122896] = 16'b0000000000000000;
	sram_mem[122897] = 16'b0000000000000000;
	sram_mem[122898] = 16'b0000000000000000;
	sram_mem[122899] = 16'b0000000000000000;
	sram_mem[122900] = 16'b0000000000000000;
	sram_mem[122901] = 16'b0000000000000000;
	sram_mem[122902] = 16'b0000000000000000;
	sram_mem[122903] = 16'b0000000000000000;
	sram_mem[122904] = 16'b0000000000000000;
	sram_mem[122905] = 16'b0000000000000000;
	sram_mem[122906] = 16'b0000000000000000;
	sram_mem[122907] = 16'b0000000000000000;
	sram_mem[122908] = 16'b0000000000000000;
	sram_mem[122909] = 16'b0000000000000000;
	sram_mem[122910] = 16'b0000000000000000;
	sram_mem[122911] = 16'b0000000000000000;
	sram_mem[122912] = 16'b0000000000000000;
	sram_mem[122913] = 16'b0000000000000000;
	sram_mem[122914] = 16'b0000000000000000;
	sram_mem[122915] = 16'b0000000000000000;
	sram_mem[122916] = 16'b0000000000000000;
	sram_mem[122917] = 16'b0000000000000000;
	sram_mem[122918] = 16'b0000000000000000;
	sram_mem[122919] = 16'b0000000000000000;
	sram_mem[122920] = 16'b0000000000000000;
	sram_mem[122921] = 16'b0000000000000000;
	sram_mem[122922] = 16'b0000000000000000;
	sram_mem[122923] = 16'b0000000000000000;
	sram_mem[122924] = 16'b0000000000000000;
	sram_mem[122925] = 16'b0000000000000000;
	sram_mem[122926] = 16'b0000000000000000;
	sram_mem[122927] = 16'b0000000000000000;
	sram_mem[122928] = 16'b0000000000000000;
	sram_mem[122929] = 16'b0000000000000000;
	sram_mem[122930] = 16'b0000000000000000;
	sram_mem[122931] = 16'b0000000000000000;
	sram_mem[122932] = 16'b0000000000000000;
	sram_mem[122933] = 16'b0000000000000000;
	sram_mem[122934] = 16'b0000000000000000;
	sram_mem[122935] = 16'b0000000000000000;
	sram_mem[122936] = 16'b0000000000000000;
	sram_mem[122937] = 16'b0000000000000000;
	sram_mem[122938] = 16'b0000000000000000;
	sram_mem[122939] = 16'b0000000000000000;
	sram_mem[122940] = 16'b0000000000000000;
	sram_mem[122941] = 16'b0000000000000000;
	sram_mem[122942] = 16'b0000000000000000;
	sram_mem[122943] = 16'b0000000000000000;
	sram_mem[122944] = 16'b0000000000000000;
	sram_mem[122945] = 16'b0000000000000000;
	sram_mem[122946] = 16'b0000000000000000;
	sram_mem[122947] = 16'b0000000000000000;
	sram_mem[122948] = 16'b0000000000000000;
	sram_mem[122949] = 16'b0000000000000000;
	sram_mem[122950] = 16'b0000000000000000;
	sram_mem[122951] = 16'b0000000000000000;
	sram_mem[122952] = 16'b0000000000000000;
	sram_mem[122953] = 16'b0000000000000000;
	sram_mem[122954] = 16'b0000000000000000;
	sram_mem[122955] = 16'b0000000000000000;
	sram_mem[122956] = 16'b0000000000000000;
	sram_mem[122957] = 16'b0000000000000000;
	sram_mem[122958] = 16'b0000000000000000;
	sram_mem[122959] = 16'b0000000000000000;
	sram_mem[122960] = 16'b0000000000000000;
	sram_mem[122961] = 16'b0000000000000000;
	sram_mem[122962] = 16'b0000000000000000;
	sram_mem[122963] = 16'b0000000000000000;
	sram_mem[122964] = 16'b0000000000000000;
	sram_mem[122965] = 16'b0000000000000000;
	sram_mem[122966] = 16'b0000000000000000;
	sram_mem[122967] = 16'b0000000000000000;
	sram_mem[122968] = 16'b0000000000000000;
	sram_mem[122969] = 16'b0000000000000000;
	sram_mem[122970] = 16'b0000000000000000;
	sram_mem[122971] = 16'b0000000000000000;
	sram_mem[122972] = 16'b0000000000000000;
	sram_mem[122973] = 16'b0000000000000000;
	sram_mem[122974] = 16'b0000000000000000;
	sram_mem[122975] = 16'b0000000000000000;
	sram_mem[122976] = 16'b0000000000000000;
	sram_mem[122977] = 16'b0000000000000000;
	sram_mem[122978] = 16'b0000000000000000;
	sram_mem[122979] = 16'b0000000000000000;
	sram_mem[122980] = 16'b0000000000000000;
	sram_mem[122981] = 16'b0000000000000000;
	sram_mem[122982] = 16'b0000000000000000;
	sram_mem[122983] = 16'b0000000000000000;
	sram_mem[122984] = 16'b0000000000000000;
	sram_mem[122985] = 16'b0000000000000000;
	sram_mem[122986] = 16'b0000000000000000;
	sram_mem[122987] = 16'b0000000000000000;
	sram_mem[122988] = 16'b0000000000000000;
	sram_mem[122989] = 16'b0000000000000000;
	sram_mem[122990] = 16'b0000000000000000;
	sram_mem[122991] = 16'b0000000000000000;
	sram_mem[122992] = 16'b0000000000000000;
	sram_mem[122993] = 16'b0000000000000000;
	sram_mem[122994] = 16'b0000000000000000;
	sram_mem[122995] = 16'b0000000000000000;
	sram_mem[122996] = 16'b0000000000000000;
	sram_mem[122997] = 16'b0000000000000000;
	sram_mem[122998] = 16'b0000000000000000;
	sram_mem[122999] = 16'b0000000000000000;
	sram_mem[123000] = 16'b0000000000000000;
	sram_mem[123001] = 16'b0000000000000000;
	sram_mem[123002] = 16'b0000000000000000;
	sram_mem[123003] = 16'b0000000000000000;
	sram_mem[123004] = 16'b0000000000000000;
	sram_mem[123005] = 16'b0000000000000000;
	sram_mem[123006] = 16'b0000000000000000;
	sram_mem[123007] = 16'b0000000000000000;
	sram_mem[123008] = 16'b0000000000000000;
	sram_mem[123009] = 16'b0000000000000000;
	sram_mem[123010] = 16'b0000000000000000;
	sram_mem[123011] = 16'b0000000000000000;
	sram_mem[123012] = 16'b0000000000000000;
	sram_mem[123013] = 16'b0000000000000000;
	sram_mem[123014] = 16'b0000000000000000;
	sram_mem[123015] = 16'b0000000000000000;
	sram_mem[123016] = 16'b0000000000000000;
	sram_mem[123017] = 16'b0000000000000000;
	sram_mem[123018] = 16'b0000000000000000;
	sram_mem[123019] = 16'b0000000000000000;
	sram_mem[123020] = 16'b0000000000000000;
	sram_mem[123021] = 16'b0000000000000000;
	sram_mem[123022] = 16'b0000000000000000;
	sram_mem[123023] = 16'b0000000000000000;
	sram_mem[123024] = 16'b0000000000000000;
	sram_mem[123025] = 16'b0000000000000000;
	sram_mem[123026] = 16'b0000000000000000;
	sram_mem[123027] = 16'b0000000000000000;
	sram_mem[123028] = 16'b0000000000000000;
	sram_mem[123029] = 16'b0000000000000000;
	sram_mem[123030] = 16'b0000000000000000;
	sram_mem[123031] = 16'b0000000000000000;
	sram_mem[123032] = 16'b0000000000000000;
	sram_mem[123033] = 16'b0000000000000000;
	sram_mem[123034] = 16'b0000000000000000;
	sram_mem[123035] = 16'b0000000000000000;
	sram_mem[123036] = 16'b0000000000000000;
	sram_mem[123037] = 16'b0000000000000000;
	sram_mem[123038] = 16'b0000000000000000;
	sram_mem[123039] = 16'b0000000000000000;
	sram_mem[123040] = 16'b0000000000000000;
	sram_mem[123041] = 16'b0000000000000000;
	sram_mem[123042] = 16'b0000000000000000;
	sram_mem[123043] = 16'b0000000000000000;
	sram_mem[123044] = 16'b0000000000000000;
	sram_mem[123045] = 16'b0000000000000000;
	sram_mem[123046] = 16'b0000000000000000;
	sram_mem[123047] = 16'b0000000000000000;
	sram_mem[123048] = 16'b0000000000000000;
	sram_mem[123049] = 16'b0000000000000000;
	sram_mem[123050] = 16'b0000000000000000;
	sram_mem[123051] = 16'b0000000000000000;
	sram_mem[123052] = 16'b0000000000000000;
	sram_mem[123053] = 16'b0000000000000000;
	sram_mem[123054] = 16'b0000000000000000;
	sram_mem[123055] = 16'b0000000000000000;
	sram_mem[123056] = 16'b0000000000000000;
	sram_mem[123057] = 16'b0000000000000000;
	sram_mem[123058] = 16'b0000000000000000;
	sram_mem[123059] = 16'b0000000000000000;
	sram_mem[123060] = 16'b0000000000000000;
	sram_mem[123061] = 16'b0000000000000000;
	sram_mem[123062] = 16'b0000000000000000;
	sram_mem[123063] = 16'b0000000000000000;
	sram_mem[123064] = 16'b0000000000000000;
	sram_mem[123065] = 16'b0000000000000000;
	sram_mem[123066] = 16'b0000000000000000;
	sram_mem[123067] = 16'b0000000000000000;
	sram_mem[123068] = 16'b0000000000000000;
	sram_mem[123069] = 16'b0000000000000000;
	sram_mem[123070] = 16'b0000000000000000;
	sram_mem[123071] = 16'b0000000000000000;
	sram_mem[123072] = 16'b0000000000000000;
	sram_mem[123073] = 16'b0000000000000000;
	sram_mem[123074] = 16'b0000000000000000;
	sram_mem[123075] = 16'b0000000000000000;
	sram_mem[123076] = 16'b0000000000000000;
	sram_mem[123077] = 16'b0000000000000000;
	sram_mem[123078] = 16'b0000000000000000;
	sram_mem[123079] = 16'b0000000000000000;
	sram_mem[123080] = 16'b0000000000000000;
	sram_mem[123081] = 16'b0000000000000000;
	sram_mem[123082] = 16'b0000000000000000;
	sram_mem[123083] = 16'b0000000000000000;
	sram_mem[123084] = 16'b0000000000000000;
	sram_mem[123085] = 16'b0000000000000000;
	sram_mem[123086] = 16'b0000000000000000;
	sram_mem[123087] = 16'b0000000000000000;
	sram_mem[123088] = 16'b0000000000000000;
	sram_mem[123089] = 16'b0000000000000000;
	sram_mem[123090] = 16'b0000000000000000;
	sram_mem[123091] = 16'b0000000000000000;
	sram_mem[123092] = 16'b0000000000000000;
	sram_mem[123093] = 16'b0000000000000000;
	sram_mem[123094] = 16'b0000000000000000;
	sram_mem[123095] = 16'b0000000000000000;
	sram_mem[123096] = 16'b0000000000000000;
	sram_mem[123097] = 16'b0000000000000000;
	sram_mem[123098] = 16'b0000000000000000;
	sram_mem[123099] = 16'b0000000000000000;
	sram_mem[123100] = 16'b0000000000000000;
	sram_mem[123101] = 16'b0000000000000000;
	sram_mem[123102] = 16'b0000000000000000;
	sram_mem[123103] = 16'b0000000000000000;
	sram_mem[123104] = 16'b0000000000000000;
	sram_mem[123105] = 16'b0000000000000000;
	sram_mem[123106] = 16'b0000000000000000;
	sram_mem[123107] = 16'b0000000000000000;
	sram_mem[123108] = 16'b0000000000000000;
	sram_mem[123109] = 16'b0000000000000000;
	sram_mem[123110] = 16'b0000000000000000;
	sram_mem[123111] = 16'b0000000000000000;
	sram_mem[123112] = 16'b0000000000000000;
	sram_mem[123113] = 16'b0000000000000000;
	sram_mem[123114] = 16'b0000000000000000;
	sram_mem[123115] = 16'b0000000000000000;
	sram_mem[123116] = 16'b0000000000000000;
	sram_mem[123117] = 16'b0000000000000000;
	sram_mem[123118] = 16'b0000000000000000;
	sram_mem[123119] = 16'b0000000000000000;
	sram_mem[123120] = 16'b0000000000000000;
	sram_mem[123121] = 16'b0000000000000000;
	sram_mem[123122] = 16'b0000000000000000;
	sram_mem[123123] = 16'b0000000000000000;
	sram_mem[123124] = 16'b0000000000000000;
	sram_mem[123125] = 16'b0000000000000000;
	sram_mem[123126] = 16'b0000000000000000;
	sram_mem[123127] = 16'b0000000000000000;
	sram_mem[123128] = 16'b0000000000000000;
	sram_mem[123129] = 16'b0000000000000000;
	sram_mem[123130] = 16'b0000000000000000;
	sram_mem[123131] = 16'b0000000000000000;
	sram_mem[123132] = 16'b0000000000000000;
	sram_mem[123133] = 16'b0000000000000000;
	sram_mem[123134] = 16'b0000000000000000;
	sram_mem[123135] = 16'b0000000000000000;
	sram_mem[123136] = 16'b0000000000000000;
	sram_mem[123137] = 16'b0000000000000000;
	sram_mem[123138] = 16'b0000000000000000;
	sram_mem[123139] = 16'b0000000000000000;
	sram_mem[123140] = 16'b0000000000000000;
	sram_mem[123141] = 16'b0000000000000000;
	sram_mem[123142] = 16'b0000000000000000;
	sram_mem[123143] = 16'b0000000000000000;
	sram_mem[123144] = 16'b0000000000000000;
	sram_mem[123145] = 16'b0000000000000000;
	sram_mem[123146] = 16'b0000000000000000;
	sram_mem[123147] = 16'b0000000000000000;
	sram_mem[123148] = 16'b0000000000000000;
	sram_mem[123149] = 16'b0000000000000000;
	sram_mem[123150] = 16'b0000000000000000;
	sram_mem[123151] = 16'b0000000000000000;
	sram_mem[123152] = 16'b0000000000000000;
	sram_mem[123153] = 16'b0000000000000000;
	sram_mem[123154] = 16'b0000000000000000;
	sram_mem[123155] = 16'b0000000000000000;
	sram_mem[123156] = 16'b0000000000000000;
	sram_mem[123157] = 16'b0000000000000000;
	sram_mem[123158] = 16'b0000000000000000;
	sram_mem[123159] = 16'b0000000000000000;
	sram_mem[123160] = 16'b0000000000000000;
	sram_mem[123161] = 16'b0000000000000000;
	sram_mem[123162] = 16'b0000000000000000;
	sram_mem[123163] = 16'b0000000000000000;
	sram_mem[123164] = 16'b0000000000000000;
	sram_mem[123165] = 16'b0000000000000000;
	sram_mem[123166] = 16'b0000000000000000;
	sram_mem[123167] = 16'b0000000000000000;
	sram_mem[123168] = 16'b0000000000000000;
	sram_mem[123169] = 16'b0000000000000000;
	sram_mem[123170] = 16'b0000000000000000;
	sram_mem[123171] = 16'b0000000000000000;
	sram_mem[123172] = 16'b0000000000000000;
	sram_mem[123173] = 16'b0000000000000000;
	sram_mem[123174] = 16'b0000000000000000;
	sram_mem[123175] = 16'b0000000000000000;
	sram_mem[123176] = 16'b0000000000000000;
	sram_mem[123177] = 16'b0000000000000000;
	sram_mem[123178] = 16'b0000000000000000;
	sram_mem[123179] = 16'b0000000000000000;
	sram_mem[123180] = 16'b0000000000000000;
	sram_mem[123181] = 16'b0000000000000000;
	sram_mem[123182] = 16'b0000000000000000;
	sram_mem[123183] = 16'b0000000000000000;
	sram_mem[123184] = 16'b0000000000000000;
	sram_mem[123185] = 16'b0000000000000000;
	sram_mem[123186] = 16'b0000000000000000;
	sram_mem[123187] = 16'b0000000000000000;
	sram_mem[123188] = 16'b0000000000000000;
	sram_mem[123189] = 16'b0000000000000000;
	sram_mem[123190] = 16'b0000000000000000;
	sram_mem[123191] = 16'b0000000000000000;
	sram_mem[123192] = 16'b0000000000000000;
	sram_mem[123193] = 16'b0000000000000000;
	sram_mem[123194] = 16'b0000000000000000;
	sram_mem[123195] = 16'b0000000000000000;
	sram_mem[123196] = 16'b0000000000000000;
	sram_mem[123197] = 16'b0000000000000000;
	sram_mem[123198] = 16'b0000000000000000;
	sram_mem[123199] = 16'b0000000000000000;
	sram_mem[123200] = 16'b0000000000000000;
	sram_mem[123201] = 16'b0000000000000000;
	sram_mem[123202] = 16'b0000000000000000;
	sram_mem[123203] = 16'b0000000000000000;
	sram_mem[123204] = 16'b0000000000000000;
	sram_mem[123205] = 16'b0000000000000000;
	sram_mem[123206] = 16'b0000000000000000;
	sram_mem[123207] = 16'b0000000000000000;
	sram_mem[123208] = 16'b0000000000000000;
	sram_mem[123209] = 16'b0000000000000000;
	sram_mem[123210] = 16'b0000000000000000;
	sram_mem[123211] = 16'b0000000000000000;
	sram_mem[123212] = 16'b0000000000000000;
	sram_mem[123213] = 16'b0000000000000000;
	sram_mem[123214] = 16'b0000000000000000;
	sram_mem[123215] = 16'b0000000000000000;
	sram_mem[123216] = 16'b0000000000000000;
	sram_mem[123217] = 16'b0000000000000000;
	sram_mem[123218] = 16'b0000000000000000;
	sram_mem[123219] = 16'b0000000000000000;
	sram_mem[123220] = 16'b0000000000000000;
	sram_mem[123221] = 16'b0000000000000000;
	sram_mem[123222] = 16'b0000000000000000;
	sram_mem[123223] = 16'b0000000000000000;
	sram_mem[123224] = 16'b0000000000000000;
	sram_mem[123225] = 16'b0000000000000000;
	sram_mem[123226] = 16'b0000000000000000;
	sram_mem[123227] = 16'b0000000000000000;
	sram_mem[123228] = 16'b0000000000000000;
	sram_mem[123229] = 16'b0000000000000000;
	sram_mem[123230] = 16'b0000000000000000;
	sram_mem[123231] = 16'b0000000000000000;
	sram_mem[123232] = 16'b0000000000000000;
	sram_mem[123233] = 16'b0000000000000000;
	sram_mem[123234] = 16'b0000000000000000;
	sram_mem[123235] = 16'b0000000000000000;
	sram_mem[123236] = 16'b0000000000000000;
	sram_mem[123237] = 16'b0000000000000000;
	sram_mem[123238] = 16'b0000000000000000;
	sram_mem[123239] = 16'b0000000000000000;
	sram_mem[123240] = 16'b0000000000000000;
	sram_mem[123241] = 16'b0000000000000000;
	sram_mem[123242] = 16'b0000000000000000;
	sram_mem[123243] = 16'b0000000000000000;
	sram_mem[123244] = 16'b0000000000000000;
	sram_mem[123245] = 16'b0000000000000000;
	sram_mem[123246] = 16'b0000000000000000;
	sram_mem[123247] = 16'b0000000000000000;
	sram_mem[123248] = 16'b0000000000000000;
	sram_mem[123249] = 16'b0000000000000000;
	sram_mem[123250] = 16'b0000000000000000;
	sram_mem[123251] = 16'b0000000000000000;
	sram_mem[123252] = 16'b0000000000000000;
	sram_mem[123253] = 16'b0000000000000000;
	sram_mem[123254] = 16'b0000000000000000;
	sram_mem[123255] = 16'b0000000000000000;
	sram_mem[123256] = 16'b0000000000000000;
	sram_mem[123257] = 16'b0000000000000000;
	sram_mem[123258] = 16'b0000000000000000;
	sram_mem[123259] = 16'b0000000000000000;
	sram_mem[123260] = 16'b0000000000000000;
	sram_mem[123261] = 16'b0000000000000000;
	sram_mem[123262] = 16'b0000000000000000;
	sram_mem[123263] = 16'b0000000000000000;
	sram_mem[123264] = 16'b0000000000000000;
	sram_mem[123265] = 16'b0000000000000000;
	sram_mem[123266] = 16'b0000000000000000;
	sram_mem[123267] = 16'b0000000000000000;
	sram_mem[123268] = 16'b0000000000000000;
	sram_mem[123269] = 16'b0000000000000000;
	sram_mem[123270] = 16'b0000000000000000;
	sram_mem[123271] = 16'b0000000000000000;
	sram_mem[123272] = 16'b0000000000000000;
	sram_mem[123273] = 16'b0000000000000000;
	sram_mem[123274] = 16'b0000000000000000;
	sram_mem[123275] = 16'b0000000000000000;
	sram_mem[123276] = 16'b0000000000000000;
	sram_mem[123277] = 16'b0000000000000000;
	sram_mem[123278] = 16'b0000000000000000;
	sram_mem[123279] = 16'b0000000000000000;
	sram_mem[123280] = 16'b0000000000000000;
	sram_mem[123281] = 16'b0000000000000000;
	sram_mem[123282] = 16'b0000000000000000;
	sram_mem[123283] = 16'b0000000000000000;
	sram_mem[123284] = 16'b0000000000000000;
	sram_mem[123285] = 16'b0000000000000000;
	sram_mem[123286] = 16'b0000000000000000;
	sram_mem[123287] = 16'b0000000000000000;
	sram_mem[123288] = 16'b0000000000000000;
	sram_mem[123289] = 16'b0000000000000000;
	sram_mem[123290] = 16'b0000000000000000;
	sram_mem[123291] = 16'b0000000000000000;
	sram_mem[123292] = 16'b0000000000000000;
	sram_mem[123293] = 16'b0000000000000000;
	sram_mem[123294] = 16'b0000000000000000;
	sram_mem[123295] = 16'b0000000000000000;
	sram_mem[123296] = 16'b0000000000000000;
	sram_mem[123297] = 16'b0000000000000000;
	sram_mem[123298] = 16'b0000000000000000;
	sram_mem[123299] = 16'b0000000000000000;
	sram_mem[123300] = 16'b0000000000000000;
	sram_mem[123301] = 16'b0000000000000000;
	sram_mem[123302] = 16'b0000000000000000;
	sram_mem[123303] = 16'b0000000000000000;
	sram_mem[123304] = 16'b0000000000000000;
	sram_mem[123305] = 16'b0000000000000000;
	sram_mem[123306] = 16'b0000000000000000;
	sram_mem[123307] = 16'b0000000000000000;
	sram_mem[123308] = 16'b0000000000000000;
	sram_mem[123309] = 16'b0000000000000000;
	sram_mem[123310] = 16'b0000000000000000;
	sram_mem[123311] = 16'b0000000000000000;
	sram_mem[123312] = 16'b0000000000000000;
	sram_mem[123313] = 16'b0000000000000000;
	sram_mem[123314] = 16'b0000000000000000;
	sram_mem[123315] = 16'b0000000000000000;
	sram_mem[123316] = 16'b0000000000000000;
	sram_mem[123317] = 16'b0000000000000000;
	sram_mem[123318] = 16'b0000000000000000;
	sram_mem[123319] = 16'b0000000000000000;
	sram_mem[123320] = 16'b0000000000000000;
	sram_mem[123321] = 16'b0000000000000000;
	sram_mem[123322] = 16'b0000000000000000;
	sram_mem[123323] = 16'b0000000000000000;
	sram_mem[123324] = 16'b0000000000000000;
	sram_mem[123325] = 16'b0000000000000000;
	sram_mem[123326] = 16'b0000000000000000;
	sram_mem[123327] = 16'b0000000000000000;
	sram_mem[123328] = 16'b0000000000000000;
	sram_mem[123329] = 16'b0000000000000000;
	sram_mem[123330] = 16'b0000000000000000;
	sram_mem[123331] = 16'b0000000000000000;
	sram_mem[123332] = 16'b0000000000000000;
	sram_mem[123333] = 16'b0000000000000000;
	sram_mem[123334] = 16'b0000000000000000;
	sram_mem[123335] = 16'b0000000000000000;
	sram_mem[123336] = 16'b0000000000000000;
	sram_mem[123337] = 16'b0000000000000000;
	sram_mem[123338] = 16'b0000000000000000;
	sram_mem[123339] = 16'b0000000000000000;
	sram_mem[123340] = 16'b0000000000000000;
	sram_mem[123341] = 16'b0000000000000000;
	sram_mem[123342] = 16'b0000000000000000;
	sram_mem[123343] = 16'b0000000000000000;
	sram_mem[123344] = 16'b0000000000000000;
	sram_mem[123345] = 16'b0000000000000000;
	sram_mem[123346] = 16'b0000000000000000;
	sram_mem[123347] = 16'b0000000000000000;
	sram_mem[123348] = 16'b0000000000000000;
	sram_mem[123349] = 16'b0000000000000000;
	sram_mem[123350] = 16'b0000000000000000;
	sram_mem[123351] = 16'b0000000000000000;
	sram_mem[123352] = 16'b0000000000000000;
	sram_mem[123353] = 16'b0000000000000000;
	sram_mem[123354] = 16'b0000000000000000;
	sram_mem[123355] = 16'b0000000000000000;
	sram_mem[123356] = 16'b0000000000000000;
	sram_mem[123357] = 16'b0000000000000000;
	sram_mem[123358] = 16'b0000000000000000;
	sram_mem[123359] = 16'b0000000000000000;
	sram_mem[123360] = 16'b0000000000000000;
	sram_mem[123361] = 16'b0000000000000000;
	sram_mem[123362] = 16'b0000000000000000;
	sram_mem[123363] = 16'b0000000000000000;
	sram_mem[123364] = 16'b0000000000000000;
	sram_mem[123365] = 16'b0000000000000000;
	sram_mem[123366] = 16'b0000000000000000;
	sram_mem[123367] = 16'b0000000000000000;
	sram_mem[123368] = 16'b0000000000000000;
	sram_mem[123369] = 16'b0000000000000000;
	sram_mem[123370] = 16'b0000000000000000;
	sram_mem[123371] = 16'b0000000000000000;
	sram_mem[123372] = 16'b0000000000000000;
	sram_mem[123373] = 16'b0000000000000000;
	sram_mem[123374] = 16'b0000000000000000;
	sram_mem[123375] = 16'b0000000000000000;
	sram_mem[123376] = 16'b0000000000000000;
	sram_mem[123377] = 16'b0000000000000000;
	sram_mem[123378] = 16'b0000000000000000;
	sram_mem[123379] = 16'b0000000000000000;
	sram_mem[123380] = 16'b0000000000000000;
	sram_mem[123381] = 16'b0000000000000000;
	sram_mem[123382] = 16'b0000000000000000;
	sram_mem[123383] = 16'b0000000000000000;
	sram_mem[123384] = 16'b0000000000000000;
	sram_mem[123385] = 16'b0000000000000000;
	sram_mem[123386] = 16'b0000000000000000;
	sram_mem[123387] = 16'b0000000000000000;
	sram_mem[123388] = 16'b0000000000000000;
	sram_mem[123389] = 16'b0000000000000000;
	sram_mem[123390] = 16'b0000000000000000;
	sram_mem[123391] = 16'b0000000000000000;
	sram_mem[123392] = 16'b0000000000000000;
	sram_mem[123393] = 16'b0000000000000000;
	sram_mem[123394] = 16'b0000000000000000;
	sram_mem[123395] = 16'b0000000000000000;
	sram_mem[123396] = 16'b0000000000000000;
	sram_mem[123397] = 16'b0000000000000000;
	sram_mem[123398] = 16'b0000000000000000;
	sram_mem[123399] = 16'b0000000000000000;
	sram_mem[123400] = 16'b0000000000000000;
	sram_mem[123401] = 16'b0000000000000000;
	sram_mem[123402] = 16'b0000000000000000;
	sram_mem[123403] = 16'b0000000000000000;
	sram_mem[123404] = 16'b0000000000000000;
	sram_mem[123405] = 16'b0000000000000000;
	sram_mem[123406] = 16'b0000000000000000;
	sram_mem[123407] = 16'b0000000000000000;
	sram_mem[123408] = 16'b0000000000000000;
	sram_mem[123409] = 16'b0000000000000000;
	sram_mem[123410] = 16'b0000000000000000;
	sram_mem[123411] = 16'b0000000000000000;
	sram_mem[123412] = 16'b0000000000000000;
	sram_mem[123413] = 16'b0000000000000000;
	sram_mem[123414] = 16'b0000000000000000;
	sram_mem[123415] = 16'b0000000000000000;
	sram_mem[123416] = 16'b0000000000000000;
	sram_mem[123417] = 16'b0000000000000000;
	sram_mem[123418] = 16'b0000000000000000;
	sram_mem[123419] = 16'b0000000000000000;
	sram_mem[123420] = 16'b0000000000000000;
	sram_mem[123421] = 16'b0000000000000000;
	sram_mem[123422] = 16'b0000000000000000;
	sram_mem[123423] = 16'b0000000000000000;
	sram_mem[123424] = 16'b0000000000000000;
	sram_mem[123425] = 16'b0000000000000000;
	sram_mem[123426] = 16'b0000000000000000;
	sram_mem[123427] = 16'b0000000000000000;
	sram_mem[123428] = 16'b0000000000000000;
	sram_mem[123429] = 16'b0000000000000000;
	sram_mem[123430] = 16'b0000000000000000;
	sram_mem[123431] = 16'b0000000000000000;
	sram_mem[123432] = 16'b0000000000000000;
	sram_mem[123433] = 16'b0000000000000000;
	sram_mem[123434] = 16'b0000000000000000;
	sram_mem[123435] = 16'b0000000000000000;
	sram_mem[123436] = 16'b0000000000000000;
	sram_mem[123437] = 16'b0000000000000000;
	sram_mem[123438] = 16'b0000000000000000;
	sram_mem[123439] = 16'b0000000000000000;
	sram_mem[123440] = 16'b0000000000000000;
	sram_mem[123441] = 16'b0000000000000000;
	sram_mem[123442] = 16'b0000000000000000;
	sram_mem[123443] = 16'b0000000000000000;
	sram_mem[123444] = 16'b0000000000000000;
	sram_mem[123445] = 16'b0000000000000000;
	sram_mem[123446] = 16'b0000000000000000;
	sram_mem[123447] = 16'b0000000000000000;
	sram_mem[123448] = 16'b0000000000000000;
	sram_mem[123449] = 16'b0000000000000000;
	sram_mem[123450] = 16'b0000000000000000;
	sram_mem[123451] = 16'b0000000000000000;
	sram_mem[123452] = 16'b0000000000000000;
	sram_mem[123453] = 16'b0000000000000000;
	sram_mem[123454] = 16'b0000000000000000;
	sram_mem[123455] = 16'b0000000000000000;
	sram_mem[123456] = 16'b0000000000000000;
	sram_mem[123457] = 16'b0000000000000000;
	sram_mem[123458] = 16'b0000000000000000;
	sram_mem[123459] = 16'b0000000000000000;
	sram_mem[123460] = 16'b0000000000000000;
	sram_mem[123461] = 16'b0000000000000000;
	sram_mem[123462] = 16'b0000000000000000;
	sram_mem[123463] = 16'b0000000000000000;
	sram_mem[123464] = 16'b0000000000000000;
	sram_mem[123465] = 16'b0000000000000000;
	sram_mem[123466] = 16'b0000000000000000;
	sram_mem[123467] = 16'b0000000000000000;
	sram_mem[123468] = 16'b0000000000000000;
	sram_mem[123469] = 16'b0000000000000000;
	sram_mem[123470] = 16'b0000000000000000;
	sram_mem[123471] = 16'b0000000000000000;
	sram_mem[123472] = 16'b0000000000000000;
	sram_mem[123473] = 16'b0000000000000000;
	sram_mem[123474] = 16'b0000000000000000;
	sram_mem[123475] = 16'b0000000000000000;
	sram_mem[123476] = 16'b0000000000000000;
	sram_mem[123477] = 16'b0000000000000000;
	sram_mem[123478] = 16'b0000000000000000;
	sram_mem[123479] = 16'b0000000000000000;
	sram_mem[123480] = 16'b0000000000000000;
	sram_mem[123481] = 16'b0000000000000000;
	sram_mem[123482] = 16'b0000000000000000;
	sram_mem[123483] = 16'b0000000000000000;
	sram_mem[123484] = 16'b0000000000000000;
	sram_mem[123485] = 16'b0000000000000000;
	sram_mem[123486] = 16'b0000000000000000;
	sram_mem[123487] = 16'b0000000000000000;
	sram_mem[123488] = 16'b0000000000000000;
	sram_mem[123489] = 16'b0000000000000000;
	sram_mem[123490] = 16'b0000000000000000;
	sram_mem[123491] = 16'b0000000000000000;
	sram_mem[123492] = 16'b0000000000000000;
	sram_mem[123493] = 16'b0000000000000000;
	sram_mem[123494] = 16'b0000000000000000;
	sram_mem[123495] = 16'b0000000000000000;
	sram_mem[123496] = 16'b0000000000000000;
	sram_mem[123497] = 16'b0000000000000000;
	sram_mem[123498] = 16'b0000000000000000;
	sram_mem[123499] = 16'b0000000000000000;
	sram_mem[123500] = 16'b0000000000000000;
	sram_mem[123501] = 16'b0000000000000000;
	sram_mem[123502] = 16'b0000000000000000;
	sram_mem[123503] = 16'b0000000000000000;
	sram_mem[123504] = 16'b0000000000000000;
	sram_mem[123505] = 16'b0000000000000000;
	sram_mem[123506] = 16'b0000000000000000;
	sram_mem[123507] = 16'b0000000000000000;
	sram_mem[123508] = 16'b0000000000000000;
	sram_mem[123509] = 16'b0000000000000000;
	sram_mem[123510] = 16'b0000000000000000;
	sram_mem[123511] = 16'b0000000000000000;
	sram_mem[123512] = 16'b0000000000000000;
	sram_mem[123513] = 16'b0000000000000000;
	sram_mem[123514] = 16'b0000000000000000;
	sram_mem[123515] = 16'b0000000000000000;
	sram_mem[123516] = 16'b0000000000000000;
	sram_mem[123517] = 16'b0000000000000000;
	sram_mem[123518] = 16'b0000000000000000;
	sram_mem[123519] = 16'b0000000000000000;
	sram_mem[123520] = 16'b0000000000000000;
	sram_mem[123521] = 16'b0000000000000000;
	sram_mem[123522] = 16'b0000000000000000;
	sram_mem[123523] = 16'b0000000000000000;
	sram_mem[123524] = 16'b0000000000000000;
	sram_mem[123525] = 16'b0000000000000000;
	sram_mem[123526] = 16'b0000000000000000;
	sram_mem[123527] = 16'b0000000000000000;
	sram_mem[123528] = 16'b0000000000000000;
	sram_mem[123529] = 16'b0000000000000000;
	sram_mem[123530] = 16'b0000000000000000;
	sram_mem[123531] = 16'b0000000000000000;
	sram_mem[123532] = 16'b0000000000000000;
	sram_mem[123533] = 16'b0000000000000000;
	sram_mem[123534] = 16'b0000000000000000;
	sram_mem[123535] = 16'b0000000000000000;
	sram_mem[123536] = 16'b0000000000000000;
	sram_mem[123537] = 16'b0000000000000000;
	sram_mem[123538] = 16'b0000000000000000;
	sram_mem[123539] = 16'b0000000000000000;
	sram_mem[123540] = 16'b0000000000000000;
	sram_mem[123541] = 16'b0000000000000000;
	sram_mem[123542] = 16'b0000000000000000;
	sram_mem[123543] = 16'b0000000000000000;
	sram_mem[123544] = 16'b0000000000000000;
	sram_mem[123545] = 16'b0000000000000000;
	sram_mem[123546] = 16'b0000000000000000;
	sram_mem[123547] = 16'b0000000000000000;
	sram_mem[123548] = 16'b0000000000000000;
	sram_mem[123549] = 16'b0000000000000000;
	sram_mem[123550] = 16'b0000000000000000;
	sram_mem[123551] = 16'b0000000000000000;
	sram_mem[123552] = 16'b0000000000000000;
	sram_mem[123553] = 16'b0000000000000000;
	sram_mem[123554] = 16'b0000000000000000;
	sram_mem[123555] = 16'b0000000000000000;
	sram_mem[123556] = 16'b0000000000000000;
	sram_mem[123557] = 16'b0000000000000000;
	sram_mem[123558] = 16'b0000000000000000;
	sram_mem[123559] = 16'b0000000000000000;
	sram_mem[123560] = 16'b0000000000000000;
	sram_mem[123561] = 16'b0000000000000000;
	sram_mem[123562] = 16'b0000000000000000;
	sram_mem[123563] = 16'b0000000000000000;
	sram_mem[123564] = 16'b0000000000000000;
	sram_mem[123565] = 16'b0000000000000000;
	sram_mem[123566] = 16'b0000000000000000;
	sram_mem[123567] = 16'b0000000000000000;
	sram_mem[123568] = 16'b0000000000000000;
	sram_mem[123569] = 16'b0000000000000000;
	sram_mem[123570] = 16'b0000000000000000;
	sram_mem[123571] = 16'b0000000000000000;
	sram_mem[123572] = 16'b0000000000000000;
	sram_mem[123573] = 16'b0000000000000000;
	sram_mem[123574] = 16'b0000000000000000;
	sram_mem[123575] = 16'b0000000000000000;
	sram_mem[123576] = 16'b0000000000000000;
	sram_mem[123577] = 16'b0000000000000000;
	sram_mem[123578] = 16'b0000000000000000;
	sram_mem[123579] = 16'b0000000000000000;
	sram_mem[123580] = 16'b0000000000000000;
	sram_mem[123581] = 16'b0000000000000000;
	sram_mem[123582] = 16'b0000000000000000;
	sram_mem[123583] = 16'b0000000000000000;
	sram_mem[123584] = 16'b0000000000000000;
	sram_mem[123585] = 16'b0000000000000000;
	sram_mem[123586] = 16'b0000000000000000;
	sram_mem[123587] = 16'b0000000000000000;
	sram_mem[123588] = 16'b0000000000000000;
	sram_mem[123589] = 16'b0000000000000000;
	sram_mem[123590] = 16'b0000000000000000;
	sram_mem[123591] = 16'b0000000000000000;
	sram_mem[123592] = 16'b0000000000000000;
	sram_mem[123593] = 16'b0000000000000000;
	sram_mem[123594] = 16'b0000000000000000;
	sram_mem[123595] = 16'b0000000000000000;
	sram_mem[123596] = 16'b0000000000000000;
	sram_mem[123597] = 16'b0000000000000000;
	sram_mem[123598] = 16'b0000000000000000;
	sram_mem[123599] = 16'b0000000000000000;
	sram_mem[123600] = 16'b0000000000000000;
	sram_mem[123601] = 16'b0000000000000000;
	sram_mem[123602] = 16'b0000000000000000;
	sram_mem[123603] = 16'b0000000000000000;
	sram_mem[123604] = 16'b0000000000000000;
	sram_mem[123605] = 16'b0000000000000000;
	sram_mem[123606] = 16'b0000000000000000;
	sram_mem[123607] = 16'b0000000000000000;
	sram_mem[123608] = 16'b0000000000000000;
	sram_mem[123609] = 16'b0000000000000000;
	sram_mem[123610] = 16'b0000000000000000;
	sram_mem[123611] = 16'b0000000000000000;
	sram_mem[123612] = 16'b0000000000000000;
	sram_mem[123613] = 16'b0000000000000000;
	sram_mem[123614] = 16'b0000000000000000;
	sram_mem[123615] = 16'b0000000000000000;
	sram_mem[123616] = 16'b0000000000000000;
	sram_mem[123617] = 16'b0000000000000000;
	sram_mem[123618] = 16'b0000000000000000;
	sram_mem[123619] = 16'b0000000000000000;
	sram_mem[123620] = 16'b0000000000000000;
	sram_mem[123621] = 16'b0000000000000000;
	sram_mem[123622] = 16'b0000000000000000;
	sram_mem[123623] = 16'b0000000000000000;
	sram_mem[123624] = 16'b0000000000000000;
	sram_mem[123625] = 16'b0000000000000000;
	sram_mem[123626] = 16'b0000000000000000;
	sram_mem[123627] = 16'b0000000000000000;
	sram_mem[123628] = 16'b0000000000000000;
	sram_mem[123629] = 16'b0000000000000000;
	sram_mem[123630] = 16'b0000000000000000;
	sram_mem[123631] = 16'b0000000000000000;
	sram_mem[123632] = 16'b0000000000000000;
	sram_mem[123633] = 16'b0000000000000000;
	sram_mem[123634] = 16'b0000000000000000;
	sram_mem[123635] = 16'b0000000000000000;
	sram_mem[123636] = 16'b0000000000000000;
	sram_mem[123637] = 16'b0000000000000000;
	sram_mem[123638] = 16'b0000000000000000;
	sram_mem[123639] = 16'b0000000000000000;
	sram_mem[123640] = 16'b0000000000000000;
	sram_mem[123641] = 16'b0000000000000000;
	sram_mem[123642] = 16'b0000000000000000;
	sram_mem[123643] = 16'b0000000000000000;
	sram_mem[123644] = 16'b0000000000000000;
	sram_mem[123645] = 16'b0000000000000000;
	sram_mem[123646] = 16'b0000000000000000;
	sram_mem[123647] = 16'b0000000000000000;
	sram_mem[123648] = 16'b0000000000000000;
	sram_mem[123649] = 16'b0000000000000000;
	sram_mem[123650] = 16'b0000000000000000;
	sram_mem[123651] = 16'b0000000000000000;
	sram_mem[123652] = 16'b0000000000000000;
	sram_mem[123653] = 16'b0000000000000000;
	sram_mem[123654] = 16'b0000000000000000;
	sram_mem[123655] = 16'b0000000000000000;
	sram_mem[123656] = 16'b0000000000000000;
	sram_mem[123657] = 16'b0000000000000000;
	sram_mem[123658] = 16'b0000000000000000;
	sram_mem[123659] = 16'b0000000000000000;
	sram_mem[123660] = 16'b0000000000000000;
	sram_mem[123661] = 16'b0000000000000000;
	sram_mem[123662] = 16'b0000000000000000;
	sram_mem[123663] = 16'b0000000000000000;
	sram_mem[123664] = 16'b0000000000000000;
	sram_mem[123665] = 16'b0000000000000000;
	sram_mem[123666] = 16'b0000000000000000;
	sram_mem[123667] = 16'b0000000000000000;
	sram_mem[123668] = 16'b0000000000000000;
	sram_mem[123669] = 16'b0000000000000000;
	sram_mem[123670] = 16'b0000000000000000;
	sram_mem[123671] = 16'b0000000000000000;
	sram_mem[123672] = 16'b0000000000000000;
	sram_mem[123673] = 16'b0000000000000000;
	sram_mem[123674] = 16'b0000000000000000;
	sram_mem[123675] = 16'b0000000000000000;
	sram_mem[123676] = 16'b0000000000000000;
	sram_mem[123677] = 16'b0000000000000000;
	sram_mem[123678] = 16'b0000000000000000;
	sram_mem[123679] = 16'b0000000000000000;
	sram_mem[123680] = 16'b0000000000000000;
	sram_mem[123681] = 16'b0000000000000000;
	sram_mem[123682] = 16'b0000000000000000;
	sram_mem[123683] = 16'b0000000000000000;
	sram_mem[123684] = 16'b0000000000000000;
	sram_mem[123685] = 16'b0000000000000000;
	sram_mem[123686] = 16'b0000000000000000;
	sram_mem[123687] = 16'b0000000000000000;
	sram_mem[123688] = 16'b0000000000000000;
	sram_mem[123689] = 16'b0000000000000000;
	sram_mem[123690] = 16'b0000000000000000;
	sram_mem[123691] = 16'b0000000000000000;
	sram_mem[123692] = 16'b0000000000000000;
	sram_mem[123693] = 16'b0000000000000000;
	sram_mem[123694] = 16'b0000000000000000;
	sram_mem[123695] = 16'b0000000000000000;
	sram_mem[123696] = 16'b0000000000000000;
	sram_mem[123697] = 16'b0000000000000000;
	sram_mem[123698] = 16'b0000000000000000;
	sram_mem[123699] = 16'b0000000000000000;
	sram_mem[123700] = 16'b0000000000000000;
	sram_mem[123701] = 16'b0000000000000000;
	sram_mem[123702] = 16'b0000000000000000;
	sram_mem[123703] = 16'b0000000000000000;
	sram_mem[123704] = 16'b0000000000000000;
	sram_mem[123705] = 16'b0000000000000000;
	sram_mem[123706] = 16'b0000000000000000;
	sram_mem[123707] = 16'b0000000000000000;
	sram_mem[123708] = 16'b0000000000000000;
	sram_mem[123709] = 16'b0000000000000000;
	sram_mem[123710] = 16'b0000000000000000;
	sram_mem[123711] = 16'b0000000000000000;
	sram_mem[123712] = 16'b0000000000000000;
	sram_mem[123713] = 16'b0000000000000000;
	sram_mem[123714] = 16'b0000000000000000;
	sram_mem[123715] = 16'b0000000000000000;
	sram_mem[123716] = 16'b0000000000000000;
	sram_mem[123717] = 16'b0000000000000000;
	sram_mem[123718] = 16'b0000000000000000;
	sram_mem[123719] = 16'b0000000000000000;
	sram_mem[123720] = 16'b0000000000000000;
	sram_mem[123721] = 16'b0000000000000000;
	sram_mem[123722] = 16'b0000000000000000;
	sram_mem[123723] = 16'b0000000000000000;
	sram_mem[123724] = 16'b0000000000000000;
	sram_mem[123725] = 16'b0000000000000000;
	sram_mem[123726] = 16'b0000000000000000;
	sram_mem[123727] = 16'b0000000000000000;
	sram_mem[123728] = 16'b0000000000000000;
	sram_mem[123729] = 16'b0000000000000000;
	sram_mem[123730] = 16'b0000000000000000;
	sram_mem[123731] = 16'b0000000000000000;
	sram_mem[123732] = 16'b0000000000000000;
	sram_mem[123733] = 16'b0000000000000000;
	sram_mem[123734] = 16'b0000000000000000;
	sram_mem[123735] = 16'b0000000000000000;
	sram_mem[123736] = 16'b0000000000000000;
	sram_mem[123737] = 16'b0000000000000000;
	sram_mem[123738] = 16'b0000000000000000;
	sram_mem[123739] = 16'b0000000000000000;
	sram_mem[123740] = 16'b0000000000000000;
	sram_mem[123741] = 16'b0000000000000000;
	sram_mem[123742] = 16'b0000000000000000;
	sram_mem[123743] = 16'b0000000000000000;
	sram_mem[123744] = 16'b0000000000000000;
	sram_mem[123745] = 16'b0000000000000000;
	sram_mem[123746] = 16'b0000000000000000;
	sram_mem[123747] = 16'b0000000000000000;
	sram_mem[123748] = 16'b0000000000000000;
	sram_mem[123749] = 16'b0000000000000000;
	sram_mem[123750] = 16'b0000000000000000;
	sram_mem[123751] = 16'b0000000000000000;
	sram_mem[123752] = 16'b0000000000000000;
	sram_mem[123753] = 16'b0000000000000000;
	sram_mem[123754] = 16'b0000000000000000;
	sram_mem[123755] = 16'b0000000000000000;
	sram_mem[123756] = 16'b0000000000000000;
	sram_mem[123757] = 16'b0000000000000000;
	sram_mem[123758] = 16'b0000000000000000;
	sram_mem[123759] = 16'b0000000000000000;
	sram_mem[123760] = 16'b0000000000000000;
	sram_mem[123761] = 16'b0000000000000000;
	sram_mem[123762] = 16'b0000000000000000;
	sram_mem[123763] = 16'b0000000000000000;
	sram_mem[123764] = 16'b0000000000000000;
	sram_mem[123765] = 16'b0000000000000000;
	sram_mem[123766] = 16'b0000000000000000;
	sram_mem[123767] = 16'b0000000000000000;
	sram_mem[123768] = 16'b0000000000000000;
	sram_mem[123769] = 16'b0000000000000000;
	sram_mem[123770] = 16'b0000000000000000;
	sram_mem[123771] = 16'b0000000000000000;
	sram_mem[123772] = 16'b0000000000000000;
	sram_mem[123773] = 16'b0000000000000000;
	sram_mem[123774] = 16'b0000000000000000;
	sram_mem[123775] = 16'b0000000000000000;
	sram_mem[123776] = 16'b0000000000000000;
	sram_mem[123777] = 16'b0000000000000000;
	sram_mem[123778] = 16'b0000000000000000;
	sram_mem[123779] = 16'b0000000000000000;
	sram_mem[123780] = 16'b0000000000000000;
	sram_mem[123781] = 16'b0000000000000000;
	sram_mem[123782] = 16'b0000000000000000;
	sram_mem[123783] = 16'b0000000000000000;
	sram_mem[123784] = 16'b0000000000000000;
	sram_mem[123785] = 16'b0000000000000000;
	sram_mem[123786] = 16'b0000000000000000;
	sram_mem[123787] = 16'b0000000000000000;
	sram_mem[123788] = 16'b0000000000000000;
	sram_mem[123789] = 16'b0000000000000000;
	sram_mem[123790] = 16'b0000000000000000;
	sram_mem[123791] = 16'b0000000000000000;
	sram_mem[123792] = 16'b0000000000000000;
	sram_mem[123793] = 16'b0000000000000000;
	sram_mem[123794] = 16'b0000000000000000;
	sram_mem[123795] = 16'b0000000000000000;
	sram_mem[123796] = 16'b0000000000000000;
	sram_mem[123797] = 16'b0000000000000000;
	sram_mem[123798] = 16'b0000000000000000;
	sram_mem[123799] = 16'b0000000000000000;
	sram_mem[123800] = 16'b0000000000000000;
	sram_mem[123801] = 16'b0000000000000000;
	sram_mem[123802] = 16'b0000000000000000;
	sram_mem[123803] = 16'b0000000000000000;
	sram_mem[123804] = 16'b0000000000000000;
	sram_mem[123805] = 16'b0000000000000000;
	sram_mem[123806] = 16'b0000000000000000;
	sram_mem[123807] = 16'b0000000000000000;
	sram_mem[123808] = 16'b0000000000000000;
	sram_mem[123809] = 16'b0000000000000000;
	sram_mem[123810] = 16'b0000000000000000;
	sram_mem[123811] = 16'b0000000000000000;
	sram_mem[123812] = 16'b0000000000000000;
	sram_mem[123813] = 16'b0000000000000000;
	sram_mem[123814] = 16'b0000000000000000;
	sram_mem[123815] = 16'b0000000000000000;
	sram_mem[123816] = 16'b0000000000000000;
	sram_mem[123817] = 16'b0000000000000000;
	sram_mem[123818] = 16'b0000000000000000;
	sram_mem[123819] = 16'b0000000000000000;
	sram_mem[123820] = 16'b0000000000000000;
	sram_mem[123821] = 16'b0000000000000000;
	sram_mem[123822] = 16'b0000000000000000;
	sram_mem[123823] = 16'b0000000000000000;
	sram_mem[123824] = 16'b0000000000000000;
	sram_mem[123825] = 16'b0000000000000000;
	sram_mem[123826] = 16'b0000000000000000;
	sram_mem[123827] = 16'b0000000000000000;
	sram_mem[123828] = 16'b0000000000000000;
	sram_mem[123829] = 16'b0000000000000000;
	sram_mem[123830] = 16'b0000000000000000;
	sram_mem[123831] = 16'b0000000000000000;
	sram_mem[123832] = 16'b0000000000000000;
	sram_mem[123833] = 16'b0000000000000000;
	sram_mem[123834] = 16'b0000000000000000;
	sram_mem[123835] = 16'b0000000000000000;
	sram_mem[123836] = 16'b0000000000000000;
	sram_mem[123837] = 16'b0000000000000000;
	sram_mem[123838] = 16'b0000000000000000;
	sram_mem[123839] = 16'b0000000000000000;
	sram_mem[123840] = 16'b0000000000000000;
	sram_mem[123841] = 16'b0000000000000000;
	sram_mem[123842] = 16'b0000000000000000;
	sram_mem[123843] = 16'b0000000000000000;
	sram_mem[123844] = 16'b0000000000000000;
	sram_mem[123845] = 16'b0000000000000000;
	sram_mem[123846] = 16'b0000000000000000;
	sram_mem[123847] = 16'b0000000000000000;
	sram_mem[123848] = 16'b0000000000000000;
	sram_mem[123849] = 16'b0000000000000000;
	sram_mem[123850] = 16'b0000000000000000;
	sram_mem[123851] = 16'b0000000000000000;
	sram_mem[123852] = 16'b0000000000000000;
	sram_mem[123853] = 16'b0000000000000000;
	sram_mem[123854] = 16'b0000000000000000;
	sram_mem[123855] = 16'b0000000000000000;
	sram_mem[123856] = 16'b0000000000000000;
	sram_mem[123857] = 16'b0000000000000000;
	sram_mem[123858] = 16'b0000000000000000;
	sram_mem[123859] = 16'b0000000000000000;
	sram_mem[123860] = 16'b0000000000000000;
	sram_mem[123861] = 16'b0000000000000000;
	sram_mem[123862] = 16'b0000000000000000;
	sram_mem[123863] = 16'b0000000000000000;
	sram_mem[123864] = 16'b0000000000000000;
	sram_mem[123865] = 16'b0000000000000000;
	sram_mem[123866] = 16'b0000000000000000;
	sram_mem[123867] = 16'b0000000000000000;
	sram_mem[123868] = 16'b0000000000000000;
	sram_mem[123869] = 16'b0000000000000000;
	sram_mem[123870] = 16'b0000000000000000;
	sram_mem[123871] = 16'b0000000000000000;
	sram_mem[123872] = 16'b0000000000000000;
	sram_mem[123873] = 16'b0000000000000000;
	sram_mem[123874] = 16'b0000000000000000;
	sram_mem[123875] = 16'b0000000000000000;
	sram_mem[123876] = 16'b0000000000000000;
	sram_mem[123877] = 16'b0000000000000000;
	sram_mem[123878] = 16'b0000000000000000;
	sram_mem[123879] = 16'b0000000000000000;
	sram_mem[123880] = 16'b0000000000000000;
	sram_mem[123881] = 16'b0000000000000000;
	sram_mem[123882] = 16'b0000000000000000;
	sram_mem[123883] = 16'b0000000000000000;
	sram_mem[123884] = 16'b0000000000000000;
	sram_mem[123885] = 16'b0000000000000000;
	sram_mem[123886] = 16'b0000000000000000;
	sram_mem[123887] = 16'b0000000000000000;
	sram_mem[123888] = 16'b0000000000000000;
	sram_mem[123889] = 16'b0000000000000000;
	sram_mem[123890] = 16'b0000000000000000;
	sram_mem[123891] = 16'b0000000000000000;
	sram_mem[123892] = 16'b0000000000000000;
	sram_mem[123893] = 16'b0000000000000000;
	sram_mem[123894] = 16'b0000000000000000;
	sram_mem[123895] = 16'b0000000000000000;
	sram_mem[123896] = 16'b0000000000000000;
	sram_mem[123897] = 16'b0000000000000000;
	sram_mem[123898] = 16'b0000000000000000;
	sram_mem[123899] = 16'b0000000000000000;
	sram_mem[123900] = 16'b0000000000000000;
	sram_mem[123901] = 16'b0000000000000000;
	sram_mem[123902] = 16'b0000000000000000;
	sram_mem[123903] = 16'b0000000000000000;
	sram_mem[123904] = 16'b0000000000000000;
	sram_mem[123905] = 16'b0000000000000000;
	sram_mem[123906] = 16'b0000000000000000;
	sram_mem[123907] = 16'b0000000000000000;
	sram_mem[123908] = 16'b0000000000000000;
	sram_mem[123909] = 16'b0000000000000000;
	sram_mem[123910] = 16'b0000000000000000;
	sram_mem[123911] = 16'b0000000000000000;
	sram_mem[123912] = 16'b0000000000000000;
	sram_mem[123913] = 16'b0000000000000000;
	sram_mem[123914] = 16'b0000000000000000;
	sram_mem[123915] = 16'b0000000000000000;
	sram_mem[123916] = 16'b0000000000000000;
	sram_mem[123917] = 16'b0000000000000000;
	sram_mem[123918] = 16'b0000000000000000;
	sram_mem[123919] = 16'b0000000000000000;
	sram_mem[123920] = 16'b0000000000000000;
	sram_mem[123921] = 16'b0000000000000000;
	sram_mem[123922] = 16'b0000000000000000;
	sram_mem[123923] = 16'b0000000000000000;
	sram_mem[123924] = 16'b0000000000000000;
	sram_mem[123925] = 16'b0000000000000000;
	sram_mem[123926] = 16'b0000000000000000;
	sram_mem[123927] = 16'b0000000000000000;
	sram_mem[123928] = 16'b0000000000000000;
	sram_mem[123929] = 16'b0000000000000000;
	sram_mem[123930] = 16'b0000000000000000;
	sram_mem[123931] = 16'b0000000000000000;
	sram_mem[123932] = 16'b0000000000000000;
	sram_mem[123933] = 16'b0000000000000000;
	sram_mem[123934] = 16'b0000000000000000;
	sram_mem[123935] = 16'b0000000000000000;
	sram_mem[123936] = 16'b0000000000000000;
	sram_mem[123937] = 16'b0000000000000000;
	sram_mem[123938] = 16'b0000000000000000;
	sram_mem[123939] = 16'b0000000000000000;
	sram_mem[123940] = 16'b0000000000000000;
	sram_mem[123941] = 16'b0000000000000000;
	sram_mem[123942] = 16'b0000000000000000;
	sram_mem[123943] = 16'b0000000000000000;
	sram_mem[123944] = 16'b0000000000000000;
	sram_mem[123945] = 16'b0000000000000000;
	sram_mem[123946] = 16'b0000000000000000;
	sram_mem[123947] = 16'b0000000000000000;
	sram_mem[123948] = 16'b0000000000000000;
	sram_mem[123949] = 16'b0000000000000000;
	sram_mem[123950] = 16'b0000000000000000;
	sram_mem[123951] = 16'b0000000000000000;
	sram_mem[123952] = 16'b0000000000000000;
	sram_mem[123953] = 16'b0000000000000000;
	sram_mem[123954] = 16'b0000000000000000;
	sram_mem[123955] = 16'b0000000000000000;
	sram_mem[123956] = 16'b0000000000000000;
	sram_mem[123957] = 16'b0000000000000000;
	sram_mem[123958] = 16'b0000000000000000;
	sram_mem[123959] = 16'b0000000000000000;
	sram_mem[123960] = 16'b0000000000000000;
	sram_mem[123961] = 16'b0000000000000000;
	sram_mem[123962] = 16'b0000000000000000;
	sram_mem[123963] = 16'b0000000000000000;
	sram_mem[123964] = 16'b0000000000000000;
	sram_mem[123965] = 16'b0000000000000000;
	sram_mem[123966] = 16'b0000000000000000;
	sram_mem[123967] = 16'b0000000000000000;
	sram_mem[123968] = 16'b0000000000000000;
	sram_mem[123969] = 16'b0000000000000000;
	sram_mem[123970] = 16'b0000000000000000;
	sram_mem[123971] = 16'b0000000000000000;
	sram_mem[123972] = 16'b0000000000000000;
	sram_mem[123973] = 16'b0000000000000000;
	sram_mem[123974] = 16'b0000000000000000;
	sram_mem[123975] = 16'b0000000000000000;
	sram_mem[123976] = 16'b0000000000000000;
	sram_mem[123977] = 16'b0000000000000000;
	sram_mem[123978] = 16'b0000000000000000;
	sram_mem[123979] = 16'b0000000000000000;
	sram_mem[123980] = 16'b0000000000000000;
	sram_mem[123981] = 16'b0000000000000000;
	sram_mem[123982] = 16'b0000000000000000;
	sram_mem[123983] = 16'b0000000000000000;
	sram_mem[123984] = 16'b0000000000000000;
	sram_mem[123985] = 16'b0000000000000000;
	sram_mem[123986] = 16'b0000000000000000;
	sram_mem[123987] = 16'b0000000000000000;
	sram_mem[123988] = 16'b0000000000000000;
	sram_mem[123989] = 16'b0000000000000000;
	sram_mem[123990] = 16'b0000000000000000;
	sram_mem[123991] = 16'b0000000000000000;
	sram_mem[123992] = 16'b0000000000000000;
	sram_mem[123993] = 16'b0000000000000000;
	sram_mem[123994] = 16'b0000000000000000;
	sram_mem[123995] = 16'b0000000000000000;
	sram_mem[123996] = 16'b0000000000000000;
	sram_mem[123997] = 16'b0000000000000000;
	sram_mem[123998] = 16'b0000000000000000;
	sram_mem[123999] = 16'b0000000000000000;
	sram_mem[124000] = 16'b0000000000000000;
	sram_mem[124001] = 16'b0000000000000000;
	sram_mem[124002] = 16'b0000000000000000;
	sram_mem[124003] = 16'b0000000000000000;
	sram_mem[124004] = 16'b0000000000000000;
	sram_mem[124005] = 16'b0000000000000000;
	sram_mem[124006] = 16'b0000000000000000;
	sram_mem[124007] = 16'b0000000000000000;
	sram_mem[124008] = 16'b0000000000000000;
	sram_mem[124009] = 16'b0000000000000000;
	sram_mem[124010] = 16'b0000000000000000;
	sram_mem[124011] = 16'b0000000000000000;
	sram_mem[124012] = 16'b0000000000000000;
	sram_mem[124013] = 16'b0000000000000000;
	sram_mem[124014] = 16'b0000000000000000;
	sram_mem[124015] = 16'b0000000000000000;
	sram_mem[124016] = 16'b0000000000000000;
	sram_mem[124017] = 16'b0000000000000000;
	sram_mem[124018] = 16'b0000000000000000;
	sram_mem[124019] = 16'b0000000000000000;
	sram_mem[124020] = 16'b0000000000000000;
	sram_mem[124021] = 16'b0000000000000000;
	sram_mem[124022] = 16'b0000000000000000;
	sram_mem[124023] = 16'b0000000000000000;
	sram_mem[124024] = 16'b0000000000000000;
	sram_mem[124025] = 16'b0000000000000000;
	sram_mem[124026] = 16'b0000000000000000;
	sram_mem[124027] = 16'b0000000000000000;
	sram_mem[124028] = 16'b0000000000000000;
	sram_mem[124029] = 16'b0000000000000000;
	sram_mem[124030] = 16'b0000000000000000;
	sram_mem[124031] = 16'b0000000000000000;
	sram_mem[124032] = 16'b0000000000000000;
	sram_mem[124033] = 16'b0000000000000000;
	sram_mem[124034] = 16'b0000000000000000;
	sram_mem[124035] = 16'b0000000000000000;
	sram_mem[124036] = 16'b0000000000000000;
	sram_mem[124037] = 16'b0000000000000000;
	sram_mem[124038] = 16'b0000000000000000;
	sram_mem[124039] = 16'b0000000000000000;
	sram_mem[124040] = 16'b0000000000000000;
	sram_mem[124041] = 16'b0000000000000000;
	sram_mem[124042] = 16'b0000000000000000;
	sram_mem[124043] = 16'b0000000000000000;
	sram_mem[124044] = 16'b0000000000000000;
	sram_mem[124045] = 16'b0000000000000000;
	sram_mem[124046] = 16'b0000000000000000;
	sram_mem[124047] = 16'b0000000000000000;
	sram_mem[124048] = 16'b0000000000000000;
	sram_mem[124049] = 16'b0000000000000000;
	sram_mem[124050] = 16'b0000000000000000;
	sram_mem[124051] = 16'b0000000000000000;
	sram_mem[124052] = 16'b0000000000000000;
	sram_mem[124053] = 16'b0000000000000000;
	sram_mem[124054] = 16'b0000000000000000;
	sram_mem[124055] = 16'b0000000000000000;
	sram_mem[124056] = 16'b0000000000000000;
	sram_mem[124057] = 16'b0000000000000000;
	sram_mem[124058] = 16'b0000000000000000;
	sram_mem[124059] = 16'b0000000000000000;
	sram_mem[124060] = 16'b0000000000000000;
	sram_mem[124061] = 16'b0000000000000000;
	sram_mem[124062] = 16'b0000000000000000;
	sram_mem[124063] = 16'b0000000000000000;
	sram_mem[124064] = 16'b0000000000000000;
	sram_mem[124065] = 16'b0000000000000000;
	sram_mem[124066] = 16'b0000000000000000;
	sram_mem[124067] = 16'b0000000000000000;
	sram_mem[124068] = 16'b0000000000000000;
	sram_mem[124069] = 16'b0000000000000000;
	sram_mem[124070] = 16'b0000000000000000;
	sram_mem[124071] = 16'b0000000000000000;
	sram_mem[124072] = 16'b0000000000000000;
	sram_mem[124073] = 16'b0000000000000000;
	sram_mem[124074] = 16'b0000000000000000;
	sram_mem[124075] = 16'b0000000000000000;
	sram_mem[124076] = 16'b0000000000000000;
	sram_mem[124077] = 16'b0000000000000000;
	sram_mem[124078] = 16'b0000000000000000;
	sram_mem[124079] = 16'b0000000000000000;
	sram_mem[124080] = 16'b0000000000000000;
	sram_mem[124081] = 16'b0000000000000000;
	sram_mem[124082] = 16'b0000000000000000;
	sram_mem[124083] = 16'b0000000000000000;
	sram_mem[124084] = 16'b0000000000000000;
	sram_mem[124085] = 16'b0000000000000000;
	sram_mem[124086] = 16'b0000000000000000;
	sram_mem[124087] = 16'b0000000000000000;
	sram_mem[124088] = 16'b0000000000000000;
	sram_mem[124089] = 16'b0000000000000000;
	sram_mem[124090] = 16'b0000000000000000;
	sram_mem[124091] = 16'b0000000000000000;
	sram_mem[124092] = 16'b0000000000000000;
	sram_mem[124093] = 16'b0000000000000000;
	sram_mem[124094] = 16'b0000000000000000;
	sram_mem[124095] = 16'b0000000000000000;
	sram_mem[124096] = 16'b0000000000000000;
	sram_mem[124097] = 16'b0000000000000000;
	sram_mem[124098] = 16'b0000000000000000;
	sram_mem[124099] = 16'b0000000000000000;
	sram_mem[124100] = 16'b0000000000000000;
	sram_mem[124101] = 16'b0000000000000000;
	sram_mem[124102] = 16'b0000000000000000;
	sram_mem[124103] = 16'b0000000000000000;
	sram_mem[124104] = 16'b0000000000000000;
	sram_mem[124105] = 16'b0000000000000000;
	sram_mem[124106] = 16'b0000000000000000;
	sram_mem[124107] = 16'b0000000000000000;
	sram_mem[124108] = 16'b0000000000000000;
	sram_mem[124109] = 16'b0000000000000000;
	sram_mem[124110] = 16'b0000000000000000;
	sram_mem[124111] = 16'b0000000000000000;
	sram_mem[124112] = 16'b0000000000000000;
	sram_mem[124113] = 16'b0000000000000000;
	sram_mem[124114] = 16'b0000000000000000;
	sram_mem[124115] = 16'b0000000000000000;
	sram_mem[124116] = 16'b0000000000000000;
	sram_mem[124117] = 16'b0000000000000000;
	sram_mem[124118] = 16'b0000000000000000;
	sram_mem[124119] = 16'b0000000000000000;
	sram_mem[124120] = 16'b0000000000000000;
	sram_mem[124121] = 16'b0000000000000000;
	sram_mem[124122] = 16'b0000000000000000;
	sram_mem[124123] = 16'b0000000000000000;
	sram_mem[124124] = 16'b0000000000000000;
	sram_mem[124125] = 16'b0000000000000000;
	sram_mem[124126] = 16'b0000000000000000;
	sram_mem[124127] = 16'b0000000000000000;
	sram_mem[124128] = 16'b0000000000000000;
	sram_mem[124129] = 16'b0000000000000000;
	sram_mem[124130] = 16'b0000000000000000;
	sram_mem[124131] = 16'b0000000000000000;
	sram_mem[124132] = 16'b0000000000000000;
	sram_mem[124133] = 16'b0000000000000000;
	sram_mem[124134] = 16'b0000000000000000;
	sram_mem[124135] = 16'b0000000000000000;
	sram_mem[124136] = 16'b0000000000000000;
	sram_mem[124137] = 16'b0000000000000000;
	sram_mem[124138] = 16'b0000000000000000;
	sram_mem[124139] = 16'b0000000000000000;
	sram_mem[124140] = 16'b0000000000000000;
	sram_mem[124141] = 16'b0000000000000000;
	sram_mem[124142] = 16'b0000000000000000;
	sram_mem[124143] = 16'b0000000000000000;
	sram_mem[124144] = 16'b0000000000000000;
	sram_mem[124145] = 16'b0000000000000000;
	sram_mem[124146] = 16'b0000000000000000;
	sram_mem[124147] = 16'b0000000000000000;
	sram_mem[124148] = 16'b0000000000000000;
	sram_mem[124149] = 16'b0000000000000000;
	sram_mem[124150] = 16'b0000000000000000;
	sram_mem[124151] = 16'b0000000000000000;
	sram_mem[124152] = 16'b0000000000000000;
	sram_mem[124153] = 16'b0000000000000000;
	sram_mem[124154] = 16'b0000000000000000;
	sram_mem[124155] = 16'b0000000000000000;
	sram_mem[124156] = 16'b0000000000000000;
	sram_mem[124157] = 16'b0000000000000000;
	sram_mem[124158] = 16'b0000000000000000;
	sram_mem[124159] = 16'b0000000000000000;
	sram_mem[124160] = 16'b0000000000000000;
	sram_mem[124161] = 16'b0000000000000000;
	sram_mem[124162] = 16'b0000000000000000;
	sram_mem[124163] = 16'b0000000000000000;
	sram_mem[124164] = 16'b0000000000000000;
	sram_mem[124165] = 16'b0000000000000000;
	sram_mem[124166] = 16'b0000000000000000;
	sram_mem[124167] = 16'b0000000000000000;
	sram_mem[124168] = 16'b0000000000000000;
	sram_mem[124169] = 16'b0000000000000000;
	sram_mem[124170] = 16'b0000000000000000;
	sram_mem[124171] = 16'b0000000000000000;
	sram_mem[124172] = 16'b0000000000000000;
	sram_mem[124173] = 16'b0000000000000000;
	sram_mem[124174] = 16'b0000000000000000;
	sram_mem[124175] = 16'b0000000000000000;
	sram_mem[124176] = 16'b0000000000000000;
	sram_mem[124177] = 16'b0000000000000000;
	sram_mem[124178] = 16'b0000000000000000;
	sram_mem[124179] = 16'b0000000000000000;
	sram_mem[124180] = 16'b0000000000000000;
	sram_mem[124181] = 16'b0000000000000000;
	sram_mem[124182] = 16'b0000000000000000;
	sram_mem[124183] = 16'b0000000000000000;
	sram_mem[124184] = 16'b0000000000000000;
	sram_mem[124185] = 16'b0000000000000000;
	sram_mem[124186] = 16'b0000000000000000;
	sram_mem[124187] = 16'b0000000000000000;
	sram_mem[124188] = 16'b0000000000000000;
	sram_mem[124189] = 16'b0000000000000000;
	sram_mem[124190] = 16'b0000000000000000;
	sram_mem[124191] = 16'b0000000000000000;
	sram_mem[124192] = 16'b0000000000000000;
	sram_mem[124193] = 16'b0000000000000000;
	sram_mem[124194] = 16'b0000000000000000;
	sram_mem[124195] = 16'b0000000000000000;
	sram_mem[124196] = 16'b0000000000000000;
	sram_mem[124197] = 16'b0000000000000000;
	sram_mem[124198] = 16'b0000000000000000;
	sram_mem[124199] = 16'b0000000000000000;
	sram_mem[124200] = 16'b0000000000000000;
	sram_mem[124201] = 16'b0000000000000000;
	sram_mem[124202] = 16'b0000000000000000;
	sram_mem[124203] = 16'b0000000000000000;
	sram_mem[124204] = 16'b0000000000000000;
	sram_mem[124205] = 16'b0000000000000000;
	sram_mem[124206] = 16'b0000000000000000;
	sram_mem[124207] = 16'b0000000000000000;
	sram_mem[124208] = 16'b0000000000000000;
	sram_mem[124209] = 16'b0000000000000000;
	sram_mem[124210] = 16'b0000000000000000;
	sram_mem[124211] = 16'b0000000000000000;
	sram_mem[124212] = 16'b0000000000000000;
	sram_mem[124213] = 16'b0000000000000000;
	sram_mem[124214] = 16'b0000000000000000;
	sram_mem[124215] = 16'b0000000000000000;
	sram_mem[124216] = 16'b0000000000000000;
	sram_mem[124217] = 16'b0000000000000000;
	sram_mem[124218] = 16'b0000000000000000;
	sram_mem[124219] = 16'b0000000000000000;
	sram_mem[124220] = 16'b0000000000000000;
	sram_mem[124221] = 16'b0000000000000000;
	sram_mem[124222] = 16'b0000000000000000;
	sram_mem[124223] = 16'b0000000000000000;
	sram_mem[124224] = 16'b0000000000000000;
	sram_mem[124225] = 16'b0000000000000000;
	sram_mem[124226] = 16'b0000000000000000;
	sram_mem[124227] = 16'b0000000000000000;
	sram_mem[124228] = 16'b0000000000000000;
	sram_mem[124229] = 16'b0000000000000000;
	sram_mem[124230] = 16'b0000000000000000;
	sram_mem[124231] = 16'b0000000000000000;
	sram_mem[124232] = 16'b0000000000000000;
	sram_mem[124233] = 16'b0000000000000000;
	sram_mem[124234] = 16'b0000000000000000;
	sram_mem[124235] = 16'b0000000000000000;
	sram_mem[124236] = 16'b0000000000000000;
	sram_mem[124237] = 16'b0000000000000000;
	sram_mem[124238] = 16'b0000000000000000;
	sram_mem[124239] = 16'b0000000000000000;
	sram_mem[124240] = 16'b0000000000000000;
	sram_mem[124241] = 16'b0000000000000000;
	sram_mem[124242] = 16'b0000000000000000;
	sram_mem[124243] = 16'b0000000000000000;
	sram_mem[124244] = 16'b0000000000000000;
	sram_mem[124245] = 16'b0000000000000000;
	sram_mem[124246] = 16'b0000000000000000;
	sram_mem[124247] = 16'b0000000000000000;
	sram_mem[124248] = 16'b0000000000000000;
	sram_mem[124249] = 16'b0000000000000000;
	sram_mem[124250] = 16'b0000000000000000;
	sram_mem[124251] = 16'b0000000000000000;
	sram_mem[124252] = 16'b0000000000000000;
	sram_mem[124253] = 16'b0000000000000000;
	sram_mem[124254] = 16'b0000000000000000;
	sram_mem[124255] = 16'b0000000000000000;
	sram_mem[124256] = 16'b0000000000000000;
	sram_mem[124257] = 16'b0000000000000000;
	sram_mem[124258] = 16'b0000000000000000;
	sram_mem[124259] = 16'b0000000000000000;
	sram_mem[124260] = 16'b0000000000000000;
	sram_mem[124261] = 16'b0000000000000000;
	sram_mem[124262] = 16'b0000000000000000;
	sram_mem[124263] = 16'b0000000000000000;
	sram_mem[124264] = 16'b0000000000000000;
	sram_mem[124265] = 16'b0000000000000000;
	sram_mem[124266] = 16'b0000000000000000;
	sram_mem[124267] = 16'b0000000000000000;
	sram_mem[124268] = 16'b0000000000000000;
	sram_mem[124269] = 16'b0000000000000000;
	sram_mem[124270] = 16'b0000000000000000;
	sram_mem[124271] = 16'b0000000000000000;
	sram_mem[124272] = 16'b0000000000000000;
	sram_mem[124273] = 16'b0000000000000000;
	sram_mem[124274] = 16'b0000000000000000;
	sram_mem[124275] = 16'b0000000000000000;
	sram_mem[124276] = 16'b0000000000000000;
	sram_mem[124277] = 16'b0000000000000000;
	sram_mem[124278] = 16'b0000000000000000;
	sram_mem[124279] = 16'b0000000000000000;
	sram_mem[124280] = 16'b0000000000000000;
	sram_mem[124281] = 16'b0000000000000000;
	sram_mem[124282] = 16'b0000000000000000;
	sram_mem[124283] = 16'b0000000000000000;
	sram_mem[124284] = 16'b0000000000000000;
	sram_mem[124285] = 16'b0000000000000000;
	sram_mem[124286] = 16'b0000000000000000;
	sram_mem[124287] = 16'b0000000000000000;
	sram_mem[124288] = 16'b0000000000000000;
	sram_mem[124289] = 16'b0000000000000000;
	sram_mem[124290] = 16'b0000000000000000;
	sram_mem[124291] = 16'b0000000000000000;
	sram_mem[124292] = 16'b0000000000000000;
	sram_mem[124293] = 16'b0000000000000000;
	sram_mem[124294] = 16'b0000000000000000;
	sram_mem[124295] = 16'b0000000000000000;
	sram_mem[124296] = 16'b0000000000000000;
	sram_mem[124297] = 16'b0000000000000000;
	sram_mem[124298] = 16'b0000000000000000;
	sram_mem[124299] = 16'b0000000000000000;
	sram_mem[124300] = 16'b0000000000000000;
	sram_mem[124301] = 16'b0000000000000000;
	sram_mem[124302] = 16'b0000000000000000;
	sram_mem[124303] = 16'b0000000000000000;
	sram_mem[124304] = 16'b0000000000000000;
	sram_mem[124305] = 16'b0000000000000000;
	sram_mem[124306] = 16'b0000000000000000;
	sram_mem[124307] = 16'b0000000000000000;
	sram_mem[124308] = 16'b0000000000000000;
	sram_mem[124309] = 16'b0000000000000000;
	sram_mem[124310] = 16'b0000000000000000;
	sram_mem[124311] = 16'b0000000000000000;
	sram_mem[124312] = 16'b0000000000000000;
	sram_mem[124313] = 16'b0000000000000000;
	sram_mem[124314] = 16'b0000000000000000;
	sram_mem[124315] = 16'b0000000000000000;
	sram_mem[124316] = 16'b0000000000000000;
	sram_mem[124317] = 16'b0000000000000000;
	sram_mem[124318] = 16'b0000000000000000;
	sram_mem[124319] = 16'b0000000000000000;
	sram_mem[124320] = 16'b0000000000000000;
	sram_mem[124321] = 16'b0000000000000000;
	sram_mem[124322] = 16'b0000000000000000;
	sram_mem[124323] = 16'b0000000000000000;
	sram_mem[124324] = 16'b0000000000000000;
	sram_mem[124325] = 16'b0000000000000000;
	sram_mem[124326] = 16'b0000000000000000;
	sram_mem[124327] = 16'b0000000000000000;
	sram_mem[124328] = 16'b0000000000000000;
	sram_mem[124329] = 16'b0000000000000000;
	sram_mem[124330] = 16'b0000000000000000;
	sram_mem[124331] = 16'b0000000000000000;
	sram_mem[124332] = 16'b0000000000000000;
	sram_mem[124333] = 16'b0000000000000000;
	sram_mem[124334] = 16'b0000000000000000;
	sram_mem[124335] = 16'b0000000000000000;
	sram_mem[124336] = 16'b0000000000000000;
	sram_mem[124337] = 16'b0000000000000000;
	sram_mem[124338] = 16'b0000000000000000;
	sram_mem[124339] = 16'b0000000000000000;
	sram_mem[124340] = 16'b0000000000000000;
	sram_mem[124341] = 16'b0000000000000000;
	sram_mem[124342] = 16'b0000000000000000;
	sram_mem[124343] = 16'b0000000000000000;
	sram_mem[124344] = 16'b0000000000000000;
	sram_mem[124345] = 16'b0000000000000000;
	sram_mem[124346] = 16'b0000000000000000;
	sram_mem[124347] = 16'b0000000000000000;
	sram_mem[124348] = 16'b0000000000000000;
	sram_mem[124349] = 16'b0000000000000000;
	sram_mem[124350] = 16'b0000000000000000;
	sram_mem[124351] = 16'b0000000000000000;
	sram_mem[124352] = 16'b0000000000000000;
	sram_mem[124353] = 16'b0000000000000000;
	sram_mem[124354] = 16'b0000000000000000;
	sram_mem[124355] = 16'b0000000000000000;
	sram_mem[124356] = 16'b0000000000000000;
	sram_mem[124357] = 16'b0000000000000000;
	sram_mem[124358] = 16'b0000000000000000;
	sram_mem[124359] = 16'b0000000000000000;
	sram_mem[124360] = 16'b0000000000000000;
	sram_mem[124361] = 16'b0000000000000000;
	sram_mem[124362] = 16'b0000000000000000;
	sram_mem[124363] = 16'b0000000000000000;
	sram_mem[124364] = 16'b0000000000000000;
	sram_mem[124365] = 16'b0000000000000000;
	sram_mem[124366] = 16'b0000000000000000;
	sram_mem[124367] = 16'b0000000000000000;
	sram_mem[124368] = 16'b0000000000000000;
	sram_mem[124369] = 16'b0000000000000000;
	sram_mem[124370] = 16'b0000000000000000;
	sram_mem[124371] = 16'b0000000000000000;
	sram_mem[124372] = 16'b0000000000000000;
	sram_mem[124373] = 16'b0000000000000000;
	sram_mem[124374] = 16'b0000000000000000;
	sram_mem[124375] = 16'b0000000000000000;
	sram_mem[124376] = 16'b0000000000000000;
	sram_mem[124377] = 16'b0000000000000000;
	sram_mem[124378] = 16'b0000000000000000;
	sram_mem[124379] = 16'b0000000000000000;
	sram_mem[124380] = 16'b0000000000000000;
	sram_mem[124381] = 16'b0000000000000000;
	sram_mem[124382] = 16'b0000000000000000;
	sram_mem[124383] = 16'b0000000000000000;
	sram_mem[124384] = 16'b0000000000000000;
	sram_mem[124385] = 16'b0000000000000000;
	sram_mem[124386] = 16'b0000000000000000;
	sram_mem[124387] = 16'b0000000000000000;
	sram_mem[124388] = 16'b0000000000000000;
	sram_mem[124389] = 16'b0000000000000000;
	sram_mem[124390] = 16'b0000000000000000;
	sram_mem[124391] = 16'b0000000000000000;
	sram_mem[124392] = 16'b0000000000000000;
	sram_mem[124393] = 16'b0000000000000000;
	sram_mem[124394] = 16'b0000000000000000;
	sram_mem[124395] = 16'b0000000000000000;
	sram_mem[124396] = 16'b0000000000000000;
	sram_mem[124397] = 16'b0000000000000000;
	sram_mem[124398] = 16'b0000000000000000;
	sram_mem[124399] = 16'b0000000000000000;
	sram_mem[124400] = 16'b0000000000000000;
	sram_mem[124401] = 16'b0000000000000000;
	sram_mem[124402] = 16'b0000000000000000;
	sram_mem[124403] = 16'b0000000000000000;
	sram_mem[124404] = 16'b0000000000000000;
	sram_mem[124405] = 16'b0000000000000000;
	sram_mem[124406] = 16'b0000000000000000;
	sram_mem[124407] = 16'b0000000000000000;
	sram_mem[124408] = 16'b0000000000000000;
	sram_mem[124409] = 16'b0000000000000000;
	sram_mem[124410] = 16'b0000000000000000;
	sram_mem[124411] = 16'b0000000000000000;
	sram_mem[124412] = 16'b0000000000000000;
	sram_mem[124413] = 16'b0000000000000000;
	sram_mem[124414] = 16'b0000000000000000;
	sram_mem[124415] = 16'b0000000000000000;
	sram_mem[124416] = 16'b0000000000000000;
	sram_mem[124417] = 16'b0000000000000000;
	sram_mem[124418] = 16'b0000000000000000;
	sram_mem[124419] = 16'b0000000000000000;
	sram_mem[124420] = 16'b0000000000000000;
	sram_mem[124421] = 16'b0000000000000000;
	sram_mem[124422] = 16'b0000000000000000;
	sram_mem[124423] = 16'b0000000000000000;
	sram_mem[124424] = 16'b0000000000000000;
	sram_mem[124425] = 16'b0000000000000000;
	sram_mem[124426] = 16'b0000000000000000;
	sram_mem[124427] = 16'b0000000000000000;
	sram_mem[124428] = 16'b0000000000000000;
	sram_mem[124429] = 16'b0000000000000000;
	sram_mem[124430] = 16'b0000000000000000;
	sram_mem[124431] = 16'b0000000000000000;
	sram_mem[124432] = 16'b0000000000000000;
	sram_mem[124433] = 16'b0000000000000000;
	sram_mem[124434] = 16'b0000000000000000;
	sram_mem[124435] = 16'b0000000000000000;
	sram_mem[124436] = 16'b0000000000000000;
	sram_mem[124437] = 16'b0000000000000000;
	sram_mem[124438] = 16'b0000000000000000;
	sram_mem[124439] = 16'b0000000000000000;
	sram_mem[124440] = 16'b0000000000000000;
	sram_mem[124441] = 16'b0000000000000000;
	sram_mem[124442] = 16'b0000000000000000;
	sram_mem[124443] = 16'b0000000000000000;
	sram_mem[124444] = 16'b0000000000000000;
	sram_mem[124445] = 16'b0000000000000000;
	sram_mem[124446] = 16'b0000000000000000;
	sram_mem[124447] = 16'b0000000000000000;
	sram_mem[124448] = 16'b0000000000000000;
	sram_mem[124449] = 16'b0000000000000000;
	sram_mem[124450] = 16'b0000000000000000;
	sram_mem[124451] = 16'b0000000000000000;
	sram_mem[124452] = 16'b0000000000000000;
	sram_mem[124453] = 16'b0000000000000000;
	sram_mem[124454] = 16'b0000000000000000;
	sram_mem[124455] = 16'b0000000000000000;
	sram_mem[124456] = 16'b0000000000000000;
	sram_mem[124457] = 16'b0000000000000000;
	sram_mem[124458] = 16'b0000000000000000;
	sram_mem[124459] = 16'b0000000000000000;
	sram_mem[124460] = 16'b0000000000000000;
	sram_mem[124461] = 16'b0000000000000000;
	sram_mem[124462] = 16'b0000000000000000;
	sram_mem[124463] = 16'b0000000000000000;
	sram_mem[124464] = 16'b0000000000000000;
	sram_mem[124465] = 16'b0000000000000000;
	sram_mem[124466] = 16'b0000000000000000;
	sram_mem[124467] = 16'b0000000000000000;
	sram_mem[124468] = 16'b0000000000000000;
	sram_mem[124469] = 16'b0000000000000000;
	sram_mem[124470] = 16'b0000000000000000;
	sram_mem[124471] = 16'b0000000000000000;
	sram_mem[124472] = 16'b0000000000000000;
	sram_mem[124473] = 16'b0000000000000000;
	sram_mem[124474] = 16'b0000000000000000;
	sram_mem[124475] = 16'b0000000000000000;
	sram_mem[124476] = 16'b0000000000000000;
	sram_mem[124477] = 16'b0000000000000000;
	sram_mem[124478] = 16'b0000000000000000;
	sram_mem[124479] = 16'b0000000000000000;
	sram_mem[124480] = 16'b0000000000000000;
	sram_mem[124481] = 16'b0000000000000000;
	sram_mem[124482] = 16'b0000000000000000;
	sram_mem[124483] = 16'b0000000000000000;
	sram_mem[124484] = 16'b0000000000000000;
	sram_mem[124485] = 16'b0000000000000000;
	sram_mem[124486] = 16'b0000000000000000;
	sram_mem[124487] = 16'b0000000000000000;
	sram_mem[124488] = 16'b0000000000000000;
	sram_mem[124489] = 16'b0000000000000000;
	sram_mem[124490] = 16'b0000000000000000;
	sram_mem[124491] = 16'b0000000000000000;
	sram_mem[124492] = 16'b0000000000000000;
	sram_mem[124493] = 16'b0000000000000000;
	sram_mem[124494] = 16'b0000000000000000;
	sram_mem[124495] = 16'b0000000000000000;
	sram_mem[124496] = 16'b0000000000000000;
	sram_mem[124497] = 16'b0000000000000000;
	sram_mem[124498] = 16'b0000000000000000;
	sram_mem[124499] = 16'b0000000000000000;
	sram_mem[124500] = 16'b0000000000000000;
	sram_mem[124501] = 16'b0000000000000000;
	sram_mem[124502] = 16'b0000000000000000;
	sram_mem[124503] = 16'b0000000000000000;
	sram_mem[124504] = 16'b0000000000000000;
	sram_mem[124505] = 16'b0000000000000000;
	sram_mem[124506] = 16'b0000000000000000;
	sram_mem[124507] = 16'b0000000000000000;
	sram_mem[124508] = 16'b0000000000000000;
	sram_mem[124509] = 16'b0000000000000000;
	sram_mem[124510] = 16'b0000000000000000;
	sram_mem[124511] = 16'b0000000000000000;
	sram_mem[124512] = 16'b0000000000000000;
	sram_mem[124513] = 16'b0000000000000000;
	sram_mem[124514] = 16'b0000000000000000;
	sram_mem[124515] = 16'b0000000000000000;
	sram_mem[124516] = 16'b0000000000000000;
	sram_mem[124517] = 16'b0000000000000000;
	sram_mem[124518] = 16'b0000000000000000;
	sram_mem[124519] = 16'b0000000000000000;
	sram_mem[124520] = 16'b0000000000000000;
	sram_mem[124521] = 16'b0000000000000000;
	sram_mem[124522] = 16'b0000000000000000;
	sram_mem[124523] = 16'b0000000000000000;
	sram_mem[124524] = 16'b0000000000000000;
	sram_mem[124525] = 16'b0000000000000000;
	sram_mem[124526] = 16'b0000000000000000;
	sram_mem[124527] = 16'b0000000000000000;
	sram_mem[124528] = 16'b0000000000000000;
	sram_mem[124529] = 16'b0000000000000000;
	sram_mem[124530] = 16'b0000000000000000;
	sram_mem[124531] = 16'b0000000000000000;
	sram_mem[124532] = 16'b0000000000000000;
	sram_mem[124533] = 16'b0000000000000000;
	sram_mem[124534] = 16'b0000000000000000;
	sram_mem[124535] = 16'b0000000000000000;
	sram_mem[124536] = 16'b0000000000000000;
	sram_mem[124537] = 16'b0000000000000000;
	sram_mem[124538] = 16'b0000000000000000;
	sram_mem[124539] = 16'b0000000000000000;
	sram_mem[124540] = 16'b0000000000000000;
	sram_mem[124541] = 16'b0000000000000000;
	sram_mem[124542] = 16'b0000000000000000;
	sram_mem[124543] = 16'b0000000000000000;
	sram_mem[124544] = 16'b0000000000000000;
	sram_mem[124545] = 16'b0000000000000000;
	sram_mem[124546] = 16'b0000000000000000;
	sram_mem[124547] = 16'b0000000000000000;
	sram_mem[124548] = 16'b0000000000000000;
	sram_mem[124549] = 16'b0000000000000000;
	sram_mem[124550] = 16'b0000000000000000;
	sram_mem[124551] = 16'b0000000000000000;
	sram_mem[124552] = 16'b0000000000000000;
	sram_mem[124553] = 16'b0000000000000000;
	sram_mem[124554] = 16'b0000000000000000;
	sram_mem[124555] = 16'b0000000000000000;
	sram_mem[124556] = 16'b0000000000000000;
	sram_mem[124557] = 16'b0000000000000000;
	sram_mem[124558] = 16'b0000000000000000;
	sram_mem[124559] = 16'b0000000000000000;
	sram_mem[124560] = 16'b0000000000000000;
	sram_mem[124561] = 16'b0000000000000000;
	sram_mem[124562] = 16'b0000000000000000;
	sram_mem[124563] = 16'b0000000000000000;
	sram_mem[124564] = 16'b0000000000000000;
	sram_mem[124565] = 16'b0000000000000000;
	sram_mem[124566] = 16'b0000000000000000;
	sram_mem[124567] = 16'b0000000000000000;
	sram_mem[124568] = 16'b0000000000000000;
	sram_mem[124569] = 16'b0000000000000000;
	sram_mem[124570] = 16'b0000000000000000;
	sram_mem[124571] = 16'b0000000000000000;
	sram_mem[124572] = 16'b0000000000000000;
	sram_mem[124573] = 16'b0000000000000000;
	sram_mem[124574] = 16'b0000000000000000;
	sram_mem[124575] = 16'b0000000000000000;
	sram_mem[124576] = 16'b0000000000000000;
	sram_mem[124577] = 16'b0000000000000000;
	sram_mem[124578] = 16'b0000000000000000;
	sram_mem[124579] = 16'b0000000000000000;
	sram_mem[124580] = 16'b0000000000000000;
	sram_mem[124581] = 16'b0000000000000000;
	sram_mem[124582] = 16'b0000000000000000;
	sram_mem[124583] = 16'b0000000000000000;
	sram_mem[124584] = 16'b0000000000000000;
	sram_mem[124585] = 16'b0000000000000000;
	sram_mem[124586] = 16'b0000000000000000;
	sram_mem[124587] = 16'b0000000000000000;
	sram_mem[124588] = 16'b0000000000000000;
	sram_mem[124589] = 16'b0000000000000000;
	sram_mem[124590] = 16'b0000000000000000;
	sram_mem[124591] = 16'b0000000000000000;
	sram_mem[124592] = 16'b0000000000000000;
	sram_mem[124593] = 16'b0000000000000000;
	sram_mem[124594] = 16'b0000000000000000;
	sram_mem[124595] = 16'b0000000000000000;
	sram_mem[124596] = 16'b0000000000000000;
	sram_mem[124597] = 16'b0000000000000000;
	sram_mem[124598] = 16'b0000000000000000;
	sram_mem[124599] = 16'b0000000000000000;
	sram_mem[124600] = 16'b0000000000000000;
	sram_mem[124601] = 16'b0000000000000000;
	sram_mem[124602] = 16'b0000000000000000;
	sram_mem[124603] = 16'b0000000000000000;
	sram_mem[124604] = 16'b0000000000000000;
	sram_mem[124605] = 16'b0000000000000000;
	sram_mem[124606] = 16'b0000000000000000;
	sram_mem[124607] = 16'b0000000000000000;
	sram_mem[124608] = 16'b0000000000000000;
	sram_mem[124609] = 16'b0000000000000000;
	sram_mem[124610] = 16'b0000000000000000;
	sram_mem[124611] = 16'b0000000000000000;
	sram_mem[124612] = 16'b0000000000000000;
	sram_mem[124613] = 16'b0000000000000000;
	sram_mem[124614] = 16'b0000000000000000;
	sram_mem[124615] = 16'b0000000000000000;
	sram_mem[124616] = 16'b0000000000000000;
	sram_mem[124617] = 16'b0000000000000000;
	sram_mem[124618] = 16'b0000000000000000;
	sram_mem[124619] = 16'b0000000000000000;
	sram_mem[124620] = 16'b0000000000000000;
	sram_mem[124621] = 16'b0000000000000000;
	sram_mem[124622] = 16'b0000000000000000;
	sram_mem[124623] = 16'b0000000000000000;
	sram_mem[124624] = 16'b0000000000000000;
	sram_mem[124625] = 16'b0000000000000000;
	sram_mem[124626] = 16'b0000000000000000;
	sram_mem[124627] = 16'b0000000000000000;
	sram_mem[124628] = 16'b0000000000000000;
	sram_mem[124629] = 16'b0000000000000000;
	sram_mem[124630] = 16'b0000000000000000;
	sram_mem[124631] = 16'b0000000000000000;
	sram_mem[124632] = 16'b0000000000000000;
	sram_mem[124633] = 16'b0000000000000000;
	sram_mem[124634] = 16'b0000000000000000;
	sram_mem[124635] = 16'b0000000000000000;
	sram_mem[124636] = 16'b0000000000000000;
	sram_mem[124637] = 16'b0000000000000000;
	sram_mem[124638] = 16'b0000000000000000;
	sram_mem[124639] = 16'b0000000000000000;
	sram_mem[124640] = 16'b0000000000000000;
	sram_mem[124641] = 16'b0000000000000000;
	sram_mem[124642] = 16'b0000000000000000;
	sram_mem[124643] = 16'b0000000000000000;
	sram_mem[124644] = 16'b0000000000000000;
	sram_mem[124645] = 16'b0000000000000000;
	sram_mem[124646] = 16'b0000000000000000;
	sram_mem[124647] = 16'b0000000000000000;
	sram_mem[124648] = 16'b0000000000000000;
	sram_mem[124649] = 16'b0000000000000000;
	sram_mem[124650] = 16'b0000000000000000;
	sram_mem[124651] = 16'b0000000000000000;
	sram_mem[124652] = 16'b0000000000000000;
	sram_mem[124653] = 16'b0000000000000000;
	sram_mem[124654] = 16'b0000000000000000;
	sram_mem[124655] = 16'b0000000000000000;
	sram_mem[124656] = 16'b0000000000000000;
	sram_mem[124657] = 16'b0000000000000000;
	sram_mem[124658] = 16'b0000000000000000;
	sram_mem[124659] = 16'b0000000000000000;
	sram_mem[124660] = 16'b0000000000000000;
	sram_mem[124661] = 16'b0000000000000000;
	sram_mem[124662] = 16'b0000000000000000;
	sram_mem[124663] = 16'b0000000000000000;
	sram_mem[124664] = 16'b0000000000000000;
	sram_mem[124665] = 16'b0000000000000000;
	sram_mem[124666] = 16'b0000000000000000;
	sram_mem[124667] = 16'b0000000000000000;
	sram_mem[124668] = 16'b0000000000000000;
	sram_mem[124669] = 16'b0000000000000000;
	sram_mem[124670] = 16'b0000000000000000;
	sram_mem[124671] = 16'b0000000000000000;
	sram_mem[124672] = 16'b0000000000000000;
	sram_mem[124673] = 16'b0000000000000000;
	sram_mem[124674] = 16'b0000000000000000;
	sram_mem[124675] = 16'b0000000000000000;
	sram_mem[124676] = 16'b0000000000000000;
	sram_mem[124677] = 16'b0000000000000000;
	sram_mem[124678] = 16'b0000000000000000;
	sram_mem[124679] = 16'b0000000000000000;
	sram_mem[124680] = 16'b0000000000000000;
	sram_mem[124681] = 16'b0000000000000000;
	sram_mem[124682] = 16'b0000000000000000;
	sram_mem[124683] = 16'b0000000000000000;
	sram_mem[124684] = 16'b0000000000000000;
	sram_mem[124685] = 16'b0000000000000000;
	sram_mem[124686] = 16'b0000000000000000;
	sram_mem[124687] = 16'b0000000000000000;
	sram_mem[124688] = 16'b0000000000000000;
	sram_mem[124689] = 16'b0000000000000000;
	sram_mem[124690] = 16'b0000000000000000;
	sram_mem[124691] = 16'b0000000000000000;
	sram_mem[124692] = 16'b0000000000000000;
	sram_mem[124693] = 16'b0000000000000000;
	sram_mem[124694] = 16'b0000000000000000;
	sram_mem[124695] = 16'b0000000000000000;
	sram_mem[124696] = 16'b0000000000000000;
	sram_mem[124697] = 16'b0000000000000000;
	sram_mem[124698] = 16'b0000000000000000;
	sram_mem[124699] = 16'b0000000000000000;
	sram_mem[124700] = 16'b0000000000000000;
	sram_mem[124701] = 16'b0000000000000000;
	sram_mem[124702] = 16'b0000000000000000;
	sram_mem[124703] = 16'b0000000000000000;
	sram_mem[124704] = 16'b0000000000000000;
	sram_mem[124705] = 16'b0000000000000000;
	sram_mem[124706] = 16'b0000000000000000;
	sram_mem[124707] = 16'b0000000000000000;
	sram_mem[124708] = 16'b0000000000000000;
	sram_mem[124709] = 16'b0000000000000000;
	sram_mem[124710] = 16'b0000000000000000;
	sram_mem[124711] = 16'b0000000000000000;
	sram_mem[124712] = 16'b0000000000000000;
	sram_mem[124713] = 16'b0000000000000000;
	sram_mem[124714] = 16'b0000000000000000;
	sram_mem[124715] = 16'b0000000000000000;
	sram_mem[124716] = 16'b0000000000000000;
	sram_mem[124717] = 16'b0000000000000000;
	sram_mem[124718] = 16'b0000000000000000;
	sram_mem[124719] = 16'b0000000000000000;
	sram_mem[124720] = 16'b0000000000000000;
	sram_mem[124721] = 16'b0000000000000000;
	sram_mem[124722] = 16'b0000000000000000;
	sram_mem[124723] = 16'b0000000000000000;
	sram_mem[124724] = 16'b0000000000000000;
	sram_mem[124725] = 16'b0000000000000000;
	sram_mem[124726] = 16'b0000000000000000;
	sram_mem[124727] = 16'b0000000000000000;
	sram_mem[124728] = 16'b0000000000000000;
	sram_mem[124729] = 16'b0000000000000000;
	sram_mem[124730] = 16'b0000000000000000;
	sram_mem[124731] = 16'b0000000000000000;
	sram_mem[124732] = 16'b0000000000000000;
	sram_mem[124733] = 16'b0000000000000000;
	sram_mem[124734] = 16'b0000000000000000;
	sram_mem[124735] = 16'b0000000000000000;
	sram_mem[124736] = 16'b0000000000000000;
	sram_mem[124737] = 16'b0000000000000000;
	sram_mem[124738] = 16'b0000000000000000;
	sram_mem[124739] = 16'b0000000000000000;
	sram_mem[124740] = 16'b0000000000000000;
	sram_mem[124741] = 16'b0000000000000000;
	sram_mem[124742] = 16'b0000000000000000;
	sram_mem[124743] = 16'b0000000000000000;
	sram_mem[124744] = 16'b0000000000000000;
	sram_mem[124745] = 16'b0000000000000000;
	sram_mem[124746] = 16'b0000000000000000;
	sram_mem[124747] = 16'b0000000000000000;
	sram_mem[124748] = 16'b0000000000000000;
	sram_mem[124749] = 16'b0000000000000000;
	sram_mem[124750] = 16'b0000000000000000;
	sram_mem[124751] = 16'b0000000000000000;
	sram_mem[124752] = 16'b0000000000000000;
	sram_mem[124753] = 16'b0000000000000000;
	sram_mem[124754] = 16'b0000000000000000;
	sram_mem[124755] = 16'b0000000000000000;
	sram_mem[124756] = 16'b0000000000000000;
	sram_mem[124757] = 16'b0000000000000000;
	sram_mem[124758] = 16'b0000000000000000;
	sram_mem[124759] = 16'b0000000000000000;
	sram_mem[124760] = 16'b0000000000000000;
	sram_mem[124761] = 16'b0000000000000000;
	sram_mem[124762] = 16'b0000000000000000;
	sram_mem[124763] = 16'b0000000000000000;
	sram_mem[124764] = 16'b0000000000000000;
	sram_mem[124765] = 16'b0000000000000000;
	sram_mem[124766] = 16'b0000000000000000;
	sram_mem[124767] = 16'b0000000000000000;
	sram_mem[124768] = 16'b0000000000000000;
	sram_mem[124769] = 16'b0000000000000000;
	sram_mem[124770] = 16'b0000000000000000;
	sram_mem[124771] = 16'b0000000000000000;
	sram_mem[124772] = 16'b0000000000000000;
	sram_mem[124773] = 16'b0000000000000000;
	sram_mem[124774] = 16'b0000000000000000;
	sram_mem[124775] = 16'b0000000000000000;
	sram_mem[124776] = 16'b0000000000000000;
	sram_mem[124777] = 16'b0000000000000000;
	sram_mem[124778] = 16'b0000000000000000;
	sram_mem[124779] = 16'b0000000000000000;
	sram_mem[124780] = 16'b0000000000000000;
	sram_mem[124781] = 16'b0000000000000000;
	sram_mem[124782] = 16'b0000000000000000;
	sram_mem[124783] = 16'b0000000000000000;
	sram_mem[124784] = 16'b0000000000000000;
	sram_mem[124785] = 16'b0000000000000000;
	sram_mem[124786] = 16'b0000000000000000;
	sram_mem[124787] = 16'b0000000000000000;
	sram_mem[124788] = 16'b0000000000000000;
	sram_mem[124789] = 16'b0000000000000000;
	sram_mem[124790] = 16'b0000000000000000;
	sram_mem[124791] = 16'b0000000000000000;
	sram_mem[124792] = 16'b0000000000000000;
	sram_mem[124793] = 16'b0000000000000000;
	sram_mem[124794] = 16'b0000000000000000;
	sram_mem[124795] = 16'b0000000000000000;
	sram_mem[124796] = 16'b0000000000000000;
	sram_mem[124797] = 16'b0000000000000000;
	sram_mem[124798] = 16'b0000000000000000;
	sram_mem[124799] = 16'b0000000000000000;
	sram_mem[124800] = 16'b0000000000000000;
	sram_mem[124801] = 16'b0000000000000000;
	sram_mem[124802] = 16'b0000000000000000;
	sram_mem[124803] = 16'b0000000000000000;
	sram_mem[124804] = 16'b0000000000000000;
	sram_mem[124805] = 16'b0000000000000000;
	sram_mem[124806] = 16'b0000000000000000;
	sram_mem[124807] = 16'b0000000000000000;
	sram_mem[124808] = 16'b0000000000000000;
	sram_mem[124809] = 16'b0000000000000000;
	sram_mem[124810] = 16'b0000000000000000;
	sram_mem[124811] = 16'b0000000000000000;
	sram_mem[124812] = 16'b0000000000000000;
	sram_mem[124813] = 16'b0000000000000000;
	sram_mem[124814] = 16'b0000000000000000;
	sram_mem[124815] = 16'b0000000000000000;
	sram_mem[124816] = 16'b0000000000000000;
	sram_mem[124817] = 16'b0000000000000000;
	sram_mem[124818] = 16'b0000000000000000;
	sram_mem[124819] = 16'b0000000000000000;
	sram_mem[124820] = 16'b0000000000000000;
	sram_mem[124821] = 16'b0000000000000000;
	sram_mem[124822] = 16'b0000000000000000;
	sram_mem[124823] = 16'b0000000000000000;
	sram_mem[124824] = 16'b0000000000000000;
	sram_mem[124825] = 16'b0000000000000000;
	sram_mem[124826] = 16'b0000000000000000;
	sram_mem[124827] = 16'b0000000000000000;
	sram_mem[124828] = 16'b0000000000000000;
	sram_mem[124829] = 16'b0000000000000000;
	sram_mem[124830] = 16'b0000000000000000;
	sram_mem[124831] = 16'b0000000000000000;
	sram_mem[124832] = 16'b0000000000000000;
	sram_mem[124833] = 16'b0000000000000000;
	sram_mem[124834] = 16'b0000000000000000;
	sram_mem[124835] = 16'b0000000000000000;
	sram_mem[124836] = 16'b0000000000000000;
	sram_mem[124837] = 16'b0000000000000000;
	sram_mem[124838] = 16'b0000000000000000;
	sram_mem[124839] = 16'b0000000000000000;
	sram_mem[124840] = 16'b0000000000000000;
	sram_mem[124841] = 16'b0000000000000000;
	sram_mem[124842] = 16'b0000000000000000;
	sram_mem[124843] = 16'b0000000000000000;
	sram_mem[124844] = 16'b0000000000000000;
	sram_mem[124845] = 16'b0000000000000000;
	sram_mem[124846] = 16'b0000000000000000;
	sram_mem[124847] = 16'b0000000000000000;
	sram_mem[124848] = 16'b0000000000000000;
	sram_mem[124849] = 16'b0000000000000000;
	sram_mem[124850] = 16'b0000000000000000;
	sram_mem[124851] = 16'b0000000000000000;
	sram_mem[124852] = 16'b0000000000000000;
	sram_mem[124853] = 16'b0000000000000000;
	sram_mem[124854] = 16'b0000000000000000;
	sram_mem[124855] = 16'b0000000000000000;
	sram_mem[124856] = 16'b0000000000000000;
	sram_mem[124857] = 16'b0000000000000000;
	sram_mem[124858] = 16'b0000000000000000;
	sram_mem[124859] = 16'b0000000000000000;
	sram_mem[124860] = 16'b0000000000000000;
	sram_mem[124861] = 16'b0000000000000000;
	sram_mem[124862] = 16'b0000000000000000;
	sram_mem[124863] = 16'b0000000000000000;
	sram_mem[124864] = 16'b0000000000000000;
	sram_mem[124865] = 16'b0000000000000000;
	sram_mem[124866] = 16'b0000000000000000;
	sram_mem[124867] = 16'b0000000000000000;
	sram_mem[124868] = 16'b0000000000000000;
	sram_mem[124869] = 16'b0000000000000000;
	sram_mem[124870] = 16'b0000000000000000;
	sram_mem[124871] = 16'b0000000000000000;
	sram_mem[124872] = 16'b0000000000000000;
	sram_mem[124873] = 16'b0000000000000000;
	sram_mem[124874] = 16'b0000000000000000;
	sram_mem[124875] = 16'b0000000000000000;
	sram_mem[124876] = 16'b0000000000000000;
	sram_mem[124877] = 16'b0000000000000000;
	sram_mem[124878] = 16'b0000000000000000;
	sram_mem[124879] = 16'b0000000000000000;
	sram_mem[124880] = 16'b0000000000000000;
	sram_mem[124881] = 16'b0000000000000000;
	sram_mem[124882] = 16'b0000000000000000;
	sram_mem[124883] = 16'b0000000000000000;
	sram_mem[124884] = 16'b0000000000000000;
	sram_mem[124885] = 16'b0000000000000000;
	sram_mem[124886] = 16'b0000000000000000;
	sram_mem[124887] = 16'b0000000000000000;
	sram_mem[124888] = 16'b0000000000000000;
	sram_mem[124889] = 16'b0000000000000000;
	sram_mem[124890] = 16'b0000000000000000;
	sram_mem[124891] = 16'b0000000000000000;
	sram_mem[124892] = 16'b0000000000000000;
	sram_mem[124893] = 16'b0000000000000000;
	sram_mem[124894] = 16'b0000000000000000;
	sram_mem[124895] = 16'b0000000000000000;
	sram_mem[124896] = 16'b0000000000000000;
	sram_mem[124897] = 16'b0000000000000000;
	sram_mem[124898] = 16'b0000000000000000;
	sram_mem[124899] = 16'b0000000000000000;
	sram_mem[124900] = 16'b0000000000000000;
	sram_mem[124901] = 16'b0000000000000000;
	sram_mem[124902] = 16'b0000000000000000;
	sram_mem[124903] = 16'b0000000000000000;
	sram_mem[124904] = 16'b0000000000000000;
	sram_mem[124905] = 16'b0000000000000000;
	sram_mem[124906] = 16'b0000000000000000;
	sram_mem[124907] = 16'b0000000000000000;
	sram_mem[124908] = 16'b0000000000000000;
	sram_mem[124909] = 16'b0000000000000000;
	sram_mem[124910] = 16'b0000000000000000;
	sram_mem[124911] = 16'b0000000000000000;
	sram_mem[124912] = 16'b0000000000000000;
	sram_mem[124913] = 16'b0000000000000000;
	sram_mem[124914] = 16'b0000000000000000;
	sram_mem[124915] = 16'b0000000000000000;
	sram_mem[124916] = 16'b0000000000000000;
	sram_mem[124917] = 16'b0000000000000000;
	sram_mem[124918] = 16'b0000000000000000;
	sram_mem[124919] = 16'b0000000000000000;
	sram_mem[124920] = 16'b0000000000000000;
	sram_mem[124921] = 16'b0000000000000000;
	sram_mem[124922] = 16'b0000000000000000;
	sram_mem[124923] = 16'b0000000000000000;
	sram_mem[124924] = 16'b0000000000000000;
	sram_mem[124925] = 16'b0000000000000000;
	sram_mem[124926] = 16'b0000000000000000;
	sram_mem[124927] = 16'b0000000000000000;
	sram_mem[124928] = 16'b0000000000000000;
	sram_mem[124929] = 16'b0000000000000000;
	sram_mem[124930] = 16'b0000000000000000;
	sram_mem[124931] = 16'b0000000000000000;
	sram_mem[124932] = 16'b0000000000000000;
	sram_mem[124933] = 16'b0000000000000000;
	sram_mem[124934] = 16'b0000000000000000;
	sram_mem[124935] = 16'b0000000000000000;
	sram_mem[124936] = 16'b0000000000000000;
	sram_mem[124937] = 16'b0000000000000000;
	sram_mem[124938] = 16'b0000000000000000;
	sram_mem[124939] = 16'b0000000000000000;
	sram_mem[124940] = 16'b0000000000000000;
	sram_mem[124941] = 16'b0000000000000000;
	sram_mem[124942] = 16'b0000000000000000;
	sram_mem[124943] = 16'b0000000000000000;
	sram_mem[124944] = 16'b0000000000000000;
	sram_mem[124945] = 16'b0000000000000000;
	sram_mem[124946] = 16'b0000000000000000;
	sram_mem[124947] = 16'b0000000000000000;
	sram_mem[124948] = 16'b0000000000000000;
	sram_mem[124949] = 16'b0000000000000000;
	sram_mem[124950] = 16'b0000000000000000;
	sram_mem[124951] = 16'b0000000000000000;
	sram_mem[124952] = 16'b0000000000000000;
	sram_mem[124953] = 16'b0000000000000000;
	sram_mem[124954] = 16'b0000000000000000;
	sram_mem[124955] = 16'b0000000000000000;
	sram_mem[124956] = 16'b0000000000000000;
	sram_mem[124957] = 16'b0000000000000000;
	sram_mem[124958] = 16'b0000000000000000;
	sram_mem[124959] = 16'b0000000000000000;
	sram_mem[124960] = 16'b0000000000000000;
	sram_mem[124961] = 16'b0000000000000000;
	sram_mem[124962] = 16'b0000000000000000;
	sram_mem[124963] = 16'b0000000000000000;
	sram_mem[124964] = 16'b0000000000000000;
	sram_mem[124965] = 16'b0000000000000000;
	sram_mem[124966] = 16'b0000000000000000;
	sram_mem[124967] = 16'b0000000000000000;
	sram_mem[124968] = 16'b0000000000000000;
	sram_mem[124969] = 16'b0000000000000000;
	sram_mem[124970] = 16'b0000000000000000;
	sram_mem[124971] = 16'b0000000000000000;
	sram_mem[124972] = 16'b0000000000000000;
	sram_mem[124973] = 16'b0000000000000000;
	sram_mem[124974] = 16'b0000000000000000;
	sram_mem[124975] = 16'b0000000000000000;
	sram_mem[124976] = 16'b0000000000000000;
	sram_mem[124977] = 16'b0000000000000000;
	sram_mem[124978] = 16'b0000000000000000;
	sram_mem[124979] = 16'b0000000000000000;
	sram_mem[124980] = 16'b0000000000000000;
	sram_mem[124981] = 16'b0000000000000000;
	sram_mem[124982] = 16'b0000000000000000;
	sram_mem[124983] = 16'b0000000000000000;
	sram_mem[124984] = 16'b0000000000000000;
	sram_mem[124985] = 16'b0000000000000000;
	sram_mem[124986] = 16'b0000000000000000;
	sram_mem[124987] = 16'b0000000000000000;
	sram_mem[124988] = 16'b0000000000000000;
	sram_mem[124989] = 16'b0000000000000000;
	sram_mem[124990] = 16'b0000000000000000;
	sram_mem[124991] = 16'b0000000000000000;
	sram_mem[124992] = 16'b0000000000000000;
	sram_mem[124993] = 16'b0000000000000000;
	sram_mem[124994] = 16'b0000000000000000;
	sram_mem[124995] = 16'b0000000000000000;
	sram_mem[124996] = 16'b0000000000000000;
	sram_mem[124997] = 16'b0000000000000000;
	sram_mem[124998] = 16'b0000000000000000;
	sram_mem[124999] = 16'b0000000000000000;
	sram_mem[125000] = 16'b0000000000000000;
	sram_mem[125001] = 16'b0000000000000000;
	sram_mem[125002] = 16'b0000000000000000;
	sram_mem[125003] = 16'b0000000000000000;
	sram_mem[125004] = 16'b0000000000000000;
	sram_mem[125005] = 16'b0000000000000000;
	sram_mem[125006] = 16'b0000000000000000;
	sram_mem[125007] = 16'b0000000000000000;
	sram_mem[125008] = 16'b0000000000000000;
	sram_mem[125009] = 16'b0000000000000000;
	sram_mem[125010] = 16'b0000000000000000;
	sram_mem[125011] = 16'b0000000000000000;
	sram_mem[125012] = 16'b0000000000000000;
	sram_mem[125013] = 16'b0000000000000000;
	sram_mem[125014] = 16'b0000000000000000;
	sram_mem[125015] = 16'b0000000000000000;
	sram_mem[125016] = 16'b0000000000000000;
	sram_mem[125017] = 16'b0000000000000000;
	sram_mem[125018] = 16'b0000000000000000;
	sram_mem[125019] = 16'b0000000000000000;
	sram_mem[125020] = 16'b0000000000000000;
	sram_mem[125021] = 16'b0000000000000000;
	sram_mem[125022] = 16'b0000000000000000;
	sram_mem[125023] = 16'b0000000000000000;
	sram_mem[125024] = 16'b0000000000000000;
	sram_mem[125025] = 16'b0000000000000000;
	sram_mem[125026] = 16'b0000000000000000;
	sram_mem[125027] = 16'b0000000000000000;
	sram_mem[125028] = 16'b0000000000000000;
	sram_mem[125029] = 16'b0000000000000000;
	sram_mem[125030] = 16'b0000000000000000;
	sram_mem[125031] = 16'b0000000000000000;
	sram_mem[125032] = 16'b0000000000000000;
	sram_mem[125033] = 16'b0000000000000000;
	sram_mem[125034] = 16'b0000000000000000;
	sram_mem[125035] = 16'b0000000000000000;
	sram_mem[125036] = 16'b0000000000000000;
	sram_mem[125037] = 16'b0000000000000000;
	sram_mem[125038] = 16'b0000000000000000;
	sram_mem[125039] = 16'b0000000000000000;
	sram_mem[125040] = 16'b0000000000000000;
	sram_mem[125041] = 16'b0000000000000000;
	sram_mem[125042] = 16'b0000000000000000;
	sram_mem[125043] = 16'b0000000000000000;
	sram_mem[125044] = 16'b0000000000000000;
	sram_mem[125045] = 16'b0000000000000000;
	sram_mem[125046] = 16'b0000000000000000;
	sram_mem[125047] = 16'b0000000000000000;
	sram_mem[125048] = 16'b0000000000000000;
	sram_mem[125049] = 16'b0000000000000000;
	sram_mem[125050] = 16'b0000000000000000;
	sram_mem[125051] = 16'b0000000000000000;
	sram_mem[125052] = 16'b0000000000000000;
	sram_mem[125053] = 16'b0000000000000000;
	sram_mem[125054] = 16'b0000000000000000;
	sram_mem[125055] = 16'b0000000000000000;
	sram_mem[125056] = 16'b0000000000000000;
	sram_mem[125057] = 16'b0000000000000000;
	sram_mem[125058] = 16'b0000000000000000;
	sram_mem[125059] = 16'b0000000000000000;
	sram_mem[125060] = 16'b0000000000000000;
	sram_mem[125061] = 16'b0000000000000000;
	sram_mem[125062] = 16'b0000000000000000;
	sram_mem[125063] = 16'b0000000000000000;
	sram_mem[125064] = 16'b0000000000000000;
	sram_mem[125065] = 16'b0000000000000000;
	sram_mem[125066] = 16'b0000000000000000;
	sram_mem[125067] = 16'b0000000000000000;
	sram_mem[125068] = 16'b0000000000000000;
	sram_mem[125069] = 16'b0000000000000000;
	sram_mem[125070] = 16'b0000000000000000;
	sram_mem[125071] = 16'b0000000000000000;
	sram_mem[125072] = 16'b0000000000000000;
	sram_mem[125073] = 16'b0000000000000000;
	sram_mem[125074] = 16'b0000000000000000;
	sram_mem[125075] = 16'b0000000000000000;
	sram_mem[125076] = 16'b0000000000000000;
	sram_mem[125077] = 16'b0000000000000000;
	sram_mem[125078] = 16'b0000000000000000;
	sram_mem[125079] = 16'b0000000000000000;
	sram_mem[125080] = 16'b0000000000000000;
	sram_mem[125081] = 16'b0000000000000000;
	sram_mem[125082] = 16'b0000000000000000;
	sram_mem[125083] = 16'b0000000000000000;
	sram_mem[125084] = 16'b0000000000000000;
	sram_mem[125085] = 16'b0000000000000000;
	sram_mem[125086] = 16'b0000000000000000;
	sram_mem[125087] = 16'b0000000000000000;
	sram_mem[125088] = 16'b0000000000000000;
	sram_mem[125089] = 16'b0000000000000000;
	sram_mem[125090] = 16'b0000000000000000;
	sram_mem[125091] = 16'b0000000000000000;
	sram_mem[125092] = 16'b0000000000000000;
	sram_mem[125093] = 16'b0000000000000000;
	sram_mem[125094] = 16'b0000000000000000;
	sram_mem[125095] = 16'b0000000000000000;
	sram_mem[125096] = 16'b0000000000000000;
	sram_mem[125097] = 16'b0000000000000000;
	sram_mem[125098] = 16'b0000000000000000;
	sram_mem[125099] = 16'b0000000000000000;
	sram_mem[125100] = 16'b0000000000000000;
	sram_mem[125101] = 16'b0000000000000000;
	sram_mem[125102] = 16'b0000000000000000;
	sram_mem[125103] = 16'b0000000000000000;
	sram_mem[125104] = 16'b0000000000000000;
	sram_mem[125105] = 16'b0000000000000000;
	sram_mem[125106] = 16'b0000000000000000;
	sram_mem[125107] = 16'b0000000000000000;
	sram_mem[125108] = 16'b0000000000000000;
	sram_mem[125109] = 16'b0000000000000000;
	sram_mem[125110] = 16'b0000000000000000;
	sram_mem[125111] = 16'b0000000000000000;
	sram_mem[125112] = 16'b0000000000000000;
	sram_mem[125113] = 16'b0000000000000000;
	sram_mem[125114] = 16'b0000000000000000;
	sram_mem[125115] = 16'b0000000000000000;
	sram_mem[125116] = 16'b0000000000000000;
	sram_mem[125117] = 16'b0000000000000000;
	sram_mem[125118] = 16'b0000000000000000;
	sram_mem[125119] = 16'b0000000000000000;
	sram_mem[125120] = 16'b0000000000000000;
	sram_mem[125121] = 16'b0000000000000000;
	sram_mem[125122] = 16'b0000000000000000;
	sram_mem[125123] = 16'b0000000000000000;
	sram_mem[125124] = 16'b0000000000000000;
	sram_mem[125125] = 16'b0000000000000000;
	sram_mem[125126] = 16'b0000000000000000;
	sram_mem[125127] = 16'b0000000000000000;
	sram_mem[125128] = 16'b0000000000000000;
	sram_mem[125129] = 16'b0000000000000000;
	sram_mem[125130] = 16'b0000000000000000;
	sram_mem[125131] = 16'b0000000000000000;
	sram_mem[125132] = 16'b0000000000000000;
	sram_mem[125133] = 16'b0000000000000000;
	sram_mem[125134] = 16'b0000000000000000;
	sram_mem[125135] = 16'b0000000000000000;
	sram_mem[125136] = 16'b0000000000000000;
	sram_mem[125137] = 16'b0000000000000000;
	sram_mem[125138] = 16'b0000000000000000;
	sram_mem[125139] = 16'b0000000000000000;
	sram_mem[125140] = 16'b0000000000000000;
	sram_mem[125141] = 16'b0000000000000000;
	sram_mem[125142] = 16'b0000000000000000;
	sram_mem[125143] = 16'b0000000000000000;
	sram_mem[125144] = 16'b0000000000000000;
	sram_mem[125145] = 16'b0000000000000000;
	sram_mem[125146] = 16'b0000000000000000;
	sram_mem[125147] = 16'b0000000000000000;
	sram_mem[125148] = 16'b0000000000000000;
	sram_mem[125149] = 16'b0000000000000000;
	sram_mem[125150] = 16'b0000000000000000;
	sram_mem[125151] = 16'b0000000000000000;
	sram_mem[125152] = 16'b0000000000000000;
	sram_mem[125153] = 16'b0000000000000000;
	sram_mem[125154] = 16'b0000000000000000;
	sram_mem[125155] = 16'b0000000000000000;
	sram_mem[125156] = 16'b0000000000000000;
	sram_mem[125157] = 16'b0000000000000000;
	sram_mem[125158] = 16'b0000000000000000;
	sram_mem[125159] = 16'b0000000000000000;
	sram_mem[125160] = 16'b0000000000000000;
	sram_mem[125161] = 16'b0000000000000000;
	sram_mem[125162] = 16'b0000000000000000;
	sram_mem[125163] = 16'b0000000000000000;
	sram_mem[125164] = 16'b0000000000000000;
	sram_mem[125165] = 16'b0000000000000000;
	sram_mem[125166] = 16'b0000000000000000;
	sram_mem[125167] = 16'b0000000000000000;
	sram_mem[125168] = 16'b0000000000000000;
	sram_mem[125169] = 16'b0000000000000000;
	sram_mem[125170] = 16'b0000000000000000;
	sram_mem[125171] = 16'b0000000000000000;
	sram_mem[125172] = 16'b0000000000000000;
	sram_mem[125173] = 16'b0000000000000000;
	sram_mem[125174] = 16'b0000000000000000;
	sram_mem[125175] = 16'b0000000000000000;
	sram_mem[125176] = 16'b0000000000000000;
	sram_mem[125177] = 16'b0000000000000000;
	sram_mem[125178] = 16'b0000000000000000;
	sram_mem[125179] = 16'b0000000000000000;
	sram_mem[125180] = 16'b0000000000000000;
	sram_mem[125181] = 16'b0000000000000000;
	sram_mem[125182] = 16'b0000000000000000;
	sram_mem[125183] = 16'b0000000000000000;
	sram_mem[125184] = 16'b0000000000000000;
	sram_mem[125185] = 16'b0000000000000000;
	sram_mem[125186] = 16'b0000000000000000;
	sram_mem[125187] = 16'b0000000000000000;
	sram_mem[125188] = 16'b0000000000000000;
	sram_mem[125189] = 16'b0000000000000000;
	sram_mem[125190] = 16'b0000000000000000;
	sram_mem[125191] = 16'b0000000000000000;
	sram_mem[125192] = 16'b0000000000000000;
	sram_mem[125193] = 16'b0000000000000000;
	sram_mem[125194] = 16'b0000000000000000;
	sram_mem[125195] = 16'b0000000000000000;
	sram_mem[125196] = 16'b0000000000000000;
	sram_mem[125197] = 16'b0000000000000000;
	sram_mem[125198] = 16'b0000000000000000;
	sram_mem[125199] = 16'b0000000000000000;
	sram_mem[125200] = 16'b0000000000000000;
	sram_mem[125201] = 16'b0000000000000000;
	sram_mem[125202] = 16'b0000000000000000;
	sram_mem[125203] = 16'b0000000000000000;
	sram_mem[125204] = 16'b0000000000000000;
	sram_mem[125205] = 16'b0000000000000000;
	sram_mem[125206] = 16'b0000000000000000;
	sram_mem[125207] = 16'b0000000000000000;
	sram_mem[125208] = 16'b0000000000000000;
	sram_mem[125209] = 16'b0000000000000000;
	sram_mem[125210] = 16'b0000000000000000;
	sram_mem[125211] = 16'b0000000000000000;
	sram_mem[125212] = 16'b0000000000000000;
	sram_mem[125213] = 16'b0000000000000000;
	sram_mem[125214] = 16'b0000000000000000;
	sram_mem[125215] = 16'b0000000000000000;
	sram_mem[125216] = 16'b0000000000000000;
	sram_mem[125217] = 16'b0000000000000000;
	sram_mem[125218] = 16'b0000000000000000;
	sram_mem[125219] = 16'b0000000000000000;
	sram_mem[125220] = 16'b0000000000000000;
	sram_mem[125221] = 16'b0000000000000000;
	sram_mem[125222] = 16'b0000000000000000;
	sram_mem[125223] = 16'b0000000000000000;
	sram_mem[125224] = 16'b0000000000000000;
	sram_mem[125225] = 16'b0000000000000000;
	sram_mem[125226] = 16'b0000000000000000;
	sram_mem[125227] = 16'b0000000000000000;
	sram_mem[125228] = 16'b0000000000000000;
	sram_mem[125229] = 16'b0000000000000000;
	sram_mem[125230] = 16'b0000000000000000;
	sram_mem[125231] = 16'b0000000000000000;
	sram_mem[125232] = 16'b0000000000000000;
	sram_mem[125233] = 16'b0000000000000000;
	sram_mem[125234] = 16'b0000000000000000;
	sram_mem[125235] = 16'b0000000000000000;
	sram_mem[125236] = 16'b0000000000000000;
	sram_mem[125237] = 16'b0000000000000000;
	sram_mem[125238] = 16'b0000000000000000;
	sram_mem[125239] = 16'b0000000000000000;
	sram_mem[125240] = 16'b0000000000000000;
	sram_mem[125241] = 16'b0000000000000000;
	sram_mem[125242] = 16'b0000000000000000;
	sram_mem[125243] = 16'b0000000000000000;
	sram_mem[125244] = 16'b0000000000000000;
	sram_mem[125245] = 16'b0000000000000000;
	sram_mem[125246] = 16'b0000000000000000;
	sram_mem[125247] = 16'b0000000000000000;
	sram_mem[125248] = 16'b0000000000000000;
	sram_mem[125249] = 16'b0000000000000000;
	sram_mem[125250] = 16'b0000000000000000;
	sram_mem[125251] = 16'b0000000000000000;
	sram_mem[125252] = 16'b0000000000000000;
	sram_mem[125253] = 16'b0000000000000000;
	sram_mem[125254] = 16'b0000000000000000;
	sram_mem[125255] = 16'b0000000000000000;
	sram_mem[125256] = 16'b0000000000000000;
	sram_mem[125257] = 16'b0000000000000000;
	sram_mem[125258] = 16'b0000000000000000;
	sram_mem[125259] = 16'b0000000000000000;
	sram_mem[125260] = 16'b0000000000000000;
	sram_mem[125261] = 16'b0000000000000000;
	sram_mem[125262] = 16'b0000000000000000;
	sram_mem[125263] = 16'b0000000000000000;
	sram_mem[125264] = 16'b0000000000000000;
	sram_mem[125265] = 16'b0000000000000000;
	sram_mem[125266] = 16'b0000000000000000;
	sram_mem[125267] = 16'b0000000000000000;
	sram_mem[125268] = 16'b0000000000000000;
	sram_mem[125269] = 16'b0000000000000000;
	sram_mem[125270] = 16'b0000000000000000;
	sram_mem[125271] = 16'b0000000000000000;
	sram_mem[125272] = 16'b0000000000000000;
	sram_mem[125273] = 16'b0000000000000000;
	sram_mem[125274] = 16'b0000000000000000;
	sram_mem[125275] = 16'b0000000000000000;
	sram_mem[125276] = 16'b0000000000000000;
	sram_mem[125277] = 16'b0000000000000000;
	sram_mem[125278] = 16'b0000000000000000;
	sram_mem[125279] = 16'b0000000000000000;
	sram_mem[125280] = 16'b0000000000000000;
	sram_mem[125281] = 16'b0000000000000000;
	sram_mem[125282] = 16'b0000000000000000;
	sram_mem[125283] = 16'b0000000000000000;
	sram_mem[125284] = 16'b0000000000000000;
	sram_mem[125285] = 16'b0000000000000000;
	sram_mem[125286] = 16'b0000000000000000;
	sram_mem[125287] = 16'b0000000000000000;
	sram_mem[125288] = 16'b0000000000000000;
	sram_mem[125289] = 16'b0000000000000000;
	sram_mem[125290] = 16'b0000000000000000;
	sram_mem[125291] = 16'b0000000000000000;
	sram_mem[125292] = 16'b0000000000000000;
	sram_mem[125293] = 16'b0000000000000000;
	sram_mem[125294] = 16'b0000000000000000;
	sram_mem[125295] = 16'b0000000000000000;
	sram_mem[125296] = 16'b0000000000000000;
	sram_mem[125297] = 16'b0000000000000000;
	sram_mem[125298] = 16'b0000000000000000;
	sram_mem[125299] = 16'b0000000000000000;
	sram_mem[125300] = 16'b0000000000000000;
	sram_mem[125301] = 16'b0000000000000000;
	sram_mem[125302] = 16'b0000000000000000;
	sram_mem[125303] = 16'b0000000000000000;
	sram_mem[125304] = 16'b0000000000000000;
	sram_mem[125305] = 16'b0000000000000000;
	sram_mem[125306] = 16'b0000000000000000;
	sram_mem[125307] = 16'b0000000000000000;
	sram_mem[125308] = 16'b0000000000000000;
	sram_mem[125309] = 16'b0000000000000000;
	sram_mem[125310] = 16'b0000000000000000;
	sram_mem[125311] = 16'b0000000000000000;
	sram_mem[125312] = 16'b0000000000000000;
	sram_mem[125313] = 16'b0000000000000000;
	sram_mem[125314] = 16'b0000000000000000;
	sram_mem[125315] = 16'b0000000000000000;
	sram_mem[125316] = 16'b0000000000000000;
	sram_mem[125317] = 16'b0000000000000000;
	sram_mem[125318] = 16'b0000000000000000;
	sram_mem[125319] = 16'b0000000000000000;
	sram_mem[125320] = 16'b0000000000000000;
	sram_mem[125321] = 16'b0000000000000000;
	sram_mem[125322] = 16'b0000000000000000;
	sram_mem[125323] = 16'b0000000000000000;
	sram_mem[125324] = 16'b0000000000000000;
	sram_mem[125325] = 16'b0000000000000000;
	sram_mem[125326] = 16'b0000000000000000;
	sram_mem[125327] = 16'b0000000000000000;
	sram_mem[125328] = 16'b0000000000000000;
	sram_mem[125329] = 16'b0000000000000000;
	sram_mem[125330] = 16'b0000000000000000;
	sram_mem[125331] = 16'b0000000000000000;
	sram_mem[125332] = 16'b0000000000000000;
	sram_mem[125333] = 16'b0000000000000000;
	sram_mem[125334] = 16'b0000000000000000;
	sram_mem[125335] = 16'b0000000000000000;
	sram_mem[125336] = 16'b0000000000000000;
	sram_mem[125337] = 16'b0000000000000000;
	sram_mem[125338] = 16'b0000000000000000;
	sram_mem[125339] = 16'b0000000000000000;
	sram_mem[125340] = 16'b0000000000000000;
	sram_mem[125341] = 16'b0000000000000000;
	sram_mem[125342] = 16'b0000000000000000;
	sram_mem[125343] = 16'b0000000000000000;
	sram_mem[125344] = 16'b0000000000000000;
	sram_mem[125345] = 16'b0000000000000000;
	sram_mem[125346] = 16'b0000000000000000;
	sram_mem[125347] = 16'b0000000000000000;
	sram_mem[125348] = 16'b0000000000000000;
	sram_mem[125349] = 16'b0000000000000000;
	sram_mem[125350] = 16'b0000000000000000;
	sram_mem[125351] = 16'b0000000000000000;
	sram_mem[125352] = 16'b0000000000000000;
	sram_mem[125353] = 16'b0000000000000000;
	sram_mem[125354] = 16'b0000000000000000;
	sram_mem[125355] = 16'b0000000000000000;
	sram_mem[125356] = 16'b0000000000000000;
	sram_mem[125357] = 16'b0000000000000000;
	sram_mem[125358] = 16'b0000000000000000;
	sram_mem[125359] = 16'b0000000000000000;
	sram_mem[125360] = 16'b0000000000000000;
	sram_mem[125361] = 16'b0000000000000000;
	sram_mem[125362] = 16'b0000000000000000;
	sram_mem[125363] = 16'b0000000000000000;
	sram_mem[125364] = 16'b0000000000000000;
	sram_mem[125365] = 16'b0000000000000000;
	sram_mem[125366] = 16'b0000000000000000;
	sram_mem[125367] = 16'b0000000000000000;
	sram_mem[125368] = 16'b0000000000000000;
	sram_mem[125369] = 16'b0000000000000000;
	sram_mem[125370] = 16'b0000000000000000;
	sram_mem[125371] = 16'b0000000000000000;
	sram_mem[125372] = 16'b0000000000000000;
	sram_mem[125373] = 16'b0000000000000000;
	sram_mem[125374] = 16'b0000000000000000;
	sram_mem[125375] = 16'b0000000000000000;
	sram_mem[125376] = 16'b0000000000000000;
	sram_mem[125377] = 16'b0000000000000000;
	sram_mem[125378] = 16'b0000000000000000;
	sram_mem[125379] = 16'b0000000000000000;
	sram_mem[125380] = 16'b0000000000000000;
	sram_mem[125381] = 16'b0000000000000000;
	sram_mem[125382] = 16'b0000000000000000;
	sram_mem[125383] = 16'b0000000000000000;
	sram_mem[125384] = 16'b0000000000000000;
	sram_mem[125385] = 16'b0000000000000000;
	sram_mem[125386] = 16'b0000000000000000;
	sram_mem[125387] = 16'b0000000000000000;
	sram_mem[125388] = 16'b0000000000000000;
	sram_mem[125389] = 16'b0000000000000000;
	sram_mem[125390] = 16'b0000000000000000;
	sram_mem[125391] = 16'b0000000000000000;
	sram_mem[125392] = 16'b0000000000000000;
	sram_mem[125393] = 16'b0000000000000000;
	sram_mem[125394] = 16'b0000000000000000;
	sram_mem[125395] = 16'b0000000000000000;
	sram_mem[125396] = 16'b0000000000000000;
	sram_mem[125397] = 16'b0000000000000000;
	sram_mem[125398] = 16'b0000000000000000;
	sram_mem[125399] = 16'b0000000000000000;
	sram_mem[125400] = 16'b0000000000000000;
	sram_mem[125401] = 16'b0000000000000000;
	sram_mem[125402] = 16'b0000000000000000;
	sram_mem[125403] = 16'b0000000000000000;
	sram_mem[125404] = 16'b0000000000000000;
	sram_mem[125405] = 16'b0000000000000000;
	sram_mem[125406] = 16'b0000000000000000;
	sram_mem[125407] = 16'b0000000000000000;
	sram_mem[125408] = 16'b0000000000000000;
	sram_mem[125409] = 16'b0000000000000000;
	sram_mem[125410] = 16'b0000000000000000;
	sram_mem[125411] = 16'b0000000000000000;
	sram_mem[125412] = 16'b0000000000000000;
	sram_mem[125413] = 16'b0000000000000000;
	sram_mem[125414] = 16'b0000000000000000;
	sram_mem[125415] = 16'b0000000000000000;
	sram_mem[125416] = 16'b0000000000000000;
	sram_mem[125417] = 16'b0000000000000000;
	sram_mem[125418] = 16'b0000000000000000;
	sram_mem[125419] = 16'b0000000000000000;
	sram_mem[125420] = 16'b0000000000000000;
	sram_mem[125421] = 16'b0000000000000000;
	sram_mem[125422] = 16'b0000000000000000;
	sram_mem[125423] = 16'b0000000000000000;
	sram_mem[125424] = 16'b0000000000000000;
	sram_mem[125425] = 16'b0000000000000000;
	sram_mem[125426] = 16'b0000000000000000;
	sram_mem[125427] = 16'b0000000000000000;
	sram_mem[125428] = 16'b0000000000000000;
	sram_mem[125429] = 16'b0000000000000000;
	sram_mem[125430] = 16'b0000000000000000;
	sram_mem[125431] = 16'b0000000000000000;
	sram_mem[125432] = 16'b0000000000000000;
	sram_mem[125433] = 16'b0000000000000000;
	sram_mem[125434] = 16'b0000000000000000;
	sram_mem[125435] = 16'b0000000000000000;
	sram_mem[125436] = 16'b0000000000000000;
	sram_mem[125437] = 16'b0000000000000000;
	sram_mem[125438] = 16'b0000000000000000;
	sram_mem[125439] = 16'b0000000000000000;
	sram_mem[125440] = 16'b0000000000000000;
	sram_mem[125441] = 16'b0000000000000000;
	sram_mem[125442] = 16'b0000000000000000;
	sram_mem[125443] = 16'b0000000000000000;
	sram_mem[125444] = 16'b0000000000000000;
	sram_mem[125445] = 16'b0000000000000000;
	sram_mem[125446] = 16'b0000000000000000;
	sram_mem[125447] = 16'b0000000000000000;
	sram_mem[125448] = 16'b0000000000000000;
	sram_mem[125449] = 16'b0000000000000000;
	sram_mem[125450] = 16'b0000000000000000;
	sram_mem[125451] = 16'b0000000000000000;
	sram_mem[125452] = 16'b0000000000000000;
	sram_mem[125453] = 16'b0000000000000000;
	sram_mem[125454] = 16'b0000000000000000;
	sram_mem[125455] = 16'b0000000000000000;
	sram_mem[125456] = 16'b0000000000000000;
	sram_mem[125457] = 16'b0000000000000000;
	sram_mem[125458] = 16'b0000000000000000;
	sram_mem[125459] = 16'b0000000000000000;
	sram_mem[125460] = 16'b0000000000000000;
	sram_mem[125461] = 16'b0000000000000000;
	sram_mem[125462] = 16'b0000000000000000;
	sram_mem[125463] = 16'b0000000000000000;
	sram_mem[125464] = 16'b0000000000000000;
	sram_mem[125465] = 16'b0000000000000000;
	sram_mem[125466] = 16'b0000000000000000;
	sram_mem[125467] = 16'b0000000000000000;
	sram_mem[125468] = 16'b0000000000000000;
	sram_mem[125469] = 16'b0000000000000000;
	sram_mem[125470] = 16'b0000000000000000;
	sram_mem[125471] = 16'b0000000000000000;
	sram_mem[125472] = 16'b0000000000000000;
	sram_mem[125473] = 16'b0000000000000000;
	sram_mem[125474] = 16'b0000000000000000;
	sram_mem[125475] = 16'b0000000000000000;
	sram_mem[125476] = 16'b0000000000000000;
	sram_mem[125477] = 16'b0000000000000000;
	sram_mem[125478] = 16'b0000000000000000;
	sram_mem[125479] = 16'b0000000000000000;
	sram_mem[125480] = 16'b0000000000000000;
	sram_mem[125481] = 16'b0000000000000000;
	sram_mem[125482] = 16'b0000000000000000;
	sram_mem[125483] = 16'b0000000000000000;
	sram_mem[125484] = 16'b0000000000000000;
	sram_mem[125485] = 16'b0000000000000000;
	sram_mem[125486] = 16'b0000000000000000;
	sram_mem[125487] = 16'b0000000000000000;
	sram_mem[125488] = 16'b0000000000000000;
	sram_mem[125489] = 16'b0000000000000000;
	sram_mem[125490] = 16'b0000000000000000;
	sram_mem[125491] = 16'b0000000000000000;
	sram_mem[125492] = 16'b0000000000000000;
	sram_mem[125493] = 16'b0000000000000000;
	sram_mem[125494] = 16'b0000000000000000;
	sram_mem[125495] = 16'b0000000000000000;
	sram_mem[125496] = 16'b0000000000000000;
	sram_mem[125497] = 16'b0000000000000000;
	sram_mem[125498] = 16'b0000000000000000;
	sram_mem[125499] = 16'b0000000000000000;
	sram_mem[125500] = 16'b0000000000000000;
	sram_mem[125501] = 16'b0000000000000000;
	sram_mem[125502] = 16'b0000000000000000;
	sram_mem[125503] = 16'b0000000000000000;
	sram_mem[125504] = 16'b0000000000000000;
	sram_mem[125505] = 16'b0000000000000000;
	sram_mem[125506] = 16'b0000000000000000;
	sram_mem[125507] = 16'b0000000000000000;
	sram_mem[125508] = 16'b0000000000000000;
	sram_mem[125509] = 16'b0000000000000000;
	sram_mem[125510] = 16'b0000000000000000;
	sram_mem[125511] = 16'b0000000000000000;
	sram_mem[125512] = 16'b0000000000000000;
	sram_mem[125513] = 16'b0000000000000000;
	sram_mem[125514] = 16'b0000000000000000;
	sram_mem[125515] = 16'b0000000000000000;
	sram_mem[125516] = 16'b0000000000000000;
	sram_mem[125517] = 16'b0000000000000000;
	sram_mem[125518] = 16'b0000000000000000;
	sram_mem[125519] = 16'b0000000000000000;
	sram_mem[125520] = 16'b0000000000000000;
	sram_mem[125521] = 16'b0000000000000000;
	sram_mem[125522] = 16'b0000000000000000;
	sram_mem[125523] = 16'b0000000000000000;
	sram_mem[125524] = 16'b0000000000000000;
	sram_mem[125525] = 16'b0000000000000000;
	sram_mem[125526] = 16'b0000000000000000;
	sram_mem[125527] = 16'b0000000000000000;
	sram_mem[125528] = 16'b0000000000000000;
	sram_mem[125529] = 16'b0000000000000000;
	sram_mem[125530] = 16'b0000000000000000;
	sram_mem[125531] = 16'b0000000000000000;
	sram_mem[125532] = 16'b0000000000000000;
	sram_mem[125533] = 16'b0000000000000000;
	sram_mem[125534] = 16'b0000000000000000;
	sram_mem[125535] = 16'b0000000000000000;
	sram_mem[125536] = 16'b0000000000000000;
	sram_mem[125537] = 16'b0000000000000000;
	sram_mem[125538] = 16'b0000000000000000;
	sram_mem[125539] = 16'b0000000000000000;
	sram_mem[125540] = 16'b0000000000000000;
	sram_mem[125541] = 16'b0000000000000000;
	sram_mem[125542] = 16'b0000000000000000;
	sram_mem[125543] = 16'b0000000000000000;
	sram_mem[125544] = 16'b0000000000000000;
	sram_mem[125545] = 16'b0000000000000000;
	sram_mem[125546] = 16'b0000000000000000;
	sram_mem[125547] = 16'b0000000000000000;
	sram_mem[125548] = 16'b0000000000000000;
	sram_mem[125549] = 16'b0000000000000000;
	sram_mem[125550] = 16'b0000000000000000;
	sram_mem[125551] = 16'b0000000000000000;
	sram_mem[125552] = 16'b0000000000000000;
	sram_mem[125553] = 16'b0000000000000000;
	sram_mem[125554] = 16'b0000000000000000;
	sram_mem[125555] = 16'b0000000000000000;
	sram_mem[125556] = 16'b0000000000000000;
	sram_mem[125557] = 16'b0000000000000000;
	sram_mem[125558] = 16'b0000000000000000;
	sram_mem[125559] = 16'b0000000000000000;
	sram_mem[125560] = 16'b0000000000000000;
	sram_mem[125561] = 16'b0000000000000000;
	sram_mem[125562] = 16'b0000000000000000;
	sram_mem[125563] = 16'b0000000000000000;
	sram_mem[125564] = 16'b0000000000000000;
	sram_mem[125565] = 16'b0000000000000000;
	sram_mem[125566] = 16'b0000000000000000;
	sram_mem[125567] = 16'b0000000000000000;
	sram_mem[125568] = 16'b0000000000000000;
	sram_mem[125569] = 16'b0000000000000000;
	sram_mem[125570] = 16'b0000000000000000;
	sram_mem[125571] = 16'b0000000000000000;
	sram_mem[125572] = 16'b0000000000000000;
	sram_mem[125573] = 16'b0000000000000000;
	sram_mem[125574] = 16'b0000000000000000;
	sram_mem[125575] = 16'b0000000000000000;
	sram_mem[125576] = 16'b0000000000000000;
	sram_mem[125577] = 16'b0000000000000000;
	sram_mem[125578] = 16'b0000000000000000;
	sram_mem[125579] = 16'b0000000000000000;
	sram_mem[125580] = 16'b0000000000000000;
	sram_mem[125581] = 16'b0000000000000000;
	sram_mem[125582] = 16'b0000000000000000;
	sram_mem[125583] = 16'b0000000000000000;
	sram_mem[125584] = 16'b0000000000000000;
	sram_mem[125585] = 16'b0000000000000000;
	sram_mem[125586] = 16'b0000000000000000;
	sram_mem[125587] = 16'b0000000000000000;
	sram_mem[125588] = 16'b0000000000000000;
	sram_mem[125589] = 16'b0000000000000000;
	sram_mem[125590] = 16'b0000000000000000;
	sram_mem[125591] = 16'b0000000000000000;
	sram_mem[125592] = 16'b0000000000000000;
	sram_mem[125593] = 16'b0000000000000000;
	sram_mem[125594] = 16'b0000000000000000;
	sram_mem[125595] = 16'b0000000000000000;
	sram_mem[125596] = 16'b0000000000000000;
	sram_mem[125597] = 16'b0000000000000000;
	sram_mem[125598] = 16'b0000000000000000;
	sram_mem[125599] = 16'b0000000000000000;
	sram_mem[125600] = 16'b0000000000000000;
	sram_mem[125601] = 16'b0000000000000000;
	sram_mem[125602] = 16'b0000000000000000;
	sram_mem[125603] = 16'b0000000000000000;
	sram_mem[125604] = 16'b0000000000000000;
	sram_mem[125605] = 16'b0000000000000000;
	sram_mem[125606] = 16'b0000000000000000;
	sram_mem[125607] = 16'b0000000000000000;
	sram_mem[125608] = 16'b0000000000000000;
	sram_mem[125609] = 16'b0000000000000000;
	sram_mem[125610] = 16'b0000000000000000;
	sram_mem[125611] = 16'b0000000000000000;
	sram_mem[125612] = 16'b0000000000000000;
	sram_mem[125613] = 16'b0000000000000000;
	sram_mem[125614] = 16'b0000000000000000;
	sram_mem[125615] = 16'b0000000000000000;
	sram_mem[125616] = 16'b0000000000000000;
	sram_mem[125617] = 16'b0000000000000000;
	sram_mem[125618] = 16'b0000000000000000;
	sram_mem[125619] = 16'b0000000000000000;
	sram_mem[125620] = 16'b0000000000000000;
	sram_mem[125621] = 16'b0000000000000000;
	sram_mem[125622] = 16'b0000000000000000;
	sram_mem[125623] = 16'b0000000000000000;
	sram_mem[125624] = 16'b0000000000000000;
	sram_mem[125625] = 16'b0000000000000000;
	sram_mem[125626] = 16'b0000000000000000;
	sram_mem[125627] = 16'b0000000000000000;
	sram_mem[125628] = 16'b0000000000000000;
	sram_mem[125629] = 16'b0000000000000000;
	sram_mem[125630] = 16'b0000000000000000;
	sram_mem[125631] = 16'b0000000000000000;
	sram_mem[125632] = 16'b0000000000000000;
	sram_mem[125633] = 16'b0000000000000000;
	sram_mem[125634] = 16'b0000000000000000;
	sram_mem[125635] = 16'b0000000000000000;
	sram_mem[125636] = 16'b0000000000000000;
	sram_mem[125637] = 16'b0000000000000000;
	sram_mem[125638] = 16'b0000000000000000;
	sram_mem[125639] = 16'b0000000000000000;
	sram_mem[125640] = 16'b0000000000000000;
	sram_mem[125641] = 16'b0000000000000000;
	sram_mem[125642] = 16'b0000000000000000;
	sram_mem[125643] = 16'b0000000000000000;
	sram_mem[125644] = 16'b0000000000000000;
	sram_mem[125645] = 16'b0000000000000000;
	sram_mem[125646] = 16'b0000000000000000;
	sram_mem[125647] = 16'b0000000000000000;
	sram_mem[125648] = 16'b0000000000000000;
	sram_mem[125649] = 16'b0000000000000000;
	sram_mem[125650] = 16'b0000000000000000;
	sram_mem[125651] = 16'b0000000000000000;
	sram_mem[125652] = 16'b0000000000000000;
	sram_mem[125653] = 16'b0000000000000000;
	sram_mem[125654] = 16'b0000000000000000;
	sram_mem[125655] = 16'b0000000000000000;
	sram_mem[125656] = 16'b0000000000000000;
	sram_mem[125657] = 16'b0000000000000000;
	sram_mem[125658] = 16'b0000000000000000;
	sram_mem[125659] = 16'b0000000000000000;
	sram_mem[125660] = 16'b0000000000000000;
	sram_mem[125661] = 16'b0000000000000000;
	sram_mem[125662] = 16'b0000000000000000;
	sram_mem[125663] = 16'b0000000000000000;
	sram_mem[125664] = 16'b0000000000000000;
	sram_mem[125665] = 16'b0000000000000000;
	sram_mem[125666] = 16'b0000000000000000;
	sram_mem[125667] = 16'b0000000000000000;
	sram_mem[125668] = 16'b0000000000000000;
	sram_mem[125669] = 16'b0000000000000000;
	sram_mem[125670] = 16'b0000000000000000;
	sram_mem[125671] = 16'b0000000000000000;
	sram_mem[125672] = 16'b0000000000000000;
	sram_mem[125673] = 16'b0000000000000000;
	sram_mem[125674] = 16'b0000000000000000;
	sram_mem[125675] = 16'b0000000000000000;
	sram_mem[125676] = 16'b0000000000000000;
	sram_mem[125677] = 16'b0000000000000000;
	sram_mem[125678] = 16'b0000000000000000;
	sram_mem[125679] = 16'b0000000000000000;
	sram_mem[125680] = 16'b0000000000000000;
	sram_mem[125681] = 16'b0000000000000000;
	sram_mem[125682] = 16'b0000000000000000;
	sram_mem[125683] = 16'b0000000000000000;
	sram_mem[125684] = 16'b0000000000000000;
	sram_mem[125685] = 16'b0000000000000000;
	sram_mem[125686] = 16'b0000000000000000;
	sram_mem[125687] = 16'b0000000000000000;
	sram_mem[125688] = 16'b0000000000000000;
	sram_mem[125689] = 16'b0000000000000000;
	sram_mem[125690] = 16'b0000000000000000;
	sram_mem[125691] = 16'b0000000000000000;
	sram_mem[125692] = 16'b0000000000000000;
	sram_mem[125693] = 16'b0000000000000000;
	sram_mem[125694] = 16'b0000000000000000;
	sram_mem[125695] = 16'b0000000000000000;
	sram_mem[125696] = 16'b0000000000000000;
	sram_mem[125697] = 16'b0000000000000000;
	sram_mem[125698] = 16'b0000000000000000;
	sram_mem[125699] = 16'b0000000000000000;
	sram_mem[125700] = 16'b0000000000000000;
	sram_mem[125701] = 16'b0000000000000000;
	sram_mem[125702] = 16'b0000000000000000;
	sram_mem[125703] = 16'b0000000000000000;
	sram_mem[125704] = 16'b0000000000000000;
	sram_mem[125705] = 16'b0000000000000000;
	sram_mem[125706] = 16'b0000000000000000;
	sram_mem[125707] = 16'b0000000000000000;
	sram_mem[125708] = 16'b0000000000000000;
	sram_mem[125709] = 16'b0000000000000000;
	sram_mem[125710] = 16'b0000000000000000;
	sram_mem[125711] = 16'b0000000000000000;
	sram_mem[125712] = 16'b0000000000000000;
	sram_mem[125713] = 16'b0000000000000000;
	sram_mem[125714] = 16'b0000000000000000;
	sram_mem[125715] = 16'b0000000000000000;
	sram_mem[125716] = 16'b0000000000000000;
	sram_mem[125717] = 16'b0000000000000000;
	sram_mem[125718] = 16'b0000000000000000;
	sram_mem[125719] = 16'b0000000000000000;
	sram_mem[125720] = 16'b0000000000000000;
	sram_mem[125721] = 16'b0000000000000000;
	sram_mem[125722] = 16'b0000000000000000;
	sram_mem[125723] = 16'b0000000000000000;
	sram_mem[125724] = 16'b0000000000000000;
	sram_mem[125725] = 16'b0000000000000000;
	sram_mem[125726] = 16'b0000000000000000;
	sram_mem[125727] = 16'b0000000000000000;
	sram_mem[125728] = 16'b0000000000000000;
	sram_mem[125729] = 16'b0000000000000000;
	sram_mem[125730] = 16'b0000000000000000;
	sram_mem[125731] = 16'b0000000000000000;
	sram_mem[125732] = 16'b0000000000000000;
	sram_mem[125733] = 16'b0000000000000000;
	sram_mem[125734] = 16'b0000000000000000;
	sram_mem[125735] = 16'b0000000000000000;
	sram_mem[125736] = 16'b0000000000000000;
	sram_mem[125737] = 16'b0000000000000000;
	sram_mem[125738] = 16'b0000000000000000;
	sram_mem[125739] = 16'b0000000000000000;
	sram_mem[125740] = 16'b0000000000000000;
	sram_mem[125741] = 16'b0000000000000000;
	sram_mem[125742] = 16'b0000000000000000;
	sram_mem[125743] = 16'b0000000000000000;
	sram_mem[125744] = 16'b0000000000000000;
	sram_mem[125745] = 16'b0000000000000000;
	sram_mem[125746] = 16'b0000000000000000;
	sram_mem[125747] = 16'b0000000000000000;
	sram_mem[125748] = 16'b0000000000000000;
	sram_mem[125749] = 16'b0000000000000000;
	sram_mem[125750] = 16'b0000000000000000;
	sram_mem[125751] = 16'b0000000000000000;
	sram_mem[125752] = 16'b0000000000000000;
	sram_mem[125753] = 16'b0000000000000000;
	sram_mem[125754] = 16'b0000000000000000;
	sram_mem[125755] = 16'b0000000000000000;
	sram_mem[125756] = 16'b0000000000000000;
	sram_mem[125757] = 16'b0000000000000000;
	sram_mem[125758] = 16'b0000000000000000;
	sram_mem[125759] = 16'b0000000000000000;
	sram_mem[125760] = 16'b0000000000000000;
	sram_mem[125761] = 16'b0000000000000000;
	sram_mem[125762] = 16'b0000000000000000;
	sram_mem[125763] = 16'b0000000000000000;
	sram_mem[125764] = 16'b0000000000000000;
	sram_mem[125765] = 16'b0000000000000000;
	sram_mem[125766] = 16'b0000000000000000;
	sram_mem[125767] = 16'b0000000000000000;
	sram_mem[125768] = 16'b0000000000000000;
	sram_mem[125769] = 16'b0000000000000000;
	sram_mem[125770] = 16'b0000000000000000;
	sram_mem[125771] = 16'b0000000000000000;
	sram_mem[125772] = 16'b0000000000000000;
	sram_mem[125773] = 16'b0000000000000000;
	sram_mem[125774] = 16'b0000000000000000;
	sram_mem[125775] = 16'b0000000000000000;
	sram_mem[125776] = 16'b0000000000000000;
	sram_mem[125777] = 16'b0000000000000000;
	sram_mem[125778] = 16'b0000000000000000;
	sram_mem[125779] = 16'b0000000000000000;
	sram_mem[125780] = 16'b0000000000000000;
	sram_mem[125781] = 16'b0000000000000000;
	sram_mem[125782] = 16'b0000000000000000;
	sram_mem[125783] = 16'b0000000000000000;
	sram_mem[125784] = 16'b0000000000000000;
	sram_mem[125785] = 16'b0000000000000000;
	sram_mem[125786] = 16'b0000000000000000;
	sram_mem[125787] = 16'b0000000000000000;
	sram_mem[125788] = 16'b0000000000000000;
	sram_mem[125789] = 16'b0000000000000000;
	sram_mem[125790] = 16'b0000000000000000;
	sram_mem[125791] = 16'b0000000000000000;
	sram_mem[125792] = 16'b0000000000000000;
	sram_mem[125793] = 16'b0000000000000000;
	sram_mem[125794] = 16'b0000000000000000;
	sram_mem[125795] = 16'b0000000000000000;
	sram_mem[125796] = 16'b0000000000000000;
	sram_mem[125797] = 16'b0000000000000000;
	sram_mem[125798] = 16'b0000000000000000;
	sram_mem[125799] = 16'b0000000000000000;
	sram_mem[125800] = 16'b0000000000000000;
	sram_mem[125801] = 16'b0000000000000000;
	sram_mem[125802] = 16'b0000000000000000;
	sram_mem[125803] = 16'b0000000000000000;
	sram_mem[125804] = 16'b0000000000000000;
	sram_mem[125805] = 16'b0000000000000000;
	sram_mem[125806] = 16'b0000000000000000;
	sram_mem[125807] = 16'b0000000000000000;
	sram_mem[125808] = 16'b0000000000000000;
	sram_mem[125809] = 16'b0000000000000000;
	sram_mem[125810] = 16'b0000000000000000;
	sram_mem[125811] = 16'b0000000000000000;
	sram_mem[125812] = 16'b0000000000000000;
	sram_mem[125813] = 16'b0000000000000000;
	sram_mem[125814] = 16'b0000000000000000;
	sram_mem[125815] = 16'b0000000000000000;
	sram_mem[125816] = 16'b0000000000000000;
	sram_mem[125817] = 16'b0000000000000000;
	sram_mem[125818] = 16'b0000000000000000;
	sram_mem[125819] = 16'b0000000000000000;
	sram_mem[125820] = 16'b0000000000000000;
	sram_mem[125821] = 16'b0000000000000000;
	sram_mem[125822] = 16'b0000000000000000;
	sram_mem[125823] = 16'b0000000000000000;
	sram_mem[125824] = 16'b0000000000000000;
	sram_mem[125825] = 16'b0000000000000000;
	sram_mem[125826] = 16'b0000000000000000;
	sram_mem[125827] = 16'b0000000000000000;
	sram_mem[125828] = 16'b0000000000000000;
	sram_mem[125829] = 16'b0000000000000000;
	sram_mem[125830] = 16'b0000000000000000;
	sram_mem[125831] = 16'b0000000000000000;
	sram_mem[125832] = 16'b0000000000000000;
	sram_mem[125833] = 16'b0000000000000000;
	sram_mem[125834] = 16'b0000000000000000;
	sram_mem[125835] = 16'b0000000000000000;
	sram_mem[125836] = 16'b0000000000000000;
	sram_mem[125837] = 16'b0000000000000000;
	sram_mem[125838] = 16'b0000000000000000;
	sram_mem[125839] = 16'b0000000000000000;
	sram_mem[125840] = 16'b0000000000000000;
	sram_mem[125841] = 16'b0000000000000000;
	sram_mem[125842] = 16'b0000000000000000;
	sram_mem[125843] = 16'b0000000000000000;
	sram_mem[125844] = 16'b0000000000000000;
	sram_mem[125845] = 16'b0000000000000000;
	sram_mem[125846] = 16'b0000000000000000;
	sram_mem[125847] = 16'b0000000000000000;
	sram_mem[125848] = 16'b0000000000000000;
	sram_mem[125849] = 16'b0000000000000000;
	sram_mem[125850] = 16'b0000000000000000;
	sram_mem[125851] = 16'b0000000000000000;
	sram_mem[125852] = 16'b0000000000000000;
	sram_mem[125853] = 16'b0000000000000000;
	sram_mem[125854] = 16'b0000000000000000;
	sram_mem[125855] = 16'b0000000000000000;
	sram_mem[125856] = 16'b0000000000000000;
	sram_mem[125857] = 16'b0000000000000000;
	sram_mem[125858] = 16'b0000000000000000;
	sram_mem[125859] = 16'b0000000000000000;
	sram_mem[125860] = 16'b0000000000000000;
	sram_mem[125861] = 16'b0000000000000000;
	sram_mem[125862] = 16'b0000000000000000;
	sram_mem[125863] = 16'b0000000000000000;
	sram_mem[125864] = 16'b0000000000000000;
	sram_mem[125865] = 16'b0000000000000000;
	sram_mem[125866] = 16'b0000000000000000;
	sram_mem[125867] = 16'b0000000000000000;
	sram_mem[125868] = 16'b0000000000000000;
	sram_mem[125869] = 16'b0000000000000000;
	sram_mem[125870] = 16'b0000000000000000;
	sram_mem[125871] = 16'b0000000000000000;
	sram_mem[125872] = 16'b0000000000000000;
	sram_mem[125873] = 16'b0000000000000000;
	sram_mem[125874] = 16'b0000000000000000;
	sram_mem[125875] = 16'b0000000000000000;
	sram_mem[125876] = 16'b0000000000000000;
	sram_mem[125877] = 16'b0000000000000000;
	sram_mem[125878] = 16'b0000000000000000;
	sram_mem[125879] = 16'b0000000000000000;
	sram_mem[125880] = 16'b0000000000000000;
	sram_mem[125881] = 16'b0000000000000000;
	sram_mem[125882] = 16'b0000000000000000;
	sram_mem[125883] = 16'b0000000000000000;
	sram_mem[125884] = 16'b0000000000000000;
	sram_mem[125885] = 16'b0000000000000000;
	sram_mem[125886] = 16'b0000000000000000;
	sram_mem[125887] = 16'b0000000000000000;
	sram_mem[125888] = 16'b0000000000000000;
	sram_mem[125889] = 16'b0000000000000000;
	sram_mem[125890] = 16'b0000000000000000;
	sram_mem[125891] = 16'b0000000000000000;
	sram_mem[125892] = 16'b0000000000000000;
	sram_mem[125893] = 16'b0000000000000000;
	sram_mem[125894] = 16'b0000000000000000;
	sram_mem[125895] = 16'b0000000000000000;
	sram_mem[125896] = 16'b0000000000000000;
	sram_mem[125897] = 16'b0000000000000000;
	sram_mem[125898] = 16'b0000000000000000;
	sram_mem[125899] = 16'b0000000000000000;
	sram_mem[125900] = 16'b0000000000000000;
	sram_mem[125901] = 16'b0000000000000000;
	sram_mem[125902] = 16'b0000000000000000;
	sram_mem[125903] = 16'b0000000000000000;
	sram_mem[125904] = 16'b0000000000000000;
	sram_mem[125905] = 16'b0000000000000000;
	sram_mem[125906] = 16'b0000000000000000;
	sram_mem[125907] = 16'b0000000000000000;
	sram_mem[125908] = 16'b0000000000000000;
	sram_mem[125909] = 16'b0000000000000000;
	sram_mem[125910] = 16'b0000000000000000;
	sram_mem[125911] = 16'b0000000000000000;
	sram_mem[125912] = 16'b0000000000000000;
	sram_mem[125913] = 16'b0000000000000000;
	sram_mem[125914] = 16'b0000000000000000;
	sram_mem[125915] = 16'b0000000000000000;
	sram_mem[125916] = 16'b0000000000000000;
	sram_mem[125917] = 16'b0000000000000000;
	sram_mem[125918] = 16'b0000000000000000;
	sram_mem[125919] = 16'b0000000000000000;
	sram_mem[125920] = 16'b0000000000000000;
	sram_mem[125921] = 16'b0000000000000000;
	sram_mem[125922] = 16'b0000000000000000;
	sram_mem[125923] = 16'b0000000000000000;
	sram_mem[125924] = 16'b0000000000000000;
	sram_mem[125925] = 16'b0000000000000000;
	sram_mem[125926] = 16'b0000000000000000;
	sram_mem[125927] = 16'b0000000000000000;
	sram_mem[125928] = 16'b0000000000000000;
	sram_mem[125929] = 16'b0000000000000000;
	sram_mem[125930] = 16'b0000000000000000;
	sram_mem[125931] = 16'b0000000000000000;
	sram_mem[125932] = 16'b0000000000000000;
	sram_mem[125933] = 16'b0000000000000000;
	sram_mem[125934] = 16'b0000000000000000;
	sram_mem[125935] = 16'b0000000000000000;
	sram_mem[125936] = 16'b0000000000000000;
	sram_mem[125937] = 16'b0000000000000000;
	sram_mem[125938] = 16'b0000000000000000;
	sram_mem[125939] = 16'b0000000000000000;
	sram_mem[125940] = 16'b0000000000000000;
	sram_mem[125941] = 16'b0000000000000000;
	sram_mem[125942] = 16'b0000000000000000;
	sram_mem[125943] = 16'b0000000000000000;
	sram_mem[125944] = 16'b0000000000000000;
	sram_mem[125945] = 16'b0000000000000000;
	sram_mem[125946] = 16'b0000000000000000;
	sram_mem[125947] = 16'b0000000000000000;
	sram_mem[125948] = 16'b0000000000000000;
	sram_mem[125949] = 16'b0000000000000000;
	sram_mem[125950] = 16'b0000000000000000;
	sram_mem[125951] = 16'b0000000000000000;
	sram_mem[125952] = 16'b0000000000000000;
	sram_mem[125953] = 16'b0000000000000000;
	sram_mem[125954] = 16'b0000000000000000;
	sram_mem[125955] = 16'b0000000000000000;
	sram_mem[125956] = 16'b0000000000000000;
	sram_mem[125957] = 16'b0000000000000000;
	sram_mem[125958] = 16'b0000000000000000;
	sram_mem[125959] = 16'b0000000000000000;
	sram_mem[125960] = 16'b0000000000000000;
	sram_mem[125961] = 16'b0000000000000000;
	sram_mem[125962] = 16'b0000000000000000;
	sram_mem[125963] = 16'b0000000000000000;
	sram_mem[125964] = 16'b0000000000000000;
	sram_mem[125965] = 16'b0000000000000000;
	sram_mem[125966] = 16'b0000000000000000;
	sram_mem[125967] = 16'b0000000000000000;
	sram_mem[125968] = 16'b0000000000000000;
	sram_mem[125969] = 16'b0000000000000000;
	sram_mem[125970] = 16'b0000000000000000;
	sram_mem[125971] = 16'b0000000000000000;
	sram_mem[125972] = 16'b0000000000000000;
	sram_mem[125973] = 16'b0000000000000000;
	sram_mem[125974] = 16'b0000000000000000;
	sram_mem[125975] = 16'b0000000000000000;
	sram_mem[125976] = 16'b0000000000000000;
	sram_mem[125977] = 16'b0000000000000000;
	sram_mem[125978] = 16'b0000000000000000;
	sram_mem[125979] = 16'b0000000000000000;
	sram_mem[125980] = 16'b0000000000000000;
	sram_mem[125981] = 16'b0000000000000000;
	sram_mem[125982] = 16'b0000000000000000;
	sram_mem[125983] = 16'b0000000000000000;
	sram_mem[125984] = 16'b0000000000000000;
	sram_mem[125985] = 16'b0000000000000000;
	sram_mem[125986] = 16'b0000000000000000;
	sram_mem[125987] = 16'b0000000000000000;
	sram_mem[125988] = 16'b0000000000000000;
	sram_mem[125989] = 16'b0000000000000000;
	sram_mem[125990] = 16'b0000000000000000;
	sram_mem[125991] = 16'b0000000000000000;
	sram_mem[125992] = 16'b0000000000000000;
	sram_mem[125993] = 16'b0000000000000000;
	sram_mem[125994] = 16'b0000000000000000;
	sram_mem[125995] = 16'b0000000000000000;
	sram_mem[125996] = 16'b0000000000000000;
	sram_mem[125997] = 16'b0000000000000000;
	sram_mem[125998] = 16'b0000000000000000;
	sram_mem[125999] = 16'b0000000000000000;
	sram_mem[126000] = 16'b0000000000000000;
	sram_mem[126001] = 16'b0000000000000000;
	sram_mem[126002] = 16'b0000000000000000;
	sram_mem[126003] = 16'b0000000000000000;
	sram_mem[126004] = 16'b0000000000000000;
	sram_mem[126005] = 16'b0000000000000000;
	sram_mem[126006] = 16'b0000000000000000;
	sram_mem[126007] = 16'b0000000000000000;
	sram_mem[126008] = 16'b0000000000000000;
	sram_mem[126009] = 16'b0000000000000000;
	sram_mem[126010] = 16'b0000000000000000;
	sram_mem[126011] = 16'b0000000000000000;
	sram_mem[126012] = 16'b0000000000000000;
	sram_mem[126013] = 16'b0000000000000000;
	sram_mem[126014] = 16'b0000000000000000;
	sram_mem[126015] = 16'b0000000000000000;
	sram_mem[126016] = 16'b0000000000000000;
	sram_mem[126017] = 16'b0000000000000000;
	sram_mem[126018] = 16'b0000000000000000;
	sram_mem[126019] = 16'b0000000000000000;
	sram_mem[126020] = 16'b0000000000000000;
	sram_mem[126021] = 16'b0000000000000000;
	sram_mem[126022] = 16'b0000000000000000;
	sram_mem[126023] = 16'b0000000000000000;
	sram_mem[126024] = 16'b0000000000000000;
	sram_mem[126025] = 16'b0000000000000000;
	sram_mem[126026] = 16'b0000000000000000;
	sram_mem[126027] = 16'b0000000000000000;
	sram_mem[126028] = 16'b0000000000000000;
	sram_mem[126029] = 16'b0000000000000000;
	sram_mem[126030] = 16'b0000000000000000;
	sram_mem[126031] = 16'b0000000000000000;
	sram_mem[126032] = 16'b0000000000000000;
	sram_mem[126033] = 16'b0000000000000000;
	sram_mem[126034] = 16'b0000000000000000;
	sram_mem[126035] = 16'b0000000000000000;
	sram_mem[126036] = 16'b0000000000000000;
	sram_mem[126037] = 16'b0000000000000000;
	sram_mem[126038] = 16'b0000000000000000;
	sram_mem[126039] = 16'b0000000000000000;
	sram_mem[126040] = 16'b0000000000000000;
	sram_mem[126041] = 16'b0000000000000000;
	sram_mem[126042] = 16'b0000000000000000;
	sram_mem[126043] = 16'b0000000000000000;
	sram_mem[126044] = 16'b0000000000000000;
	sram_mem[126045] = 16'b0000000000000000;
	sram_mem[126046] = 16'b0000000000000000;
	sram_mem[126047] = 16'b0000000000000000;
	sram_mem[126048] = 16'b0000000000000000;
	sram_mem[126049] = 16'b0000000000000000;
	sram_mem[126050] = 16'b0000000000000000;
	sram_mem[126051] = 16'b0000000000000000;
	sram_mem[126052] = 16'b0000000000000000;
	sram_mem[126053] = 16'b0000000000000000;
	sram_mem[126054] = 16'b0000000000000000;
	sram_mem[126055] = 16'b0000000000000000;
	sram_mem[126056] = 16'b0000000000000000;
	sram_mem[126057] = 16'b0000000000000000;
	sram_mem[126058] = 16'b0000000000000000;
	sram_mem[126059] = 16'b0000000000000000;
	sram_mem[126060] = 16'b0000000000000000;
	sram_mem[126061] = 16'b0000000000000000;
	sram_mem[126062] = 16'b0000000000000000;
	sram_mem[126063] = 16'b0000000000000000;
	sram_mem[126064] = 16'b0000000000000000;
	sram_mem[126065] = 16'b0000000000000000;
	sram_mem[126066] = 16'b0000000000000000;
	sram_mem[126067] = 16'b0000000000000000;
	sram_mem[126068] = 16'b0000000000000000;
	sram_mem[126069] = 16'b0000000000000000;
	sram_mem[126070] = 16'b0000000000000000;
	sram_mem[126071] = 16'b0000000000000000;
	sram_mem[126072] = 16'b0000000000000000;
	sram_mem[126073] = 16'b0000000000000000;
	sram_mem[126074] = 16'b0000000000000000;
	sram_mem[126075] = 16'b0000000000000000;
	sram_mem[126076] = 16'b0000000000000000;
	sram_mem[126077] = 16'b0000000000000000;
	sram_mem[126078] = 16'b0000000000000000;
	sram_mem[126079] = 16'b0000000000000000;
	sram_mem[126080] = 16'b0000000000000000;
	sram_mem[126081] = 16'b0000000000000000;
	sram_mem[126082] = 16'b0000000000000000;
	sram_mem[126083] = 16'b0000000000000000;
	sram_mem[126084] = 16'b0000000000000000;
	sram_mem[126085] = 16'b0000000000000000;
	sram_mem[126086] = 16'b0000000000000000;
	sram_mem[126087] = 16'b0000000000000000;
	sram_mem[126088] = 16'b0000000000000000;
	sram_mem[126089] = 16'b0000000000000000;
	sram_mem[126090] = 16'b0000000000000000;
	sram_mem[126091] = 16'b0000000000000000;
	sram_mem[126092] = 16'b0000000000000000;
	sram_mem[126093] = 16'b0000000000000000;
	sram_mem[126094] = 16'b0000000000000000;
	sram_mem[126095] = 16'b0000000000000000;
	sram_mem[126096] = 16'b0000000000000000;
	sram_mem[126097] = 16'b0000000000000000;
	sram_mem[126098] = 16'b0000000000000000;
	sram_mem[126099] = 16'b0000000000000000;
	sram_mem[126100] = 16'b0000000000000000;
	sram_mem[126101] = 16'b0000000000000000;
	sram_mem[126102] = 16'b0000000000000000;
	sram_mem[126103] = 16'b0000000000000000;
	sram_mem[126104] = 16'b0000000000000000;
	sram_mem[126105] = 16'b0000000000000000;
	sram_mem[126106] = 16'b0000000000000000;
	sram_mem[126107] = 16'b0000000000000000;
	sram_mem[126108] = 16'b0000000000000000;
	sram_mem[126109] = 16'b0000000000000000;
	sram_mem[126110] = 16'b0000000000000000;
	sram_mem[126111] = 16'b0000000000000000;
	sram_mem[126112] = 16'b0000000000000000;
	sram_mem[126113] = 16'b0000000000000000;
	sram_mem[126114] = 16'b0000000000000000;
	sram_mem[126115] = 16'b0000000000000000;
	sram_mem[126116] = 16'b0000000000000000;
	sram_mem[126117] = 16'b0000000000000000;
	sram_mem[126118] = 16'b0000000000000000;
	sram_mem[126119] = 16'b0000000000000000;
	sram_mem[126120] = 16'b0000000000000000;
	sram_mem[126121] = 16'b0000000000000000;
	sram_mem[126122] = 16'b0000000000000000;
	sram_mem[126123] = 16'b0000000000000000;
	sram_mem[126124] = 16'b0000000000000000;
	sram_mem[126125] = 16'b0000000000000000;
	sram_mem[126126] = 16'b0000000000000000;
	sram_mem[126127] = 16'b0000000000000000;
	sram_mem[126128] = 16'b0000000000000000;
	sram_mem[126129] = 16'b0000000000000000;
	sram_mem[126130] = 16'b0000000000000000;
	sram_mem[126131] = 16'b0000000000000000;
	sram_mem[126132] = 16'b0000000000000000;
	sram_mem[126133] = 16'b0000000000000000;
	sram_mem[126134] = 16'b0000000000000000;
	sram_mem[126135] = 16'b0000000000000000;
	sram_mem[126136] = 16'b0000000000000000;
	sram_mem[126137] = 16'b0000000000000000;
	sram_mem[126138] = 16'b0000000000000000;
	sram_mem[126139] = 16'b0000000000000000;
	sram_mem[126140] = 16'b0000000000000000;
	sram_mem[126141] = 16'b0000000000000000;
	sram_mem[126142] = 16'b0000000000000000;
	sram_mem[126143] = 16'b0000000000000000;
	sram_mem[126144] = 16'b0000000000000000;
	sram_mem[126145] = 16'b0000000000000000;
	sram_mem[126146] = 16'b0000000000000000;
	sram_mem[126147] = 16'b0000000000000000;
	sram_mem[126148] = 16'b0000000000000000;
	sram_mem[126149] = 16'b0000000000000000;
	sram_mem[126150] = 16'b0000000000000000;
	sram_mem[126151] = 16'b0000000000000000;
	sram_mem[126152] = 16'b0000000000000000;
	sram_mem[126153] = 16'b0000000000000000;
	sram_mem[126154] = 16'b0000000000000000;
	sram_mem[126155] = 16'b0000000000000000;
	sram_mem[126156] = 16'b0000000000000000;
	sram_mem[126157] = 16'b0000000000000000;
	sram_mem[126158] = 16'b0000000000000000;
	sram_mem[126159] = 16'b0000000000000000;
	sram_mem[126160] = 16'b0000000000000000;
	sram_mem[126161] = 16'b0000000000000000;
	sram_mem[126162] = 16'b0000000000000000;
	sram_mem[126163] = 16'b0000000000000000;
	sram_mem[126164] = 16'b0000000000000000;
	sram_mem[126165] = 16'b0000000000000000;
	sram_mem[126166] = 16'b0000000000000000;
	sram_mem[126167] = 16'b0000000000000000;
	sram_mem[126168] = 16'b0000000000000000;
	sram_mem[126169] = 16'b0000000000000000;
	sram_mem[126170] = 16'b0000000000000000;
	sram_mem[126171] = 16'b0000000000000000;
	sram_mem[126172] = 16'b0000000000000000;
	sram_mem[126173] = 16'b0000000000000000;
	sram_mem[126174] = 16'b0000000000000000;
	sram_mem[126175] = 16'b0000000000000000;
	sram_mem[126176] = 16'b0000000000000000;
	sram_mem[126177] = 16'b0000000000000000;
	sram_mem[126178] = 16'b0000000000000000;
	sram_mem[126179] = 16'b0000000000000000;
	sram_mem[126180] = 16'b0000000000000000;
	sram_mem[126181] = 16'b0000000000000000;
	sram_mem[126182] = 16'b0000000000000000;
	sram_mem[126183] = 16'b0000000000000000;
	sram_mem[126184] = 16'b0000000000000000;
	sram_mem[126185] = 16'b0000000000000000;
	sram_mem[126186] = 16'b0000000000000000;
	sram_mem[126187] = 16'b0000000000000000;
	sram_mem[126188] = 16'b0000000000000000;
	sram_mem[126189] = 16'b0000000000000000;
	sram_mem[126190] = 16'b0000000000000000;
	sram_mem[126191] = 16'b0000000000000000;
	sram_mem[126192] = 16'b0000000000000000;
	sram_mem[126193] = 16'b0000000000000000;
	sram_mem[126194] = 16'b0000000000000000;
	sram_mem[126195] = 16'b0000000000000000;
	sram_mem[126196] = 16'b0000000000000000;
	sram_mem[126197] = 16'b0000000000000000;
	sram_mem[126198] = 16'b0000000000000000;
	sram_mem[126199] = 16'b0000000000000000;
	sram_mem[126200] = 16'b0000000000000000;
	sram_mem[126201] = 16'b0000000000000000;
	sram_mem[126202] = 16'b0000000000000000;
	sram_mem[126203] = 16'b0000000000000000;
	sram_mem[126204] = 16'b0000000000000000;
	sram_mem[126205] = 16'b0000000000000000;
	sram_mem[126206] = 16'b0000000000000000;
	sram_mem[126207] = 16'b0000000000000000;
	sram_mem[126208] = 16'b0000000000000000;
	sram_mem[126209] = 16'b0000000000000000;
	sram_mem[126210] = 16'b0000000000000000;
	sram_mem[126211] = 16'b0000000000000000;
	sram_mem[126212] = 16'b0000000000000000;
	sram_mem[126213] = 16'b0000000000000000;
	sram_mem[126214] = 16'b0000000000000000;
	sram_mem[126215] = 16'b0000000000000000;
	sram_mem[126216] = 16'b0000000000000000;
	sram_mem[126217] = 16'b0000000000000000;
	sram_mem[126218] = 16'b0000000000000000;
	sram_mem[126219] = 16'b0000000000000000;
	sram_mem[126220] = 16'b0000000000000000;
	sram_mem[126221] = 16'b0000000000000000;
	sram_mem[126222] = 16'b0000000000000000;
	sram_mem[126223] = 16'b0000000000000000;
	sram_mem[126224] = 16'b0000000000000000;
	sram_mem[126225] = 16'b0000000000000000;
	sram_mem[126226] = 16'b0000000000000000;
	sram_mem[126227] = 16'b0000000000000000;
	sram_mem[126228] = 16'b0000000000000000;
	sram_mem[126229] = 16'b0000000000000000;
	sram_mem[126230] = 16'b0000000000000000;
	sram_mem[126231] = 16'b0000000000000000;
	sram_mem[126232] = 16'b0000000000000000;
	sram_mem[126233] = 16'b0000000000000000;
	sram_mem[126234] = 16'b0000000000000000;
	sram_mem[126235] = 16'b0000000000000000;
	sram_mem[126236] = 16'b0000000000000000;
	sram_mem[126237] = 16'b0000000000000000;
	sram_mem[126238] = 16'b0000000000000000;
	sram_mem[126239] = 16'b0000000000000000;
	sram_mem[126240] = 16'b0000000000000000;
	sram_mem[126241] = 16'b0000000000000000;
	sram_mem[126242] = 16'b0000000000000000;
	sram_mem[126243] = 16'b0000000000000000;
	sram_mem[126244] = 16'b0000000000000000;
	sram_mem[126245] = 16'b0000000000000000;
	sram_mem[126246] = 16'b0000000000000000;
	sram_mem[126247] = 16'b0000000000000000;
	sram_mem[126248] = 16'b0000000000000000;
	sram_mem[126249] = 16'b0000000000000000;
	sram_mem[126250] = 16'b0000000000000000;
	sram_mem[126251] = 16'b0000000000000000;
	sram_mem[126252] = 16'b0000000000000000;
	sram_mem[126253] = 16'b0000000000000000;
	sram_mem[126254] = 16'b0000000000000000;
	sram_mem[126255] = 16'b0000000000000000;
	sram_mem[126256] = 16'b0000000000000000;
	sram_mem[126257] = 16'b0000000000000000;
	sram_mem[126258] = 16'b0000000000000000;
	sram_mem[126259] = 16'b0000000000000000;
	sram_mem[126260] = 16'b0000000000000000;
	sram_mem[126261] = 16'b0000000000000000;
	sram_mem[126262] = 16'b0000000000000000;
	sram_mem[126263] = 16'b0000000000000000;
	sram_mem[126264] = 16'b0000000000000000;
	sram_mem[126265] = 16'b0000000000000000;
	sram_mem[126266] = 16'b0000000000000000;
	sram_mem[126267] = 16'b0000000000000000;
	sram_mem[126268] = 16'b0000000000000000;
	sram_mem[126269] = 16'b0000000000000000;
	sram_mem[126270] = 16'b0000000000000000;
	sram_mem[126271] = 16'b0000000000000000;
	sram_mem[126272] = 16'b0000000000000000;
	sram_mem[126273] = 16'b0000000000000000;
	sram_mem[126274] = 16'b0000000000000000;
	sram_mem[126275] = 16'b0000000000000000;
	sram_mem[126276] = 16'b0000000000000000;
	sram_mem[126277] = 16'b0000000000000000;
	sram_mem[126278] = 16'b0000000000000000;
	sram_mem[126279] = 16'b0000000000000000;
	sram_mem[126280] = 16'b0000000000000000;
	sram_mem[126281] = 16'b0000000000000000;
	sram_mem[126282] = 16'b0000000000000000;
	sram_mem[126283] = 16'b0000000000000000;
	sram_mem[126284] = 16'b0000000000000000;
	sram_mem[126285] = 16'b0000000000000000;
	sram_mem[126286] = 16'b0000000000000000;
	sram_mem[126287] = 16'b0000000000000000;
	sram_mem[126288] = 16'b0000000000000000;
	sram_mem[126289] = 16'b0000000000000000;
	sram_mem[126290] = 16'b0000000000000000;
	sram_mem[126291] = 16'b0000000000000000;
	sram_mem[126292] = 16'b0000000000000000;
	sram_mem[126293] = 16'b0000000000000000;
	sram_mem[126294] = 16'b0000000000000000;
	sram_mem[126295] = 16'b0000000000000000;
	sram_mem[126296] = 16'b0000000000000000;
	sram_mem[126297] = 16'b0000000000000000;
	sram_mem[126298] = 16'b0000000000000000;
	sram_mem[126299] = 16'b0000000000000000;
	sram_mem[126300] = 16'b0000000000000000;
	sram_mem[126301] = 16'b0000000000000000;
	sram_mem[126302] = 16'b0000000000000000;
	sram_mem[126303] = 16'b0000000000000000;
	sram_mem[126304] = 16'b0000000000000000;
	sram_mem[126305] = 16'b0000000000000000;
	sram_mem[126306] = 16'b0000000000000000;
	sram_mem[126307] = 16'b0000000000000000;
	sram_mem[126308] = 16'b0000000000000000;
	sram_mem[126309] = 16'b0000000000000000;
	sram_mem[126310] = 16'b0000000000000000;
	sram_mem[126311] = 16'b0000000000000000;
	sram_mem[126312] = 16'b0000000000000000;
	sram_mem[126313] = 16'b0000000000000000;
	sram_mem[126314] = 16'b0000000000000000;
	sram_mem[126315] = 16'b0000000000000000;
	sram_mem[126316] = 16'b0000000000000000;
	sram_mem[126317] = 16'b0000000000000000;
	sram_mem[126318] = 16'b0000000000000000;
	sram_mem[126319] = 16'b0000000000000000;
	sram_mem[126320] = 16'b0000000000000000;
	sram_mem[126321] = 16'b0000000000000000;
	sram_mem[126322] = 16'b0000000000000000;
	sram_mem[126323] = 16'b0000000000000000;
	sram_mem[126324] = 16'b0000000000000000;
	sram_mem[126325] = 16'b0000000000000000;
	sram_mem[126326] = 16'b0000000000000000;
	sram_mem[126327] = 16'b0000000000000000;
	sram_mem[126328] = 16'b0000000000000000;
	sram_mem[126329] = 16'b0000000000000000;
	sram_mem[126330] = 16'b0000000000000000;
	sram_mem[126331] = 16'b0000000000000000;
	sram_mem[126332] = 16'b0000000000000000;
	sram_mem[126333] = 16'b0000000000000000;
	sram_mem[126334] = 16'b0000000000000000;
	sram_mem[126335] = 16'b0000000000000000;
	sram_mem[126336] = 16'b0000000000000000;
	sram_mem[126337] = 16'b0000000000000000;
	sram_mem[126338] = 16'b0000000000000000;
	sram_mem[126339] = 16'b0000000000000000;
	sram_mem[126340] = 16'b0000000000000000;
	sram_mem[126341] = 16'b0000000000000000;
	sram_mem[126342] = 16'b0000000000000000;
	sram_mem[126343] = 16'b0000000000000000;
	sram_mem[126344] = 16'b0000000000000000;
	sram_mem[126345] = 16'b0000000000000000;
	sram_mem[126346] = 16'b0000000000000000;
	sram_mem[126347] = 16'b0000000000000000;
	sram_mem[126348] = 16'b0000000000000000;
	sram_mem[126349] = 16'b0000000000000000;
	sram_mem[126350] = 16'b0000000000000000;
	sram_mem[126351] = 16'b0000000000000000;
	sram_mem[126352] = 16'b0000000000000000;
	sram_mem[126353] = 16'b0000000000000000;
	sram_mem[126354] = 16'b0000000000000000;
	sram_mem[126355] = 16'b0000000000000000;
	sram_mem[126356] = 16'b0000000000000000;
	sram_mem[126357] = 16'b0000000000000000;
	sram_mem[126358] = 16'b0000000000000000;
	sram_mem[126359] = 16'b0000000000000000;
	sram_mem[126360] = 16'b0000000000000000;
	sram_mem[126361] = 16'b0000000000000000;
	sram_mem[126362] = 16'b0000000000000000;
	sram_mem[126363] = 16'b0000000000000000;
	sram_mem[126364] = 16'b0000000000000000;
	sram_mem[126365] = 16'b0000000000000000;
	sram_mem[126366] = 16'b0000000000000000;
	sram_mem[126367] = 16'b0000000000000000;
	sram_mem[126368] = 16'b0000000000000000;
	sram_mem[126369] = 16'b0000000000000000;
	sram_mem[126370] = 16'b0000000000000000;
	sram_mem[126371] = 16'b0000000000000000;
	sram_mem[126372] = 16'b0000000000000000;
	sram_mem[126373] = 16'b0000000000000000;
	sram_mem[126374] = 16'b0000000000000000;
	sram_mem[126375] = 16'b0000000000000000;
	sram_mem[126376] = 16'b0000000000000000;
	sram_mem[126377] = 16'b0000000000000000;
	sram_mem[126378] = 16'b0000000000000000;
	sram_mem[126379] = 16'b0000000000000000;
	sram_mem[126380] = 16'b0000000000000000;
	sram_mem[126381] = 16'b0000000000000000;
	sram_mem[126382] = 16'b0000000000000000;
	sram_mem[126383] = 16'b0000000000000000;
	sram_mem[126384] = 16'b0000000000000000;
	sram_mem[126385] = 16'b0000000000000000;
	sram_mem[126386] = 16'b0000000000000000;
	sram_mem[126387] = 16'b0000000000000000;
	sram_mem[126388] = 16'b0000000000000000;
	sram_mem[126389] = 16'b0000000000000000;
	sram_mem[126390] = 16'b0000000000000000;
	sram_mem[126391] = 16'b0000000000000000;
	sram_mem[126392] = 16'b0000000000000000;
	sram_mem[126393] = 16'b0000000000000000;
	sram_mem[126394] = 16'b0000000000000000;
	sram_mem[126395] = 16'b0000000000000000;
	sram_mem[126396] = 16'b0000000000000000;
	sram_mem[126397] = 16'b0000000000000000;
	sram_mem[126398] = 16'b0000000000000000;
	sram_mem[126399] = 16'b0000000000000000;
	sram_mem[126400] = 16'b0000000000000000;
	sram_mem[126401] = 16'b0000000000000000;
	sram_mem[126402] = 16'b0000000000000000;
	sram_mem[126403] = 16'b0000000000000000;
	sram_mem[126404] = 16'b0000000000000000;
	sram_mem[126405] = 16'b0000000000000000;
	sram_mem[126406] = 16'b0000000000000000;
	sram_mem[126407] = 16'b0000000000000000;
	sram_mem[126408] = 16'b0000000000000000;
	sram_mem[126409] = 16'b0000000000000000;
	sram_mem[126410] = 16'b0000000000000000;
	sram_mem[126411] = 16'b0000000000000000;
	sram_mem[126412] = 16'b0000000000000000;
	sram_mem[126413] = 16'b0000000000000000;
	sram_mem[126414] = 16'b0000000000000000;
	sram_mem[126415] = 16'b0000000000000000;
	sram_mem[126416] = 16'b0000000000000000;
	sram_mem[126417] = 16'b0000000000000000;
	sram_mem[126418] = 16'b0000000000000000;
	sram_mem[126419] = 16'b0000000000000000;
	sram_mem[126420] = 16'b0000000000000000;
	sram_mem[126421] = 16'b0000000000000000;
	sram_mem[126422] = 16'b0000000000000000;
	sram_mem[126423] = 16'b0000000000000000;
	sram_mem[126424] = 16'b0000000000000000;
	sram_mem[126425] = 16'b0000000000000000;
	sram_mem[126426] = 16'b0000000000000000;
	sram_mem[126427] = 16'b0000000000000000;
	sram_mem[126428] = 16'b0000000000000000;
	sram_mem[126429] = 16'b0000000000000000;
	sram_mem[126430] = 16'b0000000000000000;
	sram_mem[126431] = 16'b0000000000000000;
	sram_mem[126432] = 16'b0000000000000000;
	sram_mem[126433] = 16'b0000000000000000;
	sram_mem[126434] = 16'b0000000000000000;
	sram_mem[126435] = 16'b0000000000000000;
	sram_mem[126436] = 16'b0000000000000000;
	sram_mem[126437] = 16'b0000000000000000;
	sram_mem[126438] = 16'b0000000000000000;
	sram_mem[126439] = 16'b0000000000000000;
	sram_mem[126440] = 16'b0000000000000000;
	sram_mem[126441] = 16'b0000000000000000;
	sram_mem[126442] = 16'b0000000000000000;
	sram_mem[126443] = 16'b0000000000000000;
	sram_mem[126444] = 16'b0000000000000000;
	sram_mem[126445] = 16'b0000000000000000;
	sram_mem[126446] = 16'b0000000000000000;
	sram_mem[126447] = 16'b0000000000000000;
	sram_mem[126448] = 16'b0000000000000000;
	sram_mem[126449] = 16'b0000000000000000;
	sram_mem[126450] = 16'b0000000000000000;
	sram_mem[126451] = 16'b0000000000000000;
	sram_mem[126452] = 16'b0000000000000000;
	sram_mem[126453] = 16'b0000000000000000;
	sram_mem[126454] = 16'b0000000000000000;
	sram_mem[126455] = 16'b0000000000000000;
	sram_mem[126456] = 16'b0000000000000000;
	sram_mem[126457] = 16'b0000000000000000;
	sram_mem[126458] = 16'b0000000000000000;
	sram_mem[126459] = 16'b0000000000000000;
	sram_mem[126460] = 16'b0000000000000000;
	sram_mem[126461] = 16'b0000000000000000;
	sram_mem[126462] = 16'b0000000000000000;
	sram_mem[126463] = 16'b0000000000000000;
	sram_mem[126464] = 16'b0000000000000000;
	sram_mem[126465] = 16'b0000000000000000;
	sram_mem[126466] = 16'b0000000000000000;
	sram_mem[126467] = 16'b0000000000000000;
	sram_mem[126468] = 16'b0000000000000000;
	sram_mem[126469] = 16'b0000000000000000;
	sram_mem[126470] = 16'b0000000000000000;
	sram_mem[126471] = 16'b0000000000000000;
	sram_mem[126472] = 16'b0000000000000000;
	sram_mem[126473] = 16'b0000000000000000;
	sram_mem[126474] = 16'b0000000000000000;
	sram_mem[126475] = 16'b0000000000000000;
	sram_mem[126476] = 16'b0000000000000000;
	sram_mem[126477] = 16'b0000000000000000;
	sram_mem[126478] = 16'b0000000000000000;
	sram_mem[126479] = 16'b0000000000000000;
	sram_mem[126480] = 16'b0000000000000000;
	sram_mem[126481] = 16'b0000000000000000;
	sram_mem[126482] = 16'b0000000000000000;
	sram_mem[126483] = 16'b0000000000000000;
	sram_mem[126484] = 16'b0000000000000000;
	sram_mem[126485] = 16'b0000000000000000;
	sram_mem[126486] = 16'b0000000000000000;
	sram_mem[126487] = 16'b0000000000000000;
	sram_mem[126488] = 16'b0000000000000000;
	sram_mem[126489] = 16'b0000000000000000;
	sram_mem[126490] = 16'b0000000000000000;
	sram_mem[126491] = 16'b0000000000000000;
	sram_mem[126492] = 16'b0000000000000000;
	sram_mem[126493] = 16'b0000000000000000;
	sram_mem[126494] = 16'b0000000000000000;
	sram_mem[126495] = 16'b0000000000000000;
	sram_mem[126496] = 16'b0000000000000000;
	sram_mem[126497] = 16'b0000000000000000;
	sram_mem[126498] = 16'b0000000000000000;
	sram_mem[126499] = 16'b0000000000000000;
	sram_mem[126500] = 16'b0000000000000000;
	sram_mem[126501] = 16'b0000000000000000;
	sram_mem[126502] = 16'b0000000000000000;
	sram_mem[126503] = 16'b0000000000000000;
	sram_mem[126504] = 16'b0000000000000000;
	sram_mem[126505] = 16'b0000000000000000;
	sram_mem[126506] = 16'b0000000000000000;
	sram_mem[126507] = 16'b0000000000000000;
	sram_mem[126508] = 16'b0000000000000000;
	sram_mem[126509] = 16'b0000000000000000;
	sram_mem[126510] = 16'b0000000000000000;
	sram_mem[126511] = 16'b0000000000000000;
	sram_mem[126512] = 16'b0000000000000000;
	sram_mem[126513] = 16'b0000000000000000;
	sram_mem[126514] = 16'b0000000000000000;
	sram_mem[126515] = 16'b0000000000000000;
	sram_mem[126516] = 16'b0000000000000000;
	sram_mem[126517] = 16'b0000000000000000;
	sram_mem[126518] = 16'b0000000000000000;
	sram_mem[126519] = 16'b0000000000000000;
	sram_mem[126520] = 16'b0000000000000000;
	sram_mem[126521] = 16'b0000000000000000;
	sram_mem[126522] = 16'b0000000000000000;
	sram_mem[126523] = 16'b0000000000000000;
	sram_mem[126524] = 16'b0000000000000000;
	sram_mem[126525] = 16'b0000000000000000;
	sram_mem[126526] = 16'b0000000000000000;
	sram_mem[126527] = 16'b0000000000000000;
	sram_mem[126528] = 16'b0000000000000000;
	sram_mem[126529] = 16'b0000000000000000;
	sram_mem[126530] = 16'b0000000000000000;
	sram_mem[126531] = 16'b0000000000000000;
	sram_mem[126532] = 16'b0000000000000000;
	sram_mem[126533] = 16'b0000000000000000;
	sram_mem[126534] = 16'b0000000000000000;
	sram_mem[126535] = 16'b0000000000000000;
	sram_mem[126536] = 16'b0000000000000000;
	sram_mem[126537] = 16'b0000000000000000;
	sram_mem[126538] = 16'b0000000000000000;
	sram_mem[126539] = 16'b0000000000000000;
	sram_mem[126540] = 16'b0000000000000000;
	sram_mem[126541] = 16'b0000000000000000;
	sram_mem[126542] = 16'b0000000000000000;
	sram_mem[126543] = 16'b0000000000000000;
	sram_mem[126544] = 16'b0000000000000000;
	sram_mem[126545] = 16'b0000000000000000;
	sram_mem[126546] = 16'b0000000000000000;
	sram_mem[126547] = 16'b0000000000000000;
	sram_mem[126548] = 16'b0000000000000000;
	sram_mem[126549] = 16'b0000000000000000;
	sram_mem[126550] = 16'b0000000000000000;
	sram_mem[126551] = 16'b0000000000000000;
	sram_mem[126552] = 16'b0000000000000000;
	sram_mem[126553] = 16'b0000000000000000;
	sram_mem[126554] = 16'b0000000000000000;
	sram_mem[126555] = 16'b0000000000000000;
	sram_mem[126556] = 16'b0000000000000000;
	sram_mem[126557] = 16'b0000000000000000;
	sram_mem[126558] = 16'b0000000000000000;
	sram_mem[126559] = 16'b0000000000000000;
	sram_mem[126560] = 16'b0000000000000000;
	sram_mem[126561] = 16'b0000000000000000;
	sram_mem[126562] = 16'b0000000000000000;
	sram_mem[126563] = 16'b0000000000000000;
	sram_mem[126564] = 16'b0000000000000000;
	sram_mem[126565] = 16'b0000000000000000;
	sram_mem[126566] = 16'b0000000000000000;
	sram_mem[126567] = 16'b0000000000000000;
	sram_mem[126568] = 16'b0000000000000000;
	sram_mem[126569] = 16'b0000000000000000;
	sram_mem[126570] = 16'b0000000000000000;
	sram_mem[126571] = 16'b0000000000000000;
	sram_mem[126572] = 16'b0000000000000000;
	sram_mem[126573] = 16'b0000000000000000;
	sram_mem[126574] = 16'b0000000000000000;
	sram_mem[126575] = 16'b0000000000000000;
	sram_mem[126576] = 16'b0000000000000000;
	sram_mem[126577] = 16'b0000000000000000;
	sram_mem[126578] = 16'b0000000000000000;
	sram_mem[126579] = 16'b0000000000000000;
	sram_mem[126580] = 16'b0000000000000000;
	sram_mem[126581] = 16'b0000000000000000;
	sram_mem[126582] = 16'b0000000000000000;
	sram_mem[126583] = 16'b0000000000000000;
	sram_mem[126584] = 16'b0000000000000000;
	sram_mem[126585] = 16'b0000000000000000;
	sram_mem[126586] = 16'b0000000000000000;
	sram_mem[126587] = 16'b0000000000000000;
	sram_mem[126588] = 16'b0000000000000000;
	sram_mem[126589] = 16'b0000000000000000;
	sram_mem[126590] = 16'b0000000000000000;
	sram_mem[126591] = 16'b0000000000000000;
	sram_mem[126592] = 16'b0000000000000000;
	sram_mem[126593] = 16'b0000000000000000;
	sram_mem[126594] = 16'b0000000000000000;
	sram_mem[126595] = 16'b0000000000000000;
	sram_mem[126596] = 16'b0000000000000000;
	sram_mem[126597] = 16'b0000000000000000;
	sram_mem[126598] = 16'b0000000000000000;
	sram_mem[126599] = 16'b0000000000000000;
	sram_mem[126600] = 16'b0000000000000000;
	sram_mem[126601] = 16'b0000000000000000;
	sram_mem[126602] = 16'b0000000000000000;
	sram_mem[126603] = 16'b0000000000000000;
	sram_mem[126604] = 16'b0000000000000000;
	sram_mem[126605] = 16'b0000000000000000;
	sram_mem[126606] = 16'b0000000000000000;
	sram_mem[126607] = 16'b0000000000000000;
	sram_mem[126608] = 16'b0000000000000000;
	sram_mem[126609] = 16'b0000000000000000;
	sram_mem[126610] = 16'b0000000000000000;
	sram_mem[126611] = 16'b0000000000000000;
	sram_mem[126612] = 16'b0000000000000000;
	sram_mem[126613] = 16'b0000000000000000;
	sram_mem[126614] = 16'b0000000000000000;
	sram_mem[126615] = 16'b0000000000000000;
	sram_mem[126616] = 16'b0000000000000000;
	sram_mem[126617] = 16'b0000000000000000;
	sram_mem[126618] = 16'b0000000000000000;
	sram_mem[126619] = 16'b0000000000000000;
	sram_mem[126620] = 16'b0000000000000000;
	sram_mem[126621] = 16'b0000000000000000;
	sram_mem[126622] = 16'b0000000000000000;
	sram_mem[126623] = 16'b0000000000000000;
	sram_mem[126624] = 16'b0000000000000000;
	sram_mem[126625] = 16'b0000000000000000;
	sram_mem[126626] = 16'b0000000000000000;
	sram_mem[126627] = 16'b0000000000000000;
	sram_mem[126628] = 16'b0000000000000000;
	sram_mem[126629] = 16'b0000000000000000;
	sram_mem[126630] = 16'b0000000000000000;
	sram_mem[126631] = 16'b0000000000000000;
	sram_mem[126632] = 16'b0000000000000000;
	sram_mem[126633] = 16'b0000000000000000;
	sram_mem[126634] = 16'b0000000000000000;
	sram_mem[126635] = 16'b0000000000000000;
	sram_mem[126636] = 16'b0000000000000000;
	sram_mem[126637] = 16'b0000000000000000;
	sram_mem[126638] = 16'b0000000000000000;
	sram_mem[126639] = 16'b0000000000000000;
	sram_mem[126640] = 16'b0000000000000000;
	sram_mem[126641] = 16'b0000000000000000;
	sram_mem[126642] = 16'b0000000000000000;
	sram_mem[126643] = 16'b0000000000000000;
	sram_mem[126644] = 16'b0000000000000000;
	sram_mem[126645] = 16'b0000000000000000;
	sram_mem[126646] = 16'b0000000000000000;
	sram_mem[126647] = 16'b0000000000000000;
	sram_mem[126648] = 16'b0000000000000000;
	sram_mem[126649] = 16'b0000000000000000;
	sram_mem[126650] = 16'b0000000000000000;
	sram_mem[126651] = 16'b0000000000000000;
	sram_mem[126652] = 16'b0000000000000000;
	sram_mem[126653] = 16'b0000000000000000;
	sram_mem[126654] = 16'b0000000000000000;
	sram_mem[126655] = 16'b0000000000000000;
	sram_mem[126656] = 16'b0000000000000000;
	sram_mem[126657] = 16'b0000000000000000;
	sram_mem[126658] = 16'b0000000000000000;
	sram_mem[126659] = 16'b0000000000000000;
	sram_mem[126660] = 16'b0000000000000000;
	sram_mem[126661] = 16'b0000000000000000;
	sram_mem[126662] = 16'b0000000000000000;
	sram_mem[126663] = 16'b0000000000000000;
	sram_mem[126664] = 16'b0000000000000000;
	sram_mem[126665] = 16'b0000000000000000;
	sram_mem[126666] = 16'b0000000000000000;
	sram_mem[126667] = 16'b0000000000000000;
	sram_mem[126668] = 16'b0000000000000000;
	sram_mem[126669] = 16'b0000000000000000;
	sram_mem[126670] = 16'b0000000000000000;
	sram_mem[126671] = 16'b0000000000000000;
	sram_mem[126672] = 16'b0000000000000000;
	sram_mem[126673] = 16'b0000000000000000;
	sram_mem[126674] = 16'b0000000000000000;
	sram_mem[126675] = 16'b0000000000000000;
	sram_mem[126676] = 16'b0000000000000000;
	sram_mem[126677] = 16'b0000000000000000;
	sram_mem[126678] = 16'b0000000000000000;
	sram_mem[126679] = 16'b0000000000000000;
	sram_mem[126680] = 16'b0000000000000000;
	sram_mem[126681] = 16'b0000000000000000;
	sram_mem[126682] = 16'b0000000000000000;
	sram_mem[126683] = 16'b0000000000000000;
	sram_mem[126684] = 16'b0000000000000000;
	sram_mem[126685] = 16'b0000000000000000;
	sram_mem[126686] = 16'b0000000000000000;
	sram_mem[126687] = 16'b0000000000000000;
	sram_mem[126688] = 16'b0000000000000000;
	sram_mem[126689] = 16'b0000000000000000;
	sram_mem[126690] = 16'b0000000000000000;
	sram_mem[126691] = 16'b0000000000000000;
	sram_mem[126692] = 16'b0000000000000000;
	sram_mem[126693] = 16'b0000000000000000;
	sram_mem[126694] = 16'b0000000000000000;
	sram_mem[126695] = 16'b0000000000000000;
	sram_mem[126696] = 16'b0000000000000000;
	sram_mem[126697] = 16'b0000000000000000;
	sram_mem[126698] = 16'b0000000000000000;
	sram_mem[126699] = 16'b0000000000000000;
	sram_mem[126700] = 16'b0000000000000000;
	sram_mem[126701] = 16'b0000000000000000;
	sram_mem[126702] = 16'b0000000000000000;
	sram_mem[126703] = 16'b0000000000000000;
	sram_mem[126704] = 16'b0000000000000000;
	sram_mem[126705] = 16'b0000000000000000;
	sram_mem[126706] = 16'b0000000000000000;
	sram_mem[126707] = 16'b0000000000000000;
	sram_mem[126708] = 16'b0000000000000000;
	sram_mem[126709] = 16'b0000000000000000;
	sram_mem[126710] = 16'b0000000000000000;
	sram_mem[126711] = 16'b0000000000000000;
	sram_mem[126712] = 16'b0000000000000000;
	sram_mem[126713] = 16'b0000000000000000;
	sram_mem[126714] = 16'b0000000000000000;
	sram_mem[126715] = 16'b0000000000000000;
	sram_mem[126716] = 16'b0000000000000000;
	sram_mem[126717] = 16'b0000000000000000;
	sram_mem[126718] = 16'b0000000000000000;
	sram_mem[126719] = 16'b0000000000000000;
	sram_mem[126720] = 16'b0000000000000000;
	sram_mem[126721] = 16'b0000000000000000;
	sram_mem[126722] = 16'b0000000000000000;
	sram_mem[126723] = 16'b0000000000000000;
	sram_mem[126724] = 16'b0000000000000000;
	sram_mem[126725] = 16'b0000000000000000;
	sram_mem[126726] = 16'b0000000000000000;
	sram_mem[126727] = 16'b0000000000000000;
	sram_mem[126728] = 16'b0000000000000000;
	sram_mem[126729] = 16'b0000000000000000;
	sram_mem[126730] = 16'b0000000000000000;
	sram_mem[126731] = 16'b0000000000000000;
	sram_mem[126732] = 16'b0000000000000000;
	sram_mem[126733] = 16'b0000000000000000;
	sram_mem[126734] = 16'b0000000000000000;
	sram_mem[126735] = 16'b0000000000000000;
	sram_mem[126736] = 16'b0000000000000000;
	sram_mem[126737] = 16'b0000000000000000;
	sram_mem[126738] = 16'b0000000000000000;
	sram_mem[126739] = 16'b0000000000000000;
	sram_mem[126740] = 16'b0000000000000000;
	sram_mem[126741] = 16'b0000000000000000;
	sram_mem[126742] = 16'b0000000000000000;
	sram_mem[126743] = 16'b0000000000000000;
	sram_mem[126744] = 16'b0000000000000000;
	sram_mem[126745] = 16'b0000000000000000;
	sram_mem[126746] = 16'b0000000000000000;
	sram_mem[126747] = 16'b0000000000000000;
	sram_mem[126748] = 16'b0000000000000000;
	sram_mem[126749] = 16'b0000000000000000;
	sram_mem[126750] = 16'b0000000000000000;
	sram_mem[126751] = 16'b0000000000000000;
	sram_mem[126752] = 16'b0000000000000000;
	sram_mem[126753] = 16'b0000000000000000;
	sram_mem[126754] = 16'b0000000000000000;
	sram_mem[126755] = 16'b0000000000000000;
	sram_mem[126756] = 16'b0000000000000000;
	sram_mem[126757] = 16'b0000000000000000;
	sram_mem[126758] = 16'b0000000000000000;
	sram_mem[126759] = 16'b0000000000000000;
	sram_mem[126760] = 16'b0000000000000000;
	sram_mem[126761] = 16'b0000000000000000;
	sram_mem[126762] = 16'b0000000000000000;
	sram_mem[126763] = 16'b0000000000000000;
	sram_mem[126764] = 16'b0000000000000000;
	sram_mem[126765] = 16'b0000000000000000;
	sram_mem[126766] = 16'b0000000000000000;
	sram_mem[126767] = 16'b0000000000000000;
	sram_mem[126768] = 16'b0000000000000000;
	sram_mem[126769] = 16'b0000000000000000;
	sram_mem[126770] = 16'b0000000000000000;
	sram_mem[126771] = 16'b0000000000000000;
	sram_mem[126772] = 16'b0000000000000000;
	sram_mem[126773] = 16'b0000000000000000;
	sram_mem[126774] = 16'b0000000000000000;
	sram_mem[126775] = 16'b0000000000000000;
	sram_mem[126776] = 16'b0000000000000000;
	sram_mem[126777] = 16'b0000000000000000;
	sram_mem[126778] = 16'b0000000000000000;
	sram_mem[126779] = 16'b0000000000000000;
	sram_mem[126780] = 16'b0000000000000000;
	sram_mem[126781] = 16'b0000000000000000;
	sram_mem[126782] = 16'b0000000000000000;
	sram_mem[126783] = 16'b0000000000000000;
	sram_mem[126784] = 16'b0000000000000000;
	sram_mem[126785] = 16'b0000000000000000;
	sram_mem[126786] = 16'b0000000000000000;
	sram_mem[126787] = 16'b0000000000000000;
	sram_mem[126788] = 16'b0000000000000000;
	sram_mem[126789] = 16'b0000000000000000;
	sram_mem[126790] = 16'b0000000000000000;
	sram_mem[126791] = 16'b0000000000000000;
	sram_mem[126792] = 16'b0000000000000000;
	sram_mem[126793] = 16'b0000000000000000;
	sram_mem[126794] = 16'b0000000000000000;
	sram_mem[126795] = 16'b0000000000000000;
	sram_mem[126796] = 16'b0000000000000000;
	sram_mem[126797] = 16'b0000000000000000;
	sram_mem[126798] = 16'b0000000000000000;
	sram_mem[126799] = 16'b0000000000000000;
	sram_mem[126800] = 16'b0000000000000000;
	sram_mem[126801] = 16'b0000000000000000;
	sram_mem[126802] = 16'b0000000000000000;
	sram_mem[126803] = 16'b0000000000000000;
	sram_mem[126804] = 16'b0000000000000000;
	sram_mem[126805] = 16'b0000000000000000;
	sram_mem[126806] = 16'b0000000000000000;
	sram_mem[126807] = 16'b0000000000000000;
	sram_mem[126808] = 16'b0000000000000000;
	sram_mem[126809] = 16'b0000000000000000;
	sram_mem[126810] = 16'b0000000000000000;
	sram_mem[126811] = 16'b0000000000000000;
	sram_mem[126812] = 16'b0000000000000000;
	sram_mem[126813] = 16'b0000000000000000;
	sram_mem[126814] = 16'b0000000000000000;
	sram_mem[126815] = 16'b0000000000000000;
	sram_mem[126816] = 16'b0000000000000000;
	sram_mem[126817] = 16'b0000000000000000;
	sram_mem[126818] = 16'b0000000000000000;
	sram_mem[126819] = 16'b0000000000000000;
	sram_mem[126820] = 16'b0000000000000000;
	sram_mem[126821] = 16'b0000000000000000;
	sram_mem[126822] = 16'b0000000000000000;
	sram_mem[126823] = 16'b0000000000000000;
	sram_mem[126824] = 16'b0000000000000000;
	sram_mem[126825] = 16'b0000000000000000;
	sram_mem[126826] = 16'b0000000000000000;
	sram_mem[126827] = 16'b0000000000000000;
	sram_mem[126828] = 16'b0000000000000000;
	sram_mem[126829] = 16'b0000000000000000;
	sram_mem[126830] = 16'b0000000000000000;
	sram_mem[126831] = 16'b0000000000000000;
	sram_mem[126832] = 16'b0000000000000000;
	sram_mem[126833] = 16'b0000000000000000;
	sram_mem[126834] = 16'b0000000000000000;
	sram_mem[126835] = 16'b0000000000000000;
	sram_mem[126836] = 16'b0000000000000000;
	sram_mem[126837] = 16'b0000000000000000;
	sram_mem[126838] = 16'b0000000000000000;
	sram_mem[126839] = 16'b0000000000000000;
	sram_mem[126840] = 16'b0000000000000000;
	sram_mem[126841] = 16'b0000000000000000;
	sram_mem[126842] = 16'b0000000000000000;
	sram_mem[126843] = 16'b0000000000000000;
	sram_mem[126844] = 16'b0000000000000000;
	sram_mem[126845] = 16'b0000000000000000;
	sram_mem[126846] = 16'b0000000000000000;
	sram_mem[126847] = 16'b0000000000000000;
	sram_mem[126848] = 16'b0000000000000000;
	sram_mem[126849] = 16'b0000000000000000;
	sram_mem[126850] = 16'b0000000000000000;
	sram_mem[126851] = 16'b0000000000000000;
	sram_mem[126852] = 16'b0000000000000000;
	sram_mem[126853] = 16'b0000000000000000;
	sram_mem[126854] = 16'b0000000000000000;
	sram_mem[126855] = 16'b0000000000000000;
	sram_mem[126856] = 16'b0000000000000000;
	sram_mem[126857] = 16'b0000000000000000;
	sram_mem[126858] = 16'b0000000000000000;
	sram_mem[126859] = 16'b0000000000000000;
	sram_mem[126860] = 16'b0000000000000000;
	sram_mem[126861] = 16'b0000000000000000;
	sram_mem[126862] = 16'b0000000000000000;
	sram_mem[126863] = 16'b0000000000000000;
	sram_mem[126864] = 16'b0000000000000000;
	sram_mem[126865] = 16'b0000000000000000;
	sram_mem[126866] = 16'b0000000000000000;
	sram_mem[126867] = 16'b0000000000000000;
	sram_mem[126868] = 16'b0000000000000000;
	sram_mem[126869] = 16'b0000000000000000;
	sram_mem[126870] = 16'b0000000000000000;
	sram_mem[126871] = 16'b0000000000000000;
	sram_mem[126872] = 16'b0000000000000000;
	sram_mem[126873] = 16'b0000000000000000;
	sram_mem[126874] = 16'b0000000000000000;
	sram_mem[126875] = 16'b0000000000000000;
	sram_mem[126876] = 16'b0000000000000000;
	sram_mem[126877] = 16'b0000000000000000;
	sram_mem[126878] = 16'b0000000000000000;
	sram_mem[126879] = 16'b0000000000000000;
	sram_mem[126880] = 16'b0000000000000000;
	sram_mem[126881] = 16'b0000000000000000;
	sram_mem[126882] = 16'b0000000000000000;
	sram_mem[126883] = 16'b0000000000000000;
	sram_mem[126884] = 16'b0000000000000000;
	sram_mem[126885] = 16'b0000000000000000;
	sram_mem[126886] = 16'b0000000000000000;
	sram_mem[126887] = 16'b0000000000000000;
	sram_mem[126888] = 16'b0000000000000000;
	sram_mem[126889] = 16'b0000000000000000;
	sram_mem[126890] = 16'b0000000000000000;
	sram_mem[126891] = 16'b0000000000000000;
	sram_mem[126892] = 16'b0000000000000000;
	sram_mem[126893] = 16'b0000000000000000;
	sram_mem[126894] = 16'b0000000000000000;
	sram_mem[126895] = 16'b0000000000000000;
	sram_mem[126896] = 16'b0000000000000000;
	sram_mem[126897] = 16'b0000000000000000;
	sram_mem[126898] = 16'b0000000000000000;
	sram_mem[126899] = 16'b0000000000000000;
	sram_mem[126900] = 16'b0000000000000000;
	sram_mem[126901] = 16'b0000000000000000;
	sram_mem[126902] = 16'b0000000000000000;
	sram_mem[126903] = 16'b0000000000000000;
	sram_mem[126904] = 16'b0000000000000000;
	sram_mem[126905] = 16'b0000000000000000;
	sram_mem[126906] = 16'b0000000000000000;
	sram_mem[126907] = 16'b0000000000000000;
	sram_mem[126908] = 16'b0000000000000000;
	sram_mem[126909] = 16'b0000000000000000;
	sram_mem[126910] = 16'b0000000000000000;
	sram_mem[126911] = 16'b0000000000000000;
	sram_mem[126912] = 16'b0000000000000000;
	sram_mem[126913] = 16'b0000000000000000;
	sram_mem[126914] = 16'b0000000000000000;
	sram_mem[126915] = 16'b0000000000000000;
	sram_mem[126916] = 16'b0000000000000000;
	sram_mem[126917] = 16'b0000000000000000;
	sram_mem[126918] = 16'b0000000000000000;
	sram_mem[126919] = 16'b0000000000000000;
	sram_mem[126920] = 16'b0000000000000000;
	sram_mem[126921] = 16'b0000000000000000;
	sram_mem[126922] = 16'b0000000000000000;
	sram_mem[126923] = 16'b0000000000000000;
	sram_mem[126924] = 16'b0000000000000000;
	sram_mem[126925] = 16'b0000000000000000;
	sram_mem[126926] = 16'b0000000000000000;
	sram_mem[126927] = 16'b0000000000000000;
	sram_mem[126928] = 16'b0000000000000000;
	sram_mem[126929] = 16'b0000000000000000;
	sram_mem[126930] = 16'b0000000000000000;
	sram_mem[126931] = 16'b0000000000000000;
	sram_mem[126932] = 16'b0000000000000000;
	sram_mem[126933] = 16'b0000000000000000;
	sram_mem[126934] = 16'b0000000000000000;
	sram_mem[126935] = 16'b0000000000000000;
	sram_mem[126936] = 16'b0000000000000000;
	sram_mem[126937] = 16'b0000000000000000;
	sram_mem[126938] = 16'b0000000000000000;
	sram_mem[126939] = 16'b0000000000000000;
	sram_mem[126940] = 16'b0000000000000000;
	sram_mem[126941] = 16'b0000000000000000;
	sram_mem[126942] = 16'b0000000000000000;
	sram_mem[126943] = 16'b0000000000000000;
	sram_mem[126944] = 16'b0000000000000000;
	sram_mem[126945] = 16'b0000000000000000;
	sram_mem[126946] = 16'b0000000000000000;
	sram_mem[126947] = 16'b0000000000000000;
	sram_mem[126948] = 16'b0000000000000000;
	sram_mem[126949] = 16'b0000000000000000;
	sram_mem[126950] = 16'b0000000000000000;
	sram_mem[126951] = 16'b0000000000000000;
	sram_mem[126952] = 16'b0000000000000000;
	sram_mem[126953] = 16'b0000000000000000;
	sram_mem[126954] = 16'b0000000000000000;
	sram_mem[126955] = 16'b0000000000000000;
	sram_mem[126956] = 16'b0000000000000000;
	sram_mem[126957] = 16'b0000000000000000;
	sram_mem[126958] = 16'b0000000000000000;
	sram_mem[126959] = 16'b0000000000000000;
	sram_mem[126960] = 16'b0000000000000000;
	sram_mem[126961] = 16'b0000000000000000;
	sram_mem[126962] = 16'b0000000000000000;
	sram_mem[126963] = 16'b0000000000000000;
	sram_mem[126964] = 16'b0000000000000000;
	sram_mem[126965] = 16'b0000000000000000;
	sram_mem[126966] = 16'b0000000000000000;
	sram_mem[126967] = 16'b0000000000000000;
	sram_mem[126968] = 16'b0000000000000000;
	sram_mem[126969] = 16'b0000000000000000;
	sram_mem[126970] = 16'b0000000000000000;
	sram_mem[126971] = 16'b0000000000000000;
	sram_mem[126972] = 16'b0000000000000000;
	sram_mem[126973] = 16'b0000000000000000;
	sram_mem[126974] = 16'b0000000000000000;
	sram_mem[126975] = 16'b0000000000000000;
	sram_mem[126976] = 16'b0000000000000000;
	sram_mem[126977] = 16'b0000000000000000;
	sram_mem[126978] = 16'b0000000000000000;
	sram_mem[126979] = 16'b0000000000000000;
	sram_mem[126980] = 16'b0000000000000000;
	sram_mem[126981] = 16'b0000000000000000;
	sram_mem[126982] = 16'b0000000000000000;
	sram_mem[126983] = 16'b0000000000000000;
	sram_mem[126984] = 16'b0000000000000000;
	sram_mem[126985] = 16'b0000000000000000;
	sram_mem[126986] = 16'b0000000000000000;
	sram_mem[126987] = 16'b0000000000000000;
	sram_mem[126988] = 16'b0000000000000000;
	sram_mem[126989] = 16'b0000000000000000;
	sram_mem[126990] = 16'b0000000000000000;
	sram_mem[126991] = 16'b0000000000000000;
	sram_mem[126992] = 16'b0000000000000000;
	sram_mem[126993] = 16'b0000000000000000;
	sram_mem[126994] = 16'b0000000000000000;
	sram_mem[126995] = 16'b0000000000000000;
	sram_mem[126996] = 16'b0000000000000000;
	sram_mem[126997] = 16'b0000000000000000;
	sram_mem[126998] = 16'b0000000000000000;
	sram_mem[126999] = 16'b0000000000000000;
	sram_mem[127000] = 16'b0000000000000000;
	sram_mem[127001] = 16'b0000000000000000;
	sram_mem[127002] = 16'b0000000000000000;
	sram_mem[127003] = 16'b0000000000000000;
	sram_mem[127004] = 16'b0000000000000000;
	sram_mem[127005] = 16'b0000000000000000;
	sram_mem[127006] = 16'b0000000000000000;
	sram_mem[127007] = 16'b0000000000000000;
	sram_mem[127008] = 16'b0000000000000000;
	sram_mem[127009] = 16'b0000000000000000;
	sram_mem[127010] = 16'b0000000000000000;
	sram_mem[127011] = 16'b0000000000000000;
	sram_mem[127012] = 16'b0000000000000000;
	sram_mem[127013] = 16'b0000000000000000;
	sram_mem[127014] = 16'b0000000000000000;
	sram_mem[127015] = 16'b0000000000000000;
	sram_mem[127016] = 16'b0000000000000000;
	sram_mem[127017] = 16'b0000000000000000;
	sram_mem[127018] = 16'b0000000000000000;
	sram_mem[127019] = 16'b0000000000000000;
	sram_mem[127020] = 16'b0000000000000000;
	sram_mem[127021] = 16'b0000000000000000;
	sram_mem[127022] = 16'b0000000000000000;
	sram_mem[127023] = 16'b0000000000000000;
	sram_mem[127024] = 16'b0000000000000000;
	sram_mem[127025] = 16'b0000000000000000;
	sram_mem[127026] = 16'b0000000000000000;
	sram_mem[127027] = 16'b0000000000000000;
	sram_mem[127028] = 16'b0000000000000000;
	sram_mem[127029] = 16'b0000000000000000;
	sram_mem[127030] = 16'b0000000000000000;
	sram_mem[127031] = 16'b0000000000000000;
	sram_mem[127032] = 16'b0000000000000000;
	sram_mem[127033] = 16'b0000000000000000;
	sram_mem[127034] = 16'b0000000000000000;
	sram_mem[127035] = 16'b0000000000000000;
	sram_mem[127036] = 16'b0000000000000000;
	sram_mem[127037] = 16'b0000000000000000;
	sram_mem[127038] = 16'b0000000000000000;
	sram_mem[127039] = 16'b0000000000000000;
	sram_mem[127040] = 16'b0000000000000000;
	sram_mem[127041] = 16'b0000000000000000;
	sram_mem[127042] = 16'b0000000000000000;
	sram_mem[127043] = 16'b0000000000000000;
	sram_mem[127044] = 16'b0000000000000000;
	sram_mem[127045] = 16'b0000000000000000;
	sram_mem[127046] = 16'b0000000000000000;
	sram_mem[127047] = 16'b0000000000000000;
	sram_mem[127048] = 16'b0000000000000000;
	sram_mem[127049] = 16'b0000000000000000;
	sram_mem[127050] = 16'b0000000000000000;
	sram_mem[127051] = 16'b0000000000000000;
	sram_mem[127052] = 16'b0000000000000000;
	sram_mem[127053] = 16'b0000000000000000;
	sram_mem[127054] = 16'b0000000000000000;
	sram_mem[127055] = 16'b0000000000000000;
	sram_mem[127056] = 16'b0000000000000000;
	sram_mem[127057] = 16'b0000000000000000;
	sram_mem[127058] = 16'b0000000000000000;
	sram_mem[127059] = 16'b0000000000000000;
	sram_mem[127060] = 16'b0000000000000000;
	sram_mem[127061] = 16'b0000000000000000;
	sram_mem[127062] = 16'b0000000000000000;
	sram_mem[127063] = 16'b0000000000000000;
	sram_mem[127064] = 16'b0000000000000000;
	sram_mem[127065] = 16'b0000000000000000;
	sram_mem[127066] = 16'b0000000000000000;
	sram_mem[127067] = 16'b0000000000000000;
	sram_mem[127068] = 16'b0000000000000000;
	sram_mem[127069] = 16'b0000000000000000;
	sram_mem[127070] = 16'b0000000000000000;
	sram_mem[127071] = 16'b0000000000000000;
	sram_mem[127072] = 16'b0000000000000000;
	sram_mem[127073] = 16'b0000000000000000;
	sram_mem[127074] = 16'b0000000000000000;
	sram_mem[127075] = 16'b0000000000000000;
	sram_mem[127076] = 16'b0000000000000000;
	sram_mem[127077] = 16'b0000000000000000;
	sram_mem[127078] = 16'b0000000000000000;
	sram_mem[127079] = 16'b0000000000000000;
	sram_mem[127080] = 16'b0000000000000000;
	sram_mem[127081] = 16'b0000000000000000;
	sram_mem[127082] = 16'b0000000000000000;
	sram_mem[127083] = 16'b0000000000000000;
	sram_mem[127084] = 16'b0000000000000000;
	sram_mem[127085] = 16'b0000000000000000;
	sram_mem[127086] = 16'b0000000000000000;
	sram_mem[127087] = 16'b0000000000000000;
	sram_mem[127088] = 16'b0000000000000000;
	sram_mem[127089] = 16'b0000000000000000;
	sram_mem[127090] = 16'b0000000000000000;
	sram_mem[127091] = 16'b0000000000000000;
	sram_mem[127092] = 16'b0000000000000000;
	sram_mem[127093] = 16'b0000000000000000;
	sram_mem[127094] = 16'b0000000000000000;
	sram_mem[127095] = 16'b0000000000000000;
	sram_mem[127096] = 16'b0000000000000000;
	sram_mem[127097] = 16'b0000000000000000;
	sram_mem[127098] = 16'b0000000000000000;
	sram_mem[127099] = 16'b0000000000000000;
	sram_mem[127100] = 16'b0000000000000000;
	sram_mem[127101] = 16'b0000000000000000;
	sram_mem[127102] = 16'b0000000000000000;
	sram_mem[127103] = 16'b0000000000000000;
	sram_mem[127104] = 16'b0000000000000000;
	sram_mem[127105] = 16'b0000000000000000;
	sram_mem[127106] = 16'b0000000000000000;
	sram_mem[127107] = 16'b0000000000000000;
	sram_mem[127108] = 16'b0000000000000000;
	sram_mem[127109] = 16'b0000000000000000;
	sram_mem[127110] = 16'b0000000000000000;
	sram_mem[127111] = 16'b0000000000000000;
	sram_mem[127112] = 16'b0000000000000000;
	sram_mem[127113] = 16'b0000000000000000;
	sram_mem[127114] = 16'b0000000000000000;
	sram_mem[127115] = 16'b0000000000000000;
	sram_mem[127116] = 16'b0000000000000000;
	sram_mem[127117] = 16'b0000000000000000;
	sram_mem[127118] = 16'b0000000000000000;
	sram_mem[127119] = 16'b0000000000000000;
	sram_mem[127120] = 16'b0000000000000000;
	sram_mem[127121] = 16'b0000000000000000;
	sram_mem[127122] = 16'b0000000000000000;
	sram_mem[127123] = 16'b0000000000000000;
	sram_mem[127124] = 16'b0000000000000000;
	sram_mem[127125] = 16'b0000000000000000;
	sram_mem[127126] = 16'b0000000000000000;
	sram_mem[127127] = 16'b0000000000000000;
	sram_mem[127128] = 16'b0000000000000000;
	sram_mem[127129] = 16'b0000000000000000;
	sram_mem[127130] = 16'b0000000000000000;
	sram_mem[127131] = 16'b0000000000000000;
	sram_mem[127132] = 16'b0000000000000000;
	sram_mem[127133] = 16'b0000000000000000;
	sram_mem[127134] = 16'b0000000000000000;
	sram_mem[127135] = 16'b0000000000000000;
	sram_mem[127136] = 16'b0000000000000000;
	sram_mem[127137] = 16'b0000000000000000;
	sram_mem[127138] = 16'b0000000000000000;
	sram_mem[127139] = 16'b0000000000000000;
	sram_mem[127140] = 16'b0000000000000000;
	sram_mem[127141] = 16'b0000000000000000;
	sram_mem[127142] = 16'b0000000000000000;
	sram_mem[127143] = 16'b0000000000000000;
	sram_mem[127144] = 16'b0000000000000000;
	sram_mem[127145] = 16'b0000000000000000;
	sram_mem[127146] = 16'b0000000000000000;
	sram_mem[127147] = 16'b0000000000000000;
	sram_mem[127148] = 16'b0000000000000000;
	sram_mem[127149] = 16'b0000000000000000;
	sram_mem[127150] = 16'b0000000000000000;
	sram_mem[127151] = 16'b0000000000000000;
	sram_mem[127152] = 16'b0000000000000000;
	sram_mem[127153] = 16'b0000000000000000;
	sram_mem[127154] = 16'b0000000000000000;
	sram_mem[127155] = 16'b0000000000000000;
	sram_mem[127156] = 16'b0000000000000000;
	sram_mem[127157] = 16'b0000000000000000;
	sram_mem[127158] = 16'b0000000000000000;
	sram_mem[127159] = 16'b0000000000000000;
	sram_mem[127160] = 16'b0000000000000000;
	sram_mem[127161] = 16'b0000000000000000;
	sram_mem[127162] = 16'b0000000000000000;
	sram_mem[127163] = 16'b0000000000000000;
	sram_mem[127164] = 16'b0000000000000000;
	sram_mem[127165] = 16'b0000000000000000;
	sram_mem[127166] = 16'b0000000000000000;
	sram_mem[127167] = 16'b0000000000000000;
	sram_mem[127168] = 16'b0000000000000000;
	sram_mem[127169] = 16'b0000000000000000;
	sram_mem[127170] = 16'b0000000000000000;
	sram_mem[127171] = 16'b0000000000000000;
	sram_mem[127172] = 16'b0000000000000000;
	sram_mem[127173] = 16'b0000000000000000;
	sram_mem[127174] = 16'b0000000000000000;
	sram_mem[127175] = 16'b0000000000000000;
	sram_mem[127176] = 16'b0000000000000000;
	sram_mem[127177] = 16'b0000000000000000;
	sram_mem[127178] = 16'b0000000000000000;
	sram_mem[127179] = 16'b0000000000000000;
	sram_mem[127180] = 16'b0000000000000000;
	sram_mem[127181] = 16'b0000000000000000;
	sram_mem[127182] = 16'b0000000000000000;
	sram_mem[127183] = 16'b0000000000000000;
	sram_mem[127184] = 16'b0000000000000000;
	sram_mem[127185] = 16'b0000000000000000;
	sram_mem[127186] = 16'b0000000000000000;
	sram_mem[127187] = 16'b0000000000000000;
	sram_mem[127188] = 16'b0000000000000000;
	sram_mem[127189] = 16'b0000000000000000;
	sram_mem[127190] = 16'b0000000000000000;
	sram_mem[127191] = 16'b0000000000000000;
	sram_mem[127192] = 16'b0000000000000000;
	sram_mem[127193] = 16'b0000000000000000;
	sram_mem[127194] = 16'b0000000000000000;
	sram_mem[127195] = 16'b0000000000000000;
	sram_mem[127196] = 16'b0000000000000000;
	sram_mem[127197] = 16'b0000000000000000;
	sram_mem[127198] = 16'b0000000000000000;
	sram_mem[127199] = 16'b0000000000000000;
	sram_mem[127200] = 16'b0000000000000000;
	sram_mem[127201] = 16'b0000000000000000;
	sram_mem[127202] = 16'b0000000000000000;
	sram_mem[127203] = 16'b0000000000000000;
	sram_mem[127204] = 16'b0000000000000000;
	sram_mem[127205] = 16'b0000000000000000;
	sram_mem[127206] = 16'b0000000000000000;
	sram_mem[127207] = 16'b0000000000000000;
	sram_mem[127208] = 16'b0000000000000000;
	sram_mem[127209] = 16'b0000000000000000;
	sram_mem[127210] = 16'b0000000000000000;
	sram_mem[127211] = 16'b0000000000000000;
	sram_mem[127212] = 16'b0000000000000000;
	sram_mem[127213] = 16'b0000000000000000;
	sram_mem[127214] = 16'b0000000000000000;
	sram_mem[127215] = 16'b0000000000000000;
	sram_mem[127216] = 16'b0000000000000000;
	sram_mem[127217] = 16'b0000000000000000;
	sram_mem[127218] = 16'b0000000000000000;
	sram_mem[127219] = 16'b0000000000000000;
	sram_mem[127220] = 16'b0000000000000000;
	sram_mem[127221] = 16'b0000000000000000;
	sram_mem[127222] = 16'b0000000000000000;
	sram_mem[127223] = 16'b0000000000000000;
	sram_mem[127224] = 16'b0000000000000000;
	sram_mem[127225] = 16'b0000000000000000;
	sram_mem[127226] = 16'b0000000000000000;
	sram_mem[127227] = 16'b0000000000000000;
	sram_mem[127228] = 16'b0000000000000000;
	sram_mem[127229] = 16'b0000000000000000;
	sram_mem[127230] = 16'b0000000000000000;
	sram_mem[127231] = 16'b0000000000000000;
	sram_mem[127232] = 16'b0000000000000000;
	sram_mem[127233] = 16'b0000000000000000;
	sram_mem[127234] = 16'b0000000000000000;
	sram_mem[127235] = 16'b0000000000000000;
	sram_mem[127236] = 16'b0000000000000000;
	sram_mem[127237] = 16'b0000000000000000;
	sram_mem[127238] = 16'b0000000000000000;
	sram_mem[127239] = 16'b0000000000000000;
	sram_mem[127240] = 16'b0000000000000000;
	sram_mem[127241] = 16'b0000000000000000;
	sram_mem[127242] = 16'b0000000000000000;
	sram_mem[127243] = 16'b0000000000000000;
	sram_mem[127244] = 16'b0000000000000000;
	sram_mem[127245] = 16'b0000000000000000;
	sram_mem[127246] = 16'b0000000000000000;
	sram_mem[127247] = 16'b0000000000000000;
	sram_mem[127248] = 16'b0000000000000000;
	sram_mem[127249] = 16'b0000000000000000;
	sram_mem[127250] = 16'b0000000000000000;
	sram_mem[127251] = 16'b0000000000000000;
	sram_mem[127252] = 16'b0000000000000000;
	sram_mem[127253] = 16'b0000000000000000;
	sram_mem[127254] = 16'b0000000000000000;
	sram_mem[127255] = 16'b0000000000000000;
	sram_mem[127256] = 16'b0000000000000000;
	sram_mem[127257] = 16'b0000000000000000;
	sram_mem[127258] = 16'b0000000000000000;
	sram_mem[127259] = 16'b0000000000000000;
	sram_mem[127260] = 16'b0000000000000000;
	sram_mem[127261] = 16'b0000000000000000;
	sram_mem[127262] = 16'b0000000000000000;
	sram_mem[127263] = 16'b0000000000000000;
	sram_mem[127264] = 16'b0000000000000000;
	sram_mem[127265] = 16'b0000000000000000;
	sram_mem[127266] = 16'b0000000000000000;
	sram_mem[127267] = 16'b0000000000000000;
	sram_mem[127268] = 16'b0000000000000000;
	sram_mem[127269] = 16'b0000000000000000;
	sram_mem[127270] = 16'b0000000000000000;
	sram_mem[127271] = 16'b0000000000000000;
	sram_mem[127272] = 16'b0000000000000000;
	sram_mem[127273] = 16'b0000000000000000;
	sram_mem[127274] = 16'b0000000000000000;
	sram_mem[127275] = 16'b0000000000000000;
	sram_mem[127276] = 16'b0000000000000000;
	sram_mem[127277] = 16'b0000000000000000;
	sram_mem[127278] = 16'b0000000000000000;
	sram_mem[127279] = 16'b0000000000000000;
	sram_mem[127280] = 16'b0000000000000000;
	sram_mem[127281] = 16'b0000000000000000;
	sram_mem[127282] = 16'b0000000000000000;
	sram_mem[127283] = 16'b0000000000000000;
	sram_mem[127284] = 16'b0000000000000000;
	sram_mem[127285] = 16'b0000000000000000;
	sram_mem[127286] = 16'b0000000000000000;
	sram_mem[127287] = 16'b0000000000000000;
	sram_mem[127288] = 16'b0000000000000000;
	sram_mem[127289] = 16'b0000000000000000;
	sram_mem[127290] = 16'b0000000000000000;
	sram_mem[127291] = 16'b0000000000000000;
	sram_mem[127292] = 16'b0000000000000000;
	sram_mem[127293] = 16'b0000000000000000;
	sram_mem[127294] = 16'b0000000000000000;
	sram_mem[127295] = 16'b0000000000000000;
	sram_mem[127296] = 16'b0000000000000000;
	sram_mem[127297] = 16'b0000000000000000;
	sram_mem[127298] = 16'b0000000000000000;
	sram_mem[127299] = 16'b0000000000000000;
	sram_mem[127300] = 16'b0000000000000000;
	sram_mem[127301] = 16'b0000000000000000;
	sram_mem[127302] = 16'b0000000000000000;
	sram_mem[127303] = 16'b0000000000000000;
	sram_mem[127304] = 16'b0000000000000000;
	sram_mem[127305] = 16'b0000000000000000;
	sram_mem[127306] = 16'b0000000000000000;
	sram_mem[127307] = 16'b0000000000000000;
	sram_mem[127308] = 16'b0000000000000000;
	sram_mem[127309] = 16'b0000000000000000;
	sram_mem[127310] = 16'b0000000000000000;
	sram_mem[127311] = 16'b0000000000000000;
	sram_mem[127312] = 16'b0000000000000000;
	sram_mem[127313] = 16'b0000000000000000;
	sram_mem[127314] = 16'b0000000000000000;
	sram_mem[127315] = 16'b0000000000000000;
	sram_mem[127316] = 16'b0000000000000000;
	sram_mem[127317] = 16'b0000000000000000;
	sram_mem[127318] = 16'b0000000000000000;
	sram_mem[127319] = 16'b0000000000000000;
	sram_mem[127320] = 16'b0000000000000000;
	sram_mem[127321] = 16'b0000000000000000;
	sram_mem[127322] = 16'b0000000000000000;
	sram_mem[127323] = 16'b0000000000000000;
	sram_mem[127324] = 16'b0000000000000000;
	sram_mem[127325] = 16'b0000000000000000;
	sram_mem[127326] = 16'b0000000000000000;
	sram_mem[127327] = 16'b0000000000000000;
	sram_mem[127328] = 16'b0000000000000000;
	sram_mem[127329] = 16'b0000000000000000;
	sram_mem[127330] = 16'b0000000000000000;
	sram_mem[127331] = 16'b0000000000000000;
	sram_mem[127332] = 16'b0000000000000000;
	sram_mem[127333] = 16'b0000000000000000;
	sram_mem[127334] = 16'b0000000000000000;
	sram_mem[127335] = 16'b0000000000000000;
	sram_mem[127336] = 16'b0000000000000000;
	sram_mem[127337] = 16'b0000000000000000;
	sram_mem[127338] = 16'b0000000000000000;
	sram_mem[127339] = 16'b0000000000000000;
	sram_mem[127340] = 16'b0000000000000000;
	sram_mem[127341] = 16'b0000000000000000;
	sram_mem[127342] = 16'b0000000000000000;
	sram_mem[127343] = 16'b0000000000000000;
	sram_mem[127344] = 16'b0000000000000000;
	sram_mem[127345] = 16'b0000000000000000;
	sram_mem[127346] = 16'b0000000000000000;
	sram_mem[127347] = 16'b0000000000000000;
	sram_mem[127348] = 16'b0000000000000000;
	sram_mem[127349] = 16'b0000000000000000;
	sram_mem[127350] = 16'b0000000000000000;
	sram_mem[127351] = 16'b0000000000000000;
	sram_mem[127352] = 16'b0000000000000000;
	sram_mem[127353] = 16'b0000000000000000;
	sram_mem[127354] = 16'b0000000000000000;
	sram_mem[127355] = 16'b0000000000000000;
	sram_mem[127356] = 16'b0000000000000000;
	sram_mem[127357] = 16'b0000000000000000;
	sram_mem[127358] = 16'b0000000000000000;
	sram_mem[127359] = 16'b0000000000000000;
	sram_mem[127360] = 16'b0000000000000000;
	sram_mem[127361] = 16'b0000000000000000;
	sram_mem[127362] = 16'b0000000000000000;
	sram_mem[127363] = 16'b0000000000000000;
	sram_mem[127364] = 16'b0000000000000000;
	sram_mem[127365] = 16'b0000000000000000;
	sram_mem[127366] = 16'b0000000000000000;
	sram_mem[127367] = 16'b0000000000000000;
	sram_mem[127368] = 16'b0000000000000000;
	sram_mem[127369] = 16'b0000000000000000;
	sram_mem[127370] = 16'b0000000000000000;
	sram_mem[127371] = 16'b0000000000000000;
	sram_mem[127372] = 16'b0000000000000000;
	sram_mem[127373] = 16'b0000000000000000;
	sram_mem[127374] = 16'b0000000000000000;
	sram_mem[127375] = 16'b0000000000000000;
	sram_mem[127376] = 16'b0000000000000000;
	sram_mem[127377] = 16'b0000000000000000;
	sram_mem[127378] = 16'b0000000000000000;
	sram_mem[127379] = 16'b0000000000000000;
	sram_mem[127380] = 16'b0000000000000000;
	sram_mem[127381] = 16'b0000000000000000;
	sram_mem[127382] = 16'b0000000000000000;
	sram_mem[127383] = 16'b0000000000000000;
	sram_mem[127384] = 16'b0000000000000000;
	sram_mem[127385] = 16'b0000000000000000;
	sram_mem[127386] = 16'b0000000000000000;
	sram_mem[127387] = 16'b0000000000000000;
	sram_mem[127388] = 16'b0000000000000000;
	sram_mem[127389] = 16'b0000000000000000;
	sram_mem[127390] = 16'b0000000000000000;
	sram_mem[127391] = 16'b0000000000000000;
	sram_mem[127392] = 16'b0000000000000000;
	sram_mem[127393] = 16'b0000000000000000;
	sram_mem[127394] = 16'b0000000000000000;
	sram_mem[127395] = 16'b0000000000000000;
	sram_mem[127396] = 16'b0000000000000000;
	sram_mem[127397] = 16'b0000000000000000;
	sram_mem[127398] = 16'b0000000000000000;
	sram_mem[127399] = 16'b0000000000000000;
	sram_mem[127400] = 16'b0000000000000000;
	sram_mem[127401] = 16'b0000000000000000;
	sram_mem[127402] = 16'b0000000000000000;
	sram_mem[127403] = 16'b0000000000000000;
	sram_mem[127404] = 16'b0000000000000000;
	sram_mem[127405] = 16'b0000000000000000;
	sram_mem[127406] = 16'b0000000000000000;
	sram_mem[127407] = 16'b0000000000000000;
	sram_mem[127408] = 16'b0000000000000000;
	sram_mem[127409] = 16'b0000000000000000;
	sram_mem[127410] = 16'b0000000000000000;
	sram_mem[127411] = 16'b0000000000000000;
	sram_mem[127412] = 16'b0000000000000000;
	sram_mem[127413] = 16'b0000000000000000;
	sram_mem[127414] = 16'b0000000000000000;
	sram_mem[127415] = 16'b0000000000000000;
	sram_mem[127416] = 16'b0000000000000000;
	sram_mem[127417] = 16'b0000000000000000;
	sram_mem[127418] = 16'b0000000000000000;
	sram_mem[127419] = 16'b0000000000000000;
	sram_mem[127420] = 16'b0000000000000000;
	sram_mem[127421] = 16'b0000000000000000;
	sram_mem[127422] = 16'b0000000000000000;
	sram_mem[127423] = 16'b0000000000000000;
	sram_mem[127424] = 16'b0000000000000000;
	sram_mem[127425] = 16'b0000000000000000;
	sram_mem[127426] = 16'b0000000000000000;
	sram_mem[127427] = 16'b0000000000000000;
	sram_mem[127428] = 16'b0000000000000000;
	sram_mem[127429] = 16'b0000000000000000;
	sram_mem[127430] = 16'b0000000000000000;
	sram_mem[127431] = 16'b0000000000000000;
	sram_mem[127432] = 16'b0000000000000000;
	sram_mem[127433] = 16'b0000000000000000;
	sram_mem[127434] = 16'b0000000000000000;
	sram_mem[127435] = 16'b0000000000000000;
	sram_mem[127436] = 16'b0000000000000000;
	sram_mem[127437] = 16'b0000000000000000;
	sram_mem[127438] = 16'b0000000000000000;
	sram_mem[127439] = 16'b0000000000000000;
	sram_mem[127440] = 16'b0000000000000000;
	sram_mem[127441] = 16'b0000000000000000;
	sram_mem[127442] = 16'b0000000000000000;
	sram_mem[127443] = 16'b0000000000000000;
	sram_mem[127444] = 16'b0000000000000000;
	sram_mem[127445] = 16'b0000000000000000;
	sram_mem[127446] = 16'b0000000000000000;
	sram_mem[127447] = 16'b0000000000000000;
	sram_mem[127448] = 16'b0000000000000000;
	sram_mem[127449] = 16'b0000000000000000;
	sram_mem[127450] = 16'b0000000000000000;
	sram_mem[127451] = 16'b0000000000000000;
	sram_mem[127452] = 16'b0000000000000000;
	sram_mem[127453] = 16'b0000000000000000;
	sram_mem[127454] = 16'b0000000000000000;
	sram_mem[127455] = 16'b0000000000000000;
	sram_mem[127456] = 16'b0000000000000000;
	sram_mem[127457] = 16'b0000000000000000;
	sram_mem[127458] = 16'b0000000000000000;
	sram_mem[127459] = 16'b0000000000000000;
	sram_mem[127460] = 16'b0000000000000000;
	sram_mem[127461] = 16'b0000000000000000;
	sram_mem[127462] = 16'b0000000000000000;
	sram_mem[127463] = 16'b0000000000000000;
	sram_mem[127464] = 16'b0000000000000000;
	sram_mem[127465] = 16'b0000000000000000;
	sram_mem[127466] = 16'b0000000000000000;
	sram_mem[127467] = 16'b0000000000000000;
	sram_mem[127468] = 16'b0000000000000000;
	sram_mem[127469] = 16'b0000000000000000;
	sram_mem[127470] = 16'b0000000000000000;
	sram_mem[127471] = 16'b0000000000000000;
	sram_mem[127472] = 16'b0000000000000000;
	sram_mem[127473] = 16'b0000000000000000;
	sram_mem[127474] = 16'b0000000000000000;
	sram_mem[127475] = 16'b0000000000000000;
	sram_mem[127476] = 16'b0000000000000000;
	sram_mem[127477] = 16'b0000000000000000;
	sram_mem[127478] = 16'b0000000000000000;
	sram_mem[127479] = 16'b0000000000000000;
	sram_mem[127480] = 16'b0000000000000000;
	sram_mem[127481] = 16'b0000000000000000;
	sram_mem[127482] = 16'b0000000000000000;
	sram_mem[127483] = 16'b0000000000000000;
	sram_mem[127484] = 16'b0000000000000000;
	sram_mem[127485] = 16'b0000000000000000;
	sram_mem[127486] = 16'b0000000000000000;
	sram_mem[127487] = 16'b0000000000000000;
	sram_mem[127488] = 16'b0000000000000000;
	sram_mem[127489] = 16'b0000000000000000;
	sram_mem[127490] = 16'b0000000000000000;
	sram_mem[127491] = 16'b0000000000000000;
	sram_mem[127492] = 16'b0000000000000000;
	sram_mem[127493] = 16'b0000000000000000;
	sram_mem[127494] = 16'b0000000000000000;
	sram_mem[127495] = 16'b0000000000000000;
	sram_mem[127496] = 16'b0000000000000000;
	sram_mem[127497] = 16'b0000000000000000;
	sram_mem[127498] = 16'b0000000000000000;
	sram_mem[127499] = 16'b0000000000000000;
	sram_mem[127500] = 16'b0000000000000000;
	sram_mem[127501] = 16'b0000000000000000;
	sram_mem[127502] = 16'b0000000000000000;
	sram_mem[127503] = 16'b0000000000000000;
	sram_mem[127504] = 16'b0000000000000000;
	sram_mem[127505] = 16'b0000000000000000;
	sram_mem[127506] = 16'b0000000000000000;
	sram_mem[127507] = 16'b0000000000000000;
	sram_mem[127508] = 16'b0000000000000000;
	sram_mem[127509] = 16'b0000000000000000;
	sram_mem[127510] = 16'b0000000000000000;
	sram_mem[127511] = 16'b0000000000000000;
	sram_mem[127512] = 16'b0000000000000000;
	sram_mem[127513] = 16'b0000000000000000;
	sram_mem[127514] = 16'b0000000000000000;
	sram_mem[127515] = 16'b0000000000000000;
	sram_mem[127516] = 16'b0000000000000000;
	sram_mem[127517] = 16'b0000000000000000;
	sram_mem[127518] = 16'b0000000000000000;
	sram_mem[127519] = 16'b0000000000000000;
	sram_mem[127520] = 16'b0000000000000000;
	sram_mem[127521] = 16'b0000000000000000;
	sram_mem[127522] = 16'b0000000000000000;
	sram_mem[127523] = 16'b0000000000000000;
	sram_mem[127524] = 16'b0000000000000000;
	sram_mem[127525] = 16'b0000000000000000;
	sram_mem[127526] = 16'b0000000000000000;
	sram_mem[127527] = 16'b0000000000000000;
	sram_mem[127528] = 16'b0000000000000000;
	sram_mem[127529] = 16'b0000000000000000;
	sram_mem[127530] = 16'b0000000000000000;
	sram_mem[127531] = 16'b0000000000000000;
	sram_mem[127532] = 16'b0000000000000000;
	sram_mem[127533] = 16'b0000000000000000;
	sram_mem[127534] = 16'b0000000000000000;
	sram_mem[127535] = 16'b0000000000000000;
	sram_mem[127536] = 16'b0000000000000000;
	sram_mem[127537] = 16'b0000000000000000;
	sram_mem[127538] = 16'b0000000000000000;
	sram_mem[127539] = 16'b0000000000000000;
	sram_mem[127540] = 16'b0000000000000000;
	sram_mem[127541] = 16'b0000000000000000;
	sram_mem[127542] = 16'b0000000000000000;
	sram_mem[127543] = 16'b0000000000000000;
	sram_mem[127544] = 16'b0000000000000000;
	sram_mem[127545] = 16'b0000000000000000;
	sram_mem[127546] = 16'b0000000000000000;
	sram_mem[127547] = 16'b0000000000000000;
	sram_mem[127548] = 16'b0000000000000000;
	sram_mem[127549] = 16'b0000000000000000;
	sram_mem[127550] = 16'b0000000000000000;
	sram_mem[127551] = 16'b0000000000000000;
	sram_mem[127552] = 16'b0000000000000000;
	sram_mem[127553] = 16'b0000000000000000;
	sram_mem[127554] = 16'b0000000000000000;
	sram_mem[127555] = 16'b0000000000000000;
	sram_mem[127556] = 16'b0000000000000000;
	sram_mem[127557] = 16'b0000000000000000;
	sram_mem[127558] = 16'b0000000000000000;
	sram_mem[127559] = 16'b0000000000000000;
	sram_mem[127560] = 16'b0000000000000000;
	sram_mem[127561] = 16'b0000000000000000;
	sram_mem[127562] = 16'b0000000000000000;
	sram_mem[127563] = 16'b0000000000000000;
	sram_mem[127564] = 16'b0000000000000000;
	sram_mem[127565] = 16'b0000000000000000;
	sram_mem[127566] = 16'b0000000000000000;
	sram_mem[127567] = 16'b0000000000000000;
	sram_mem[127568] = 16'b0000000000000000;
	sram_mem[127569] = 16'b0000000000000000;
	sram_mem[127570] = 16'b0000000000000000;
	sram_mem[127571] = 16'b0000000000000000;
	sram_mem[127572] = 16'b0000000000000000;
	sram_mem[127573] = 16'b0000000000000000;
	sram_mem[127574] = 16'b0000000000000000;
	sram_mem[127575] = 16'b0000000000000000;
	sram_mem[127576] = 16'b0000000000000000;
	sram_mem[127577] = 16'b0000000000000000;
	sram_mem[127578] = 16'b0000000000000000;
	sram_mem[127579] = 16'b0000000000000000;
	sram_mem[127580] = 16'b0000000000000000;
	sram_mem[127581] = 16'b0000000000000000;
	sram_mem[127582] = 16'b0000000000000000;
	sram_mem[127583] = 16'b0000000000000000;
	sram_mem[127584] = 16'b0000000000000000;
	sram_mem[127585] = 16'b0000000000000000;
	sram_mem[127586] = 16'b0000000000000000;
	sram_mem[127587] = 16'b0000000000000000;
	sram_mem[127588] = 16'b0000000000000000;
	sram_mem[127589] = 16'b0000000000000000;
	sram_mem[127590] = 16'b0000000000000000;
	sram_mem[127591] = 16'b0000000000000000;
	sram_mem[127592] = 16'b0000000000000000;
	sram_mem[127593] = 16'b0000000000000000;
	sram_mem[127594] = 16'b0000000000000000;
	sram_mem[127595] = 16'b0000000000000000;
	sram_mem[127596] = 16'b0000000000000000;
	sram_mem[127597] = 16'b0000000000000000;
	sram_mem[127598] = 16'b0000000000000000;
	sram_mem[127599] = 16'b0000000000000000;
	sram_mem[127600] = 16'b0000000000000000;
	sram_mem[127601] = 16'b0000000000000000;
	sram_mem[127602] = 16'b0000000000000000;
	sram_mem[127603] = 16'b0000000000000000;
	sram_mem[127604] = 16'b0000000000000000;
	sram_mem[127605] = 16'b0000000000000000;
	sram_mem[127606] = 16'b0000000000000000;
	sram_mem[127607] = 16'b0000000000000000;
	sram_mem[127608] = 16'b0000000000000000;
	sram_mem[127609] = 16'b0000000000000000;
	sram_mem[127610] = 16'b0000000000000000;
	sram_mem[127611] = 16'b0000000000000000;
	sram_mem[127612] = 16'b0000000000000000;
	sram_mem[127613] = 16'b0000000000000000;
	sram_mem[127614] = 16'b0000000000000000;
	sram_mem[127615] = 16'b0000000000000000;
	sram_mem[127616] = 16'b0000000000000000;
	sram_mem[127617] = 16'b0000000000000000;
	sram_mem[127618] = 16'b0000000000000000;
	sram_mem[127619] = 16'b0000000000000000;
	sram_mem[127620] = 16'b0000000000000000;
	sram_mem[127621] = 16'b0000000000000000;
	sram_mem[127622] = 16'b0000000000000000;
	sram_mem[127623] = 16'b0000000000000000;
	sram_mem[127624] = 16'b0000000000000000;
	sram_mem[127625] = 16'b0000000000000000;
	sram_mem[127626] = 16'b0000000000000000;
	sram_mem[127627] = 16'b0000000000000000;
	sram_mem[127628] = 16'b0000000000000000;
	sram_mem[127629] = 16'b0000000000000000;
	sram_mem[127630] = 16'b0000000000000000;
	sram_mem[127631] = 16'b0000000000000000;
	sram_mem[127632] = 16'b0000000000000000;
	sram_mem[127633] = 16'b0000000000000000;
	sram_mem[127634] = 16'b0000000000000000;
	sram_mem[127635] = 16'b0000000000000000;
	sram_mem[127636] = 16'b0000000000000000;
	sram_mem[127637] = 16'b0000000000000000;
	sram_mem[127638] = 16'b0000000000000000;
	sram_mem[127639] = 16'b0000000000000000;
	sram_mem[127640] = 16'b0000000000000000;
	sram_mem[127641] = 16'b0000000000000000;
	sram_mem[127642] = 16'b0000000000000000;
	sram_mem[127643] = 16'b0000000000000000;
	sram_mem[127644] = 16'b0000000000000000;
	sram_mem[127645] = 16'b0000000000000000;
	sram_mem[127646] = 16'b0000000000000000;
	sram_mem[127647] = 16'b0000000000000000;
	sram_mem[127648] = 16'b0000000000000000;
	sram_mem[127649] = 16'b0000000000000000;
	sram_mem[127650] = 16'b0000000000000000;
	sram_mem[127651] = 16'b0000000000000000;
	sram_mem[127652] = 16'b0000000000000000;
	sram_mem[127653] = 16'b0000000000000000;
	sram_mem[127654] = 16'b0000000000000000;
	sram_mem[127655] = 16'b0000000000000000;
	sram_mem[127656] = 16'b0000000000000000;
	sram_mem[127657] = 16'b0000000000000000;
	sram_mem[127658] = 16'b0000000000000000;
	sram_mem[127659] = 16'b0000000000000000;
	sram_mem[127660] = 16'b0000000000000000;
	sram_mem[127661] = 16'b0000000000000000;
	sram_mem[127662] = 16'b0000000000000000;
	sram_mem[127663] = 16'b0000000000000000;
	sram_mem[127664] = 16'b0000000000000000;
	sram_mem[127665] = 16'b0000000000000000;
	sram_mem[127666] = 16'b0000000000000000;
	sram_mem[127667] = 16'b0000000000000000;
	sram_mem[127668] = 16'b0000000000000000;
	sram_mem[127669] = 16'b0000000000000000;
	sram_mem[127670] = 16'b0000000000000000;
	sram_mem[127671] = 16'b0000000000000000;
	sram_mem[127672] = 16'b0000000000000000;
	sram_mem[127673] = 16'b0000000000000000;
	sram_mem[127674] = 16'b0000000000000000;
	sram_mem[127675] = 16'b0000000000000000;
	sram_mem[127676] = 16'b0000000000000000;
	sram_mem[127677] = 16'b0000000000000000;
	sram_mem[127678] = 16'b0000000000000000;
	sram_mem[127679] = 16'b0000000000000000;
	sram_mem[127680] = 16'b0000000000000000;
	sram_mem[127681] = 16'b0000000000000000;
	sram_mem[127682] = 16'b0000000000000000;
	sram_mem[127683] = 16'b0000000000000000;
	sram_mem[127684] = 16'b0000000000000000;
	sram_mem[127685] = 16'b0000000000000000;
	sram_mem[127686] = 16'b0000000000000000;
	sram_mem[127687] = 16'b0000000000000000;
	sram_mem[127688] = 16'b0000000000000000;
	sram_mem[127689] = 16'b0000000000000000;
	sram_mem[127690] = 16'b0000000000000000;
	sram_mem[127691] = 16'b0000000000000000;
	sram_mem[127692] = 16'b0000000000000000;
	sram_mem[127693] = 16'b0000000000000000;
	sram_mem[127694] = 16'b0000000000000000;
	sram_mem[127695] = 16'b0000000000000000;
	sram_mem[127696] = 16'b0000000000000000;
	sram_mem[127697] = 16'b0000000000000000;
	sram_mem[127698] = 16'b0000000000000000;
	sram_mem[127699] = 16'b0000000000000000;
	sram_mem[127700] = 16'b0000000000000000;
	sram_mem[127701] = 16'b0000000000000000;
	sram_mem[127702] = 16'b0000000000000000;
	sram_mem[127703] = 16'b0000000000000000;
	sram_mem[127704] = 16'b0000000000000000;
	sram_mem[127705] = 16'b0000000000000000;
	sram_mem[127706] = 16'b0000000000000000;
	sram_mem[127707] = 16'b0000000000000000;
	sram_mem[127708] = 16'b0000000000000000;
	sram_mem[127709] = 16'b0000000000000000;
	sram_mem[127710] = 16'b0000000000000000;
	sram_mem[127711] = 16'b0000000000000000;
	sram_mem[127712] = 16'b0000000000000000;
	sram_mem[127713] = 16'b0000000000000000;
	sram_mem[127714] = 16'b0000000000000000;
	sram_mem[127715] = 16'b0000000000000000;
	sram_mem[127716] = 16'b0000000000000000;
	sram_mem[127717] = 16'b0000000000000000;
	sram_mem[127718] = 16'b0000000000000000;
	sram_mem[127719] = 16'b0000000000000000;
	sram_mem[127720] = 16'b0000000000000000;
	sram_mem[127721] = 16'b0000000000000000;
	sram_mem[127722] = 16'b0000000000000000;
	sram_mem[127723] = 16'b0000000000000000;
	sram_mem[127724] = 16'b0000000000000000;
	sram_mem[127725] = 16'b0000000000000000;
	sram_mem[127726] = 16'b0000000000000000;
	sram_mem[127727] = 16'b0000000000000000;
	sram_mem[127728] = 16'b0000000000000000;
	sram_mem[127729] = 16'b0000000000000000;
	sram_mem[127730] = 16'b0000000000000000;
	sram_mem[127731] = 16'b0000000000000000;
	sram_mem[127732] = 16'b0000000000000000;
	sram_mem[127733] = 16'b0000000000000000;
	sram_mem[127734] = 16'b0000000000000000;
	sram_mem[127735] = 16'b0000000000000000;
	sram_mem[127736] = 16'b0000000000000000;
	sram_mem[127737] = 16'b0000000000000000;
	sram_mem[127738] = 16'b0000000000000000;
	sram_mem[127739] = 16'b0000000000000000;
	sram_mem[127740] = 16'b0000000000000000;
	sram_mem[127741] = 16'b0000000000000000;
	sram_mem[127742] = 16'b0000000000000000;
	sram_mem[127743] = 16'b0000000000000000;
	sram_mem[127744] = 16'b0000000000000000;
	sram_mem[127745] = 16'b0000000000000000;
	sram_mem[127746] = 16'b0000000000000000;
	sram_mem[127747] = 16'b0000000000000000;
	sram_mem[127748] = 16'b0000000000000000;
	sram_mem[127749] = 16'b0000000000000000;
	sram_mem[127750] = 16'b0000000000000000;
	sram_mem[127751] = 16'b0000000000000000;
	sram_mem[127752] = 16'b0000000000000000;
	sram_mem[127753] = 16'b0000000000000000;
	sram_mem[127754] = 16'b0000000000000000;
	sram_mem[127755] = 16'b0000000000000000;
	sram_mem[127756] = 16'b0000000000000000;
	sram_mem[127757] = 16'b0000000000000000;
	sram_mem[127758] = 16'b0000000000000000;
	sram_mem[127759] = 16'b0000000000000000;
	sram_mem[127760] = 16'b0000000000000000;
	sram_mem[127761] = 16'b0000000000000000;
	sram_mem[127762] = 16'b0000000000000000;
	sram_mem[127763] = 16'b0000000000000000;
	sram_mem[127764] = 16'b0000000000000000;
	sram_mem[127765] = 16'b0000000000000000;
	sram_mem[127766] = 16'b0000000000000000;
	sram_mem[127767] = 16'b0000000000000000;
	sram_mem[127768] = 16'b0000000000000000;
	sram_mem[127769] = 16'b0000000000000000;
	sram_mem[127770] = 16'b0000000000000000;
	sram_mem[127771] = 16'b0000000000000000;
	sram_mem[127772] = 16'b0000000000000000;
	sram_mem[127773] = 16'b0000000000000000;
	sram_mem[127774] = 16'b0000000000000000;
	sram_mem[127775] = 16'b0000000000000000;
	sram_mem[127776] = 16'b0000000000000000;
	sram_mem[127777] = 16'b0000000000000000;
	sram_mem[127778] = 16'b0000000000000000;
	sram_mem[127779] = 16'b0000000000000000;
	sram_mem[127780] = 16'b0000000000000000;
	sram_mem[127781] = 16'b0000000000000000;
	sram_mem[127782] = 16'b0000000000000000;
	sram_mem[127783] = 16'b0000000000000000;
	sram_mem[127784] = 16'b0000000000000000;
	sram_mem[127785] = 16'b0000000000000000;
	sram_mem[127786] = 16'b0000000000000000;
	sram_mem[127787] = 16'b0000000000000000;
	sram_mem[127788] = 16'b0000000000000000;
	sram_mem[127789] = 16'b0000000000000000;
	sram_mem[127790] = 16'b0000000000000000;
	sram_mem[127791] = 16'b0000000000000000;
	sram_mem[127792] = 16'b0000000000000000;
	sram_mem[127793] = 16'b0000000000000000;
	sram_mem[127794] = 16'b0000000000000000;
	sram_mem[127795] = 16'b0000000000000000;
	sram_mem[127796] = 16'b0000000000000000;
	sram_mem[127797] = 16'b0000000000000000;
	sram_mem[127798] = 16'b0000000000000000;
	sram_mem[127799] = 16'b0000000000000000;
	sram_mem[127800] = 16'b0000000000000000;
	sram_mem[127801] = 16'b0000000000000000;
	sram_mem[127802] = 16'b0000000000000000;
	sram_mem[127803] = 16'b0000000000000000;
	sram_mem[127804] = 16'b0000000000000000;
	sram_mem[127805] = 16'b0000000000000000;
	sram_mem[127806] = 16'b0000000000000000;
	sram_mem[127807] = 16'b0000000000000000;
	sram_mem[127808] = 16'b0000000000000000;
	sram_mem[127809] = 16'b0000000000000000;
	sram_mem[127810] = 16'b0000000000000000;
	sram_mem[127811] = 16'b0000000000000000;
	sram_mem[127812] = 16'b0000000000000000;
	sram_mem[127813] = 16'b0000000000000000;
	sram_mem[127814] = 16'b0000000000000000;
	sram_mem[127815] = 16'b0000000000000000;
	sram_mem[127816] = 16'b0000000000000000;
	sram_mem[127817] = 16'b0000000000000000;
	sram_mem[127818] = 16'b0000000000000000;
	sram_mem[127819] = 16'b0000000000000000;
	sram_mem[127820] = 16'b0000000000000000;
	sram_mem[127821] = 16'b0000000000000000;
	sram_mem[127822] = 16'b0000000000000000;
	sram_mem[127823] = 16'b0000000000000000;
	sram_mem[127824] = 16'b0000000000000000;
	sram_mem[127825] = 16'b0000000000000000;
	sram_mem[127826] = 16'b0000000000000000;
	sram_mem[127827] = 16'b0000000000000000;
	sram_mem[127828] = 16'b0000000000000000;
	sram_mem[127829] = 16'b0000000000000000;
	sram_mem[127830] = 16'b0000000000000000;
	sram_mem[127831] = 16'b0000000000000000;
	sram_mem[127832] = 16'b0000000000000000;
	sram_mem[127833] = 16'b0000000000000000;
	sram_mem[127834] = 16'b0000000000000000;
	sram_mem[127835] = 16'b0000000000000000;
	sram_mem[127836] = 16'b0000000000000000;
	sram_mem[127837] = 16'b0000000000000000;
	sram_mem[127838] = 16'b0000000000000000;
	sram_mem[127839] = 16'b0000000000000000;
	sram_mem[127840] = 16'b0000000000000000;
	sram_mem[127841] = 16'b0000000000000000;
	sram_mem[127842] = 16'b0000000000000000;
	sram_mem[127843] = 16'b0000000000000000;
	sram_mem[127844] = 16'b0000000000000000;
	sram_mem[127845] = 16'b0000000000000000;
	sram_mem[127846] = 16'b0000000000000000;
	sram_mem[127847] = 16'b0000000000000000;
	sram_mem[127848] = 16'b0000000000000000;
	sram_mem[127849] = 16'b0000000000000000;
	sram_mem[127850] = 16'b0000000000000000;
	sram_mem[127851] = 16'b0000000000000000;
	sram_mem[127852] = 16'b0000000000000000;
	sram_mem[127853] = 16'b0000000000000000;
	sram_mem[127854] = 16'b0000000000000000;
	sram_mem[127855] = 16'b0000000000000000;
	sram_mem[127856] = 16'b0000000000000000;
	sram_mem[127857] = 16'b0000000000000000;
	sram_mem[127858] = 16'b0000000000000000;
	sram_mem[127859] = 16'b0000000000000000;
	sram_mem[127860] = 16'b0000000000000000;
	sram_mem[127861] = 16'b0000000000000000;
	sram_mem[127862] = 16'b0000000000000000;
	sram_mem[127863] = 16'b0000000000000000;
	sram_mem[127864] = 16'b0000000000000000;
	sram_mem[127865] = 16'b0000000000000000;
	sram_mem[127866] = 16'b0000000000000000;
	sram_mem[127867] = 16'b0000000000000000;
	sram_mem[127868] = 16'b0000000000000000;
	sram_mem[127869] = 16'b0000000000000000;
	sram_mem[127870] = 16'b0000000000000000;
	sram_mem[127871] = 16'b0000000000000000;
	sram_mem[127872] = 16'b0000000000000000;
	sram_mem[127873] = 16'b0000000000000000;
	sram_mem[127874] = 16'b0000000000000000;
	sram_mem[127875] = 16'b0000000000000000;
	sram_mem[127876] = 16'b0000000000000000;
	sram_mem[127877] = 16'b0000000000000000;
	sram_mem[127878] = 16'b0000000000000000;
	sram_mem[127879] = 16'b0000000000000000;
	sram_mem[127880] = 16'b0000000000000000;
	sram_mem[127881] = 16'b0000000000000000;
	sram_mem[127882] = 16'b0000000000000000;
	sram_mem[127883] = 16'b0000000000000000;
	sram_mem[127884] = 16'b0000000000000000;
	sram_mem[127885] = 16'b0000000000000000;
	sram_mem[127886] = 16'b0000000000000000;
	sram_mem[127887] = 16'b0000000000000000;
	sram_mem[127888] = 16'b0000000000000000;
	sram_mem[127889] = 16'b0000000000000000;
	sram_mem[127890] = 16'b0000000000000000;
	sram_mem[127891] = 16'b0000000000000000;
	sram_mem[127892] = 16'b0000000000000000;
	sram_mem[127893] = 16'b0000000000000000;
	sram_mem[127894] = 16'b0000000000000000;
	sram_mem[127895] = 16'b0000000000000000;
	sram_mem[127896] = 16'b0000000000000000;
	sram_mem[127897] = 16'b0000000000000000;
	sram_mem[127898] = 16'b0000000000000000;
	sram_mem[127899] = 16'b0000000000000000;
	sram_mem[127900] = 16'b0000000000000000;
	sram_mem[127901] = 16'b0000000000000000;
	sram_mem[127902] = 16'b0000000000000000;
	sram_mem[127903] = 16'b0000000000000000;
	sram_mem[127904] = 16'b0000000000000000;
	sram_mem[127905] = 16'b0000000000000000;
	sram_mem[127906] = 16'b0000000000000000;
	sram_mem[127907] = 16'b0000000000000000;
	sram_mem[127908] = 16'b0000000000000000;
	sram_mem[127909] = 16'b0000000000000000;
	sram_mem[127910] = 16'b0000000000000000;
	sram_mem[127911] = 16'b0000000000000000;
	sram_mem[127912] = 16'b0000000000000000;
	sram_mem[127913] = 16'b0000000000000000;
	sram_mem[127914] = 16'b0000000000000000;
	sram_mem[127915] = 16'b0000000000000000;
	sram_mem[127916] = 16'b0000000000000000;
	sram_mem[127917] = 16'b0000000000000000;
	sram_mem[127918] = 16'b0000000000000000;
	sram_mem[127919] = 16'b0000000000000000;
	sram_mem[127920] = 16'b0000000000000000;
	sram_mem[127921] = 16'b0000000000000000;
	sram_mem[127922] = 16'b0000000000000000;
	sram_mem[127923] = 16'b0000000000000000;
	sram_mem[127924] = 16'b0000000000000000;
	sram_mem[127925] = 16'b0000000000000000;
	sram_mem[127926] = 16'b0000000000000000;
	sram_mem[127927] = 16'b0000000000000000;
	sram_mem[127928] = 16'b0000000000000000;
	sram_mem[127929] = 16'b0000000000000000;
	sram_mem[127930] = 16'b0000000000000000;
	sram_mem[127931] = 16'b0000000000000000;
	sram_mem[127932] = 16'b0000000000000000;
	sram_mem[127933] = 16'b0000000000000000;
	sram_mem[127934] = 16'b0000000000000000;
	sram_mem[127935] = 16'b0000000000000000;
	sram_mem[127936] = 16'b0000000000000000;
	sram_mem[127937] = 16'b0000000000000000;
	sram_mem[127938] = 16'b0000000000000000;
	sram_mem[127939] = 16'b0000000000000000;
	sram_mem[127940] = 16'b0000000000000000;
	sram_mem[127941] = 16'b0000000000000000;
	sram_mem[127942] = 16'b0000000000000000;
	sram_mem[127943] = 16'b0000000000000000;
	sram_mem[127944] = 16'b0000000000000000;
	sram_mem[127945] = 16'b0000000000000000;
	sram_mem[127946] = 16'b0000000000000000;
	sram_mem[127947] = 16'b0000000000000000;
	sram_mem[127948] = 16'b0000000000000000;
	sram_mem[127949] = 16'b0000000000000000;
	sram_mem[127950] = 16'b0000000000000000;
	sram_mem[127951] = 16'b0000000000000000;
	sram_mem[127952] = 16'b0000000000000000;
	sram_mem[127953] = 16'b0000000000000000;
	sram_mem[127954] = 16'b0000000000000000;
	sram_mem[127955] = 16'b0000000000000000;
	sram_mem[127956] = 16'b0000000000000000;
	sram_mem[127957] = 16'b0000000000000000;
	sram_mem[127958] = 16'b0000000000000000;
	sram_mem[127959] = 16'b0000000000000000;
	sram_mem[127960] = 16'b0000000000000000;
	sram_mem[127961] = 16'b0000000000000000;
	sram_mem[127962] = 16'b0000000000000000;
	sram_mem[127963] = 16'b0000000000000000;
	sram_mem[127964] = 16'b0000000000000000;
	sram_mem[127965] = 16'b0000000000000000;
	sram_mem[127966] = 16'b0000000000000000;
	sram_mem[127967] = 16'b0000000000000000;
	sram_mem[127968] = 16'b0000000000000000;
	sram_mem[127969] = 16'b0000000000000000;
	sram_mem[127970] = 16'b0000000000000000;
	sram_mem[127971] = 16'b0000000000000000;
	sram_mem[127972] = 16'b0000000000000000;
	sram_mem[127973] = 16'b0000000000000000;
	sram_mem[127974] = 16'b0000000000000000;
	sram_mem[127975] = 16'b0000000000000000;
	sram_mem[127976] = 16'b0000000000000000;
	sram_mem[127977] = 16'b0000000000000000;
	sram_mem[127978] = 16'b0000000000000000;
	sram_mem[127979] = 16'b0000000000000000;
	sram_mem[127980] = 16'b0000000000000000;
	sram_mem[127981] = 16'b0000000000000000;
	sram_mem[127982] = 16'b0000000000000000;
	sram_mem[127983] = 16'b0000000000000000;
	sram_mem[127984] = 16'b0000000000000000;
	sram_mem[127985] = 16'b0000000000000000;
	sram_mem[127986] = 16'b0000000000000000;
	sram_mem[127987] = 16'b0000000000000000;
	sram_mem[127988] = 16'b0000000000000000;
	sram_mem[127989] = 16'b0000000000000000;
	sram_mem[127990] = 16'b0000000000000000;
	sram_mem[127991] = 16'b0000000000000000;
	sram_mem[127992] = 16'b0000000000000000;
	sram_mem[127993] = 16'b0000000000000000;
	sram_mem[127994] = 16'b0000000000000000;
	sram_mem[127995] = 16'b0000000000000000;
	sram_mem[127996] = 16'b0000000000000000;
	sram_mem[127997] = 16'b0000000000000000;
	sram_mem[127998] = 16'b0000000000000000;
	sram_mem[127999] = 16'b0000000000000000;
	sram_mem[128000] = 16'b0000000000000000;
	sram_mem[128001] = 16'b0000000000000000;
	sram_mem[128002] = 16'b0000000000000000;
	sram_mem[128003] = 16'b0000000000000000;
	sram_mem[128004] = 16'b0000000000000000;
	sram_mem[128005] = 16'b0000000000000000;
	sram_mem[128006] = 16'b0000000000000000;
	sram_mem[128007] = 16'b0000000000000000;
	sram_mem[128008] = 16'b0000000000000000;
	sram_mem[128009] = 16'b0000000000000000;
	sram_mem[128010] = 16'b0000000000000000;
	sram_mem[128011] = 16'b0000000000000000;
	sram_mem[128012] = 16'b0000000000000000;
	sram_mem[128013] = 16'b0000000000000000;
	sram_mem[128014] = 16'b0000000000000000;
	sram_mem[128015] = 16'b0000000000000000;
	sram_mem[128016] = 16'b0000000000000000;
	sram_mem[128017] = 16'b0000000000000000;
	sram_mem[128018] = 16'b0000000000000000;
	sram_mem[128019] = 16'b0000000000000000;
	sram_mem[128020] = 16'b0000000000000000;
	sram_mem[128021] = 16'b0000000000000000;
	sram_mem[128022] = 16'b0000000000000000;
	sram_mem[128023] = 16'b0000000000000000;
	sram_mem[128024] = 16'b0000000000000000;
	sram_mem[128025] = 16'b0000000000000000;
	sram_mem[128026] = 16'b0000000000000000;
	sram_mem[128027] = 16'b0000000000000000;
	sram_mem[128028] = 16'b0000000000000000;
	sram_mem[128029] = 16'b0000000000000000;
	sram_mem[128030] = 16'b0000000000000000;
	sram_mem[128031] = 16'b0000000000000000;
	sram_mem[128032] = 16'b0000000000000000;
	sram_mem[128033] = 16'b0000000000000000;
	sram_mem[128034] = 16'b0000000000000000;
	sram_mem[128035] = 16'b0000000000000000;
	sram_mem[128036] = 16'b0000000000000000;
	sram_mem[128037] = 16'b0000000000000000;
	sram_mem[128038] = 16'b0000000000000000;
	sram_mem[128039] = 16'b0000000000000000;
	sram_mem[128040] = 16'b0000000000000000;
	sram_mem[128041] = 16'b0000000000000000;
	sram_mem[128042] = 16'b0000000000000000;
	sram_mem[128043] = 16'b0000000000000000;
	sram_mem[128044] = 16'b0000000000000000;
	sram_mem[128045] = 16'b0000000000000000;
	sram_mem[128046] = 16'b0000000000000000;
	sram_mem[128047] = 16'b0000000000000000;
	sram_mem[128048] = 16'b0000000000000000;
	sram_mem[128049] = 16'b0000000000000000;
	sram_mem[128050] = 16'b0000000000000000;
	sram_mem[128051] = 16'b0000000000000000;
	sram_mem[128052] = 16'b0000000000000000;
	sram_mem[128053] = 16'b0000000000000000;
	sram_mem[128054] = 16'b0000000000000000;
	sram_mem[128055] = 16'b0000000000000000;
	sram_mem[128056] = 16'b0000000000000000;
	sram_mem[128057] = 16'b0000000000000000;
	sram_mem[128058] = 16'b0000000000000000;
	sram_mem[128059] = 16'b0000000000000000;
	sram_mem[128060] = 16'b0000000000000000;
	sram_mem[128061] = 16'b0000000000000000;
	sram_mem[128062] = 16'b0000000000000000;
	sram_mem[128063] = 16'b0000000000000000;
	sram_mem[128064] = 16'b0000000000000000;
	sram_mem[128065] = 16'b0000000000000000;
	sram_mem[128066] = 16'b0000000000000000;
	sram_mem[128067] = 16'b0000000000000000;
	sram_mem[128068] = 16'b0000000000000000;
	sram_mem[128069] = 16'b0000000000000000;
	sram_mem[128070] = 16'b0000000000000000;
	sram_mem[128071] = 16'b0000000000000000;
	sram_mem[128072] = 16'b0000000000000000;
	sram_mem[128073] = 16'b0000000000000000;
	sram_mem[128074] = 16'b0000000000000000;
	sram_mem[128075] = 16'b0000000000000000;
	sram_mem[128076] = 16'b0000000000000000;
	sram_mem[128077] = 16'b0000000000000000;
	sram_mem[128078] = 16'b0000000000000000;
	sram_mem[128079] = 16'b0000000000000000;
	sram_mem[128080] = 16'b0000000000000000;
	sram_mem[128081] = 16'b0000000000000000;
	sram_mem[128082] = 16'b0000000000000000;
	sram_mem[128083] = 16'b0000000000000000;
	sram_mem[128084] = 16'b0000000000000000;
	sram_mem[128085] = 16'b0000000000000000;
	sram_mem[128086] = 16'b0000000000000000;
	sram_mem[128087] = 16'b0000000000000000;
	sram_mem[128088] = 16'b0000000000000000;
	sram_mem[128089] = 16'b0000000000000000;
	sram_mem[128090] = 16'b0000000000000000;
	sram_mem[128091] = 16'b0000000000000000;
	sram_mem[128092] = 16'b0000000000000000;
	sram_mem[128093] = 16'b0000000000000000;
	sram_mem[128094] = 16'b0000000000000000;
	sram_mem[128095] = 16'b0000000000000000;
	sram_mem[128096] = 16'b0000000000000000;
	sram_mem[128097] = 16'b0000000000000000;
	sram_mem[128098] = 16'b0000000000000000;
	sram_mem[128099] = 16'b0000000000000000;
	sram_mem[128100] = 16'b0000000000000000;
	sram_mem[128101] = 16'b0000000000000000;
	sram_mem[128102] = 16'b0000000000000000;
	sram_mem[128103] = 16'b0000000000000000;
	sram_mem[128104] = 16'b0000000000000000;
	sram_mem[128105] = 16'b0000000000000000;
	sram_mem[128106] = 16'b0000000000000000;
	sram_mem[128107] = 16'b0000000000000000;
	sram_mem[128108] = 16'b0000000000000000;
	sram_mem[128109] = 16'b0000000000000000;
	sram_mem[128110] = 16'b0000000000000000;
	sram_mem[128111] = 16'b0000000000000000;
	sram_mem[128112] = 16'b0000000000000000;
	sram_mem[128113] = 16'b0000000000000000;
	sram_mem[128114] = 16'b0000000000000000;
	sram_mem[128115] = 16'b0000000000000000;
	sram_mem[128116] = 16'b0000000000000000;
	sram_mem[128117] = 16'b0000000000000000;
	sram_mem[128118] = 16'b0000000000000000;
	sram_mem[128119] = 16'b0000000000000000;
	sram_mem[128120] = 16'b0000000000000000;
	sram_mem[128121] = 16'b0000000000000000;
	sram_mem[128122] = 16'b0000000000000000;
	sram_mem[128123] = 16'b0000000000000000;
	sram_mem[128124] = 16'b0000000000000000;
	sram_mem[128125] = 16'b0000000000000000;
	sram_mem[128126] = 16'b0000000000000000;
	sram_mem[128127] = 16'b0000000000000000;
	sram_mem[128128] = 16'b0000000000000000;
	sram_mem[128129] = 16'b0000000000000000;
	sram_mem[128130] = 16'b0000000000000000;
	sram_mem[128131] = 16'b0000000000000000;
	sram_mem[128132] = 16'b0000000000000000;
	sram_mem[128133] = 16'b0000000000000000;
	sram_mem[128134] = 16'b0000000000000000;
	sram_mem[128135] = 16'b0000000000000000;
	sram_mem[128136] = 16'b0000000000000000;
	sram_mem[128137] = 16'b0000000000000000;
	sram_mem[128138] = 16'b0000000000000000;
	sram_mem[128139] = 16'b0000000000000000;
	sram_mem[128140] = 16'b0000000000000000;
	sram_mem[128141] = 16'b0000000000000000;
	sram_mem[128142] = 16'b0000000000000000;
	sram_mem[128143] = 16'b0000000000000000;
	sram_mem[128144] = 16'b0000000000000000;
	sram_mem[128145] = 16'b0000000000000000;
	sram_mem[128146] = 16'b0000000000000000;
	sram_mem[128147] = 16'b0000000000000000;
	sram_mem[128148] = 16'b0000000000000000;
	sram_mem[128149] = 16'b0000000000000000;
	sram_mem[128150] = 16'b0000000000000000;
	sram_mem[128151] = 16'b0000000000000000;
	sram_mem[128152] = 16'b0000000000000000;
	sram_mem[128153] = 16'b0000000000000000;
	sram_mem[128154] = 16'b0000000000000000;
	sram_mem[128155] = 16'b0000000000000000;
	sram_mem[128156] = 16'b0000000000000000;
	sram_mem[128157] = 16'b0000000000000000;
	sram_mem[128158] = 16'b0000000000000000;
	sram_mem[128159] = 16'b0000000000000000;
	sram_mem[128160] = 16'b0000000000000000;
	sram_mem[128161] = 16'b0000000000000000;
	sram_mem[128162] = 16'b0000000000000000;
	sram_mem[128163] = 16'b0000000000000000;
	sram_mem[128164] = 16'b0000000000000000;
	sram_mem[128165] = 16'b0000000000000000;
	sram_mem[128166] = 16'b0000000000000000;
	sram_mem[128167] = 16'b0000000000000000;
	sram_mem[128168] = 16'b0000000000000000;
	sram_mem[128169] = 16'b0000000000000000;
	sram_mem[128170] = 16'b0000000000000000;
	sram_mem[128171] = 16'b0000000000000000;
	sram_mem[128172] = 16'b0000000000000000;
	sram_mem[128173] = 16'b0000000000000000;
	sram_mem[128174] = 16'b0000000000000000;
	sram_mem[128175] = 16'b0000000000000000;
	sram_mem[128176] = 16'b0000000000000000;
	sram_mem[128177] = 16'b0000000000000000;
	sram_mem[128178] = 16'b0000000000000000;
	sram_mem[128179] = 16'b0000000000000000;
	sram_mem[128180] = 16'b0000000000000000;
	sram_mem[128181] = 16'b0000000000000000;
	sram_mem[128182] = 16'b0000000000000000;
	sram_mem[128183] = 16'b0000000000000000;
	sram_mem[128184] = 16'b0000000000000000;
	sram_mem[128185] = 16'b0000000000000000;
	sram_mem[128186] = 16'b0000000000000000;
	sram_mem[128187] = 16'b0000000000000000;
	sram_mem[128188] = 16'b0000000000000000;
	sram_mem[128189] = 16'b0000000000000000;
	sram_mem[128190] = 16'b0000000000000000;
	sram_mem[128191] = 16'b0000000000000000;
	sram_mem[128192] = 16'b0000000000000000;
	sram_mem[128193] = 16'b0000000000000000;
	sram_mem[128194] = 16'b0000000000000000;
	sram_mem[128195] = 16'b0000000000000000;
	sram_mem[128196] = 16'b0000000000000000;
	sram_mem[128197] = 16'b0000000000000000;
	sram_mem[128198] = 16'b0000000000000000;
	sram_mem[128199] = 16'b0000000000000000;
	sram_mem[128200] = 16'b0000000000000000;
	sram_mem[128201] = 16'b0000000000000000;
	sram_mem[128202] = 16'b0000000000000000;
	sram_mem[128203] = 16'b0000000000000000;
	sram_mem[128204] = 16'b0000000000000000;
	sram_mem[128205] = 16'b0000000000000000;
	sram_mem[128206] = 16'b0000000000000000;
	sram_mem[128207] = 16'b0000000000000000;
	sram_mem[128208] = 16'b0000000000000000;
	sram_mem[128209] = 16'b0000000000000000;
	sram_mem[128210] = 16'b0000000000000000;
	sram_mem[128211] = 16'b0000000000000000;
	sram_mem[128212] = 16'b0000000000000000;
	sram_mem[128213] = 16'b0000000000000000;
	sram_mem[128214] = 16'b0000000000000000;
	sram_mem[128215] = 16'b0000000000000000;
	sram_mem[128216] = 16'b0000000000000000;
	sram_mem[128217] = 16'b0000000000000000;
	sram_mem[128218] = 16'b0000000000000000;
	sram_mem[128219] = 16'b0000000000000000;
	sram_mem[128220] = 16'b0000000000000000;
	sram_mem[128221] = 16'b0000000000000000;
	sram_mem[128222] = 16'b0000000000000000;
	sram_mem[128223] = 16'b0000000000000000;
	sram_mem[128224] = 16'b0000000000000000;
	sram_mem[128225] = 16'b0000000000000000;
	sram_mem[128226] = 16'b0000000000000000;
	sram_mem[128227] = 16'b0000000000000000;
	sram_mem[128228] = 16'b0000000000000000;
	sram_mem[128229] = 16'b0000000000000000;
	sram_mem[128230] = 16'b0000000000000000;
	sram_mem[128231] = 16'b0000000000000000;
	sram_mem[128232] = 16'b0000000000000000;
	sram_mem[128233] = 16'b0000000000000000;
	sram_mem[128234] = 16'b0000000000000000;
	sram_mem[128235] = 16'b0000000000000000;
	sram_mem[128236] = 16'b0000000000000000;
	sram_mem[128237] = 16'b0000000000000000;
	sram_mem[128238] = 16'b0000000000000000;
	sram_mem[128239] = 16'b0000000000000000;
	sram_mem[128240] = 16'b0000000000000000;
	sram_mem[128241] = 16'b0000000000000000;
	sram_mem[128242] = 16'b0000000000000000;
	sram_mem[128243] = 16'b0000000000000000;
	sram_mem[128244] = 16'b0000000000000000;
	sram_mem[128245] = 16'b0000000000000000;
	sram_mem[128246] = 16'b0000000000000000;
	sram_mem[128247] = 16'b0000000000000000;
	sram_mem[128248] = 16'b0000000000000000;
	sram_mem[128249] = 16'b0000000000000000;
	sram_mem[128250] = 16'b0000000000000000;
	sram_mem[128251] = 16'b0000000000000000;
	sram_mem[128252] = 16'b0000000000000000;
	sram_mem[128253] = 16'b0000000000000000;
	sram_mem[128254] = 16'b0000000000000000;
	sram_mem[128255] = 16'b0000000000000000;
	sram_mem[128256] = 16'b0000000000000000;
	sram_mem[128257] = 16'b0000000000000000;
	sram_mem[128258] = 16'b0000000000000000;
	sram_mem[128259] = 16'b0000000000000000;
	sram_mem[128260] = 16'b0000000000000000;
	sram_mem[128261] = 16'b0000000000000000;
	sram_mem[128262] = 16'b0000000000000000;
	sram_mem[128263] = 16'b0000000000000000;
	sram_mem[128264] = 16'b0000000000000000;
	sram_mem[128265] = 16'b0000000000000000;
	sram_mem[128266] = 16'b0000000000000000;
	sram_mem[128267] = 16'b0000000000000000;
	sram_mem[128268] = 16'b0000000000000000;
	sram_mem[128269] = 16'b0000000000000000;
	sram_mem[128270] = 16'b0000000000000000;
	sram_mem[128271] = 16'b0000000000000000;
	sram_mem[128272] = 16'b0000000000000000;
	sram_mem[128273] = 16'b0000000000000000;
	sram_mem[128274] = 16'b0000000000000000;
	sram_mem[128275] = 16'b0000000000000000;
	sram_mem[128276] = 16'b0000000000000000;
	sram_mem[128277] = 16'b0000000000000000;
	sram_mem[128278] = 16'b0000000000000000;
	sram_mem[128279] = 16'b0000000000000000;
	sram_mem[128280] = 16'b0000000000000000;
	sram_mem[128281] = 16'b0000000000000000;
	sram_mem[128282] = 16'b0000000000000000;
	sram_mem[128283] = 16'b0000000000000000;
	sram_mem[128284] = 16'b0000000000000000;
	sram_mem[128285] = 16'b0000000000000000;
	sram_mem[128286] = 16'b0000000000000000;
	sram_mem[128287] = 16'b0000000000000000;
	sram_mem[128288] = 16'b0000000000000000;
	sram_mem[128289] = 16'b0000000000000000;
	sram_mem[128290] = 16'b0000000000000000;
	sram_mem[128291] = 16'b0000000000000000;
	sram_mem[128292] = 16'b0000000000000000;
	sram_mem[128293] = 16'b0000000000000000;
	sram_mem[128294] = 16'b0000000000000000;
	sram_mem[128295] = 16'b0000000000000000;
	sram_mem[128296] = 16'b0000000000000000;
	sram_mem[128297] = 16'b0000000000000000;
	sram_mem[128298] = 16'b0000000000000000;
	sram_mem[128299] = 16'b0000000000000000;
	sram_mem[128300] = 16'b0000000000000000;
	sram_mem[128301] = 16'b0000000000000000;
	sram_mem[128302] = 16'b0000000000000000;
	sram_mem[128303] = 16'b0000000000000000;
	sram_mem[128304] = 16'b0000000000000000;
	sram_mem[128305] = 16'b0000000000000000;
	sram_mem[128306] = 16'b0000000000000000;
	sram_mem[128307] = 16'b0000000000000000;
	sram_mem[128308] = 16'b0000000000000000;
	sram_mem[128309] = 16'b0000000000000000;
	sram_mem[128310] = 16'b0000000000000000;
	sram_mem[128311] = 16'b0000000000000000;
	sram_mem[128312] = 16'b0000000000000000;
	sram_mem[128313] = 16'b0000000000000000;
	sram_mem[128314] = 16'b0000000000000000;
	sram_mem[128315] = 16'b0000000000000000;
	sram_mem[128316] = 16'b0000000000000000;
	sram_mem[128317] = 16'b0000000000000000;
	sram_mem[128318] = 16'b0000000000000000;
	sram_mem[128319] = 16'b0000000000000000;
	sram_mem[128320] = 16'b0000000000000000;
	sram_mem[128321] = 16'b0000000000000000;
	sram_mem[128322] = 16'b0000000000000000;
	sram_mem[128323] = 16'b0000000000000000;
	sram_mem[128324] = 16'b0000000000000000;
	sram_mem[128325] = 16'b0000000000000000;
	sram_mem[128326] = 16'b0000000000000000;
	sram_mem[128327] = 16'b0000000000000000;
	sram_mem[128328] = 16'b0000000000000000;
	sram_mem[128329] = 16'b0000000000000000;
	sram_mem[128330] = 16'b0000000000000000;
	sram_mem[128331] = 16'b0000000000000000;
	sram_mem[128332] = 16'b0000000000000000;
	sram_mem[128333] = 16'b0000000000000000;
	sram_mem[128334] = 16'b0000000000000000;
	sram_mem[128335] = 16'b0000000000000000;
	sram_mem[128336] = 16'b0000000000000000;
	sram_mem[128337] = 16'b0000000000000000;
	sram_mem[128338] = 16'b0000000000000000;
	sram_mem[128339] = 16'b0000000000000000;
	sram_mem[128340] = 16'b0000000000000000;
	sram_mem[128341] = 16'b0000000000000000;
	sram_mem[128342] = 16'b0000000000000000;
	sram_mem[128343] = 16'b0000000000000000;
	sram_mem[128344] = 16'b0000000000000000;
	sram_mem[128345] = 16'b0000000000000000;
	sram_mem[128346] = 16'b0000000000000000;
	sram_mem[128347] = 16'b0000000000000000;
	sram_mem[128348] = 16'b0000000000000000;
	sram_mem[128349] = 16'b0000000000000000;
	sram_mem[128350] = 16'b0000000000000000;
	sram_mem[128351] = 16'b0000000000000000;
	sram_mem[128352] = 16'b0000000000000000;
	sram_mem[128353] = 16'b0000000000000000;
	sram_mem[128354] = 16'b0000000000000000;
	sram_mem[128355] = 16'b0000000000000000;
	sram_mem[128356] = 16'b0000000000000000;
	sram_mem[128357] = 16'b0000000000000000;
	sram_mem[128358] = 16'b0000000000000000;
	sram_mem[128359] = 16'b0000000000000000;
	sram_mem[128360] = 16'b0000000000000000;
	sram_mem[128361] = 16'b0000000000000000;
	sram_mem[128362] = 16'b0000000000000000;
	sram_mem[128363] = 16'b0000000000000000;
	sram_mem[128364] = 16'b0000000000000000;
	sram_mem[128365] = 16'b0000000000000000;
	sram_mem[128366] = 16'b0000000000000000;
	sram_mem[128367] = 16'b0000000000000000;
	sram_mem[128368] = 16'b0000000000000000;
	sram_mem[128369] = 16'b0000000000000000;
	sram_mem[128370] = 16'b0000000000000000;
	sram_mem[128371] = 16'b0000000000000000;
	sram_mem[128372] = 16'b0000000000000000;
	sram_mem[128373] = 16'b0000000000000000;
	sram_mem[128374] = 16'b0000000000000000;
	sram_mem[128375] = 16'b0000000000000000;
	sram_mem[128376] = 16'b0000000000000000;
	sram_mem[128377] = 16'b0000000000000000;
	sram_mem[128378] = 16'b0000000000000000;
	sram_mem[128379] = 16'b0000000000000000;
	sram_mem[128380] = 16'b0000000000000000;
	sram_mem[128381] = 16'b0000000000000000;
	sram_mem[128382] = 16'b0000000000000000;
	sram_mem[128383] = 16'b0000000000000000;
	sram_mem[128384] = 16'b0000000000000000;
	sram_mem[128385] = 16'b0000000000000000;
	sram_mem[128386] = 16'b0000000000000000;
	sram_mem[128387] = 16'b0000000000000000;
	sram_mem[128388] = 16'b0000000000000000;
	sram_mem[128389] = 16'b0000000000000000;
	sram_mem[128390] = 16'b0000000000000000;
	sram_mem[128391] = 16'b0000000000000000;
	sram_mem[128392] = 16'b0000000000000000;
	sram_mem[128393] = 16'b0000000000000000;
	sram_mem[128394] = 16'b0000000000000000;
	sram_mem[128395] = 16'b0000000000000000;
	sram_mem[128396] = 16'b0000000000000000;
	sram_mem[128397] = 16'b0000000000000000;
	sram_mem[128398] = 16'b0000000000000000;
	sram_mem[128399] = 16'b0000000000000000;
	sram_mem[128400] = 16'b0000000000000000;
	sram_mem[128401] = 16'b0000000000000000;
	sram_mem[128402] = 16'b0000000000000000;
	sram_mem[128403] = 16'b0000000000000000;
	sram_mem[128404] = 16'b0000000000000000;
	sram_mem[128405] = 16'b0000000000000000;
	sram_mem[128406] = 16'b0000000000000000;
	sram_mem[128407] = 16'b0000000000000000;
	sram_mem[128408] = 16'b0000000000000000;
	sram_mem[128409] = 16'b0000000000000000;
	sram_mem[128410] = 16'b0000000000000000;
	sram_mem[128411] = 16'b0000000000000000;
	sram_mem[128412] = 16'b0000000000000000;
	sram_mem[128413] = 16'b0000000000000000;
	sram_mem[128414] = 16'b0000000000000000;
	sram_mem[128415] = 16'b0000000000000000;
	sram_mem[128416] = 16'b0000000000000000;
	sram_mem[128417] = 16'b0000000000000000;
	sram_mem[128418] = 16'b0000000000000000;
	sram_mem[128419] = 16'b0000000000000000;
	sram_mem[128420] = 16'b0000000000000000;
	sram_mem[128421] = 16'b0000000000000000;
	sram_mem[128422] = 16'b0000000000000000;
	sram_mem[128423] = 16'b0000000000000000;
	sram_mem[128424] = 16'b0000000000000000;
	sram_mem[128425] = 16'b0000000000000000;
	sram_mem[128426] = 16'b0000000000000000;
	sram_mem[128427] = 16'b0000000000000000;
	sram_mem[128428] = 16'b0000000000000000;
	sram_mem[128429] = 16'b0000000000000000;
	sram_mem[128430] = 16'b0000000000000000;
	sram_mem[128431] = 16'b0000000000000000;
	sram_mem[128432] = 16'b0000000000000000;
	sram_mem[128433] = 16'b0000000000000000;
	sram_mem[128434] = 16'b0000000000000000;
	sram_mem[128435] = 16'b0000000000000000;
	sram_mem[128436] = 16'b0000000000000000;
	sram_mem[128437] = 16'b0000000000000000;
	sram_mem[128438] = 16'b0000000000000000;
	sram_mem[128439] = 16'b0000000000000000;
	sram_mem[128440] = 16'b0000000000000000;
	sram_mem[128441] = 16'b0000000000000000;
	sram_mem[128442] = 16'b0000000000000000;
	sram_mem[128443] = 16'b0000000000000000;
	sram_mem[128444] = 16'b0000000000000000;
	sram_mem[128445] = 16'b0000000000000000;
	sram_mem[128446] = 16'b0000000000000000;
	sram_mem[128447] = 16'b0000000000000000;
	sram_mem[128448] = 16'b0000000000000000;
	sram_mem[128449] = 16'b0000000000000000;
	sram_mem[128450] = 16'b0000000000000000;
	sram_mem[128451] = 16'b0000000000000000;
	sram_mem[128452] = 16'b0000000000000000;
	sram_mem[128453] = 16'b0000000000000000;
	sram_mem[128454] = 16'b0000000000000000;
	sram_mem[128455] = 16'b0000000000000000;
	sram_mem[128456] = 16'b0000000000000000;
	sram_mem[128457] = 16'b0000000000000000;
	sram_mem[128458] = 16'b0000000000000000;
	sram_mem[128459] = 16'b0000000000000000;
	sram_mem[128460] = 16'b0000000000000000;
	sram_mem[128461] = 16'b0000000000000000;
	sram_mem[128462] = 16'b0000000000000000;
	sram_mem[128463] = 16'b0000000000000000;
	sram_mem[128464] = 16'b0000000000000000;
	sram_mem[128465] = 16'b0000000000000000;
	sram_mem[128466] = 16'b0000000000000000;
	sram_mem[128467] = 16'b0000000000000000;
	sram_mem[128468] = 16'b0000000000000000;
	sram_mem[128469] = 16'b0000000000000000;
	sram_mem[128470] = 16'b0000000000000000;
	sram_mem[128471] = 16'b0000000000000000;
	sram_mem[128472] = 16'b0000000000000000;
	sram_mem[128473] = 16'b0000000000000000;
	sram_mem[128474] = 16'b0000000000000000;
	sram_mem[128475] = 16'b0000000000000000;
	sram_mem[128476] = 16'b0000000000000000;
	sram_mem[128477] = 16'b0000000000000000;
	sram_mem[128478] = 16'b0000000000000000;
	sram_mem[128479] = 16'b0000000000000000;
	sram_mem[128480] = 16'b0000000000000000;
	sram_mem[128481] = 16'b0000000000000000;
	sram_mem[128482] = 16'b0000000000000000;
	sram_mem[128483] = 16'b0000000000000000;
	sram_mem[128484] = 16'b0000000000000000;
	sram_mem[128485] = 16'b0000000000000000;
	sram_mem[128486] = 16'b0000000000000000;
	sram_mem[128487] = 16'b0000000000000000;
	sram_mem[128488] = 16'b0000000000000000;
	sram_mem[128489] = 16'b0000000000000000;
	sram_mem[128490] = 16'b0000000000000000;
	sram_mem[128491] = 16'b0000000000000000;
	sram_mem[128492] = 16'b0000000000000000;
	sram_mem[128493] = 16'b0000000000000000;
	sram_mem[128494] = 16'b0000000000000000;
	sram_mem[128495] = 16'b0000000000000000;
	sram_mem[128496] = 16'b0000000000000000;
	sram_mem[128497] = 16'b0000000000000000;
	sram_mem[128498] = 16'b0000000000000000;
	sram_mem[128499] = 16'b0000000000000000;
	sram_mem[128500] = 16'b0000000000000000;
	sram_mem[128501] = 16'b0000000000000000;
	sram_mem[128502] = 16'b0000000000000000;
	sram_mem[128503] = 16'b0000000000000000;
	sram_mem[128504] = 16'b0000000000000000;
	sram_mem[128505] = 16'b0000000000000000;
	sram_mem[128506] = 16'b0000000000000000;
	sram_mem[128507] = 16'b0000000000000000;
	sram_mem[128508] = 16'b0000000000000000;
	sram_mem[128509] = 16'b0000000000000000;
	sram_mem[128510] = 16'b0000000000000000;
	sram_mem[128511] = 16'b0000000000000000;
	sram_mem[128512] = 16'b0000000000000000;
	sram_mem[128513] = 16'b0000000000000000;
	sram_mem[128514] = 16'b0000000000000000;
	sram_mem[128515] = 16'b0000000000000000;
	sram_mem[128516] = 16'b0000000000000000;
	sram_mem[128517] = 16'b0000000000000000;
	sram_mem[128518] = 16'b0000000000000000;
	sram_mem[128519] = 16'b0000000000000000;
	sram_mem[128520] = 16'b0000000000000000;
	sram_mem[128521] = 16'b0000000000000000;
	sram_mem[128522] = 16'b0000000000000000;
	sram_mem[128523] = 16'b0000000000000000;
	sram_mem[128524] = 16'b0000000000000000;
	sram_mem[128525] = 16'b0000000000000000;
	sram_mem[128526] = 16'b0000000000000000;
	sram_mem[128527] = 16'b0000000000000000;
	sram_mem[128528] = 16'b0000000000000000;
	sram_mem[128529] = 16'b0000000000000000;
	sram_mem[128530] = 16'b0000000000000000;
	sram_mem[128531] = 16'b0000000000000000;
	sram_mem[128532] = 16'b0000000000000000;
	sram_mem[128533] = 16'b0000000000000000;
	sram_mem[128534] = 16'b0000000000000000;
	sram_mem[128535] = 16'b0000000000000000;
	sram_mem[128536] = 16'b0000000000000000;
	sram_mem[128537] = 16'b0000000000000000;
	sram_mem[128538] = 16'b0000000000000000;
	sram_mem[128539] = 16'b0000000000000000;
	sram_mem[128540] = 16'b0000000000000000;
	sram_mem[128541] = 16'b0000000000000000;
	sram_mem[128542] = 16'b0000000000000000;
	sram_mem[128543] = 16'b0000000000000000;
	sram_mem[128544] = 16'b0000000000000000;
	sram_mem[128545] = 16'b0000000000000000;
	sram_mem[128546] = 16'b0000000000000000;
	sram_mem[128547] = 16'b0000000000000000;
	sram_mem[128548] = 16'b0000000000000000;
	sram_mem[128549] = 16'b0000000000000000;
	sram_mem[128550] = 16'b0000000000000000;
	sram_mem[128551] = 16'b0000000000000000;
	sram_mem[128552] = 16'b0000000000000000;
	sram_mem[128553] = 16'b0000000000000000;
	sram_mem[128554] = 16'b0000000000000000;
	sram_mem[128555] = 16'b0000000000000000;
	sram_mem[128556] = 16'b0000000000000000;
	sram_mem[128557] = 16'b0000000000000000;
	sram_mem[128558] = 16'b0000000000000000;
	sram_mem[128559] = 16'b0000000000000000;
	sram_mem[128560] = 16'b0000000000000000;
	sram_mem[128561] = 16'b0000000000000000;
	sram_mem[128562] = 16'b0000000000000000;
	sram_mem[128563] = 16'b0000000000000000;
	sram_mem[128564] = 16'b0000000000000000;
	sram_mem[128565] = 16'b0000000000000000;
	sram_mem[128566] = 16'b0000000000000000;
	sram_mem[128567] = 16'b0000000000000000;
	sram_mem[128568] = 16'b0000000000000000;
	sram_mem[128569] = 16'b0000000000000000;
	sram_mem[128570] = 16'b0000000000000000;
	sram_mem[128571] = 16'b0000000000000000;
	sram_mem[128572] = 16'b0000000000000000;
	sram_mem[128573] = 16'b0000000000000000;
	sram_mem[128574] = 16'b0000000000000000;
	sram_mem[128575] = 16'b0000000000000000;
	sram_mem[128576] = 16'b0000000000000000;
	sram_mem[128577] = 16'b0000000000000000;
	sram_mem[128578] = 16'b0000000000000000;
	sram_mem[128579] = 16'b0000000000000000;
	sram_mem[128580] = 16'b0000000000000000;
	sram_mem[128581] = 16'b0000000000000000;
	sram_mem[128582] = 16'b0000000000000000;
	sram_mem[128583] = 16'b0000000000000000;
	sram_mem[128584] = 16'b0000000000000000;
	sram_mem[128585] = 16'b0000000000000000;
	sram_mem[128586] = 16'b0000000000000000;
	sram_mem[128587] = 16'b0000000000000000;
	sram_mem[128588] = 16'b0000000000000000;
	sram_mem[128589] = 16'b0000000000000000;
	sram_mem[128590] = 16'b0000000000000000;
	sram_mem[128591] = 16'b0000000000000000;
	sram_mem[128592] = 16'b0000000000000000;
	sram_mem[128593] = 16'b0000000000000000;
	sram_mem[128594] = 16'b0000000000000000;
	sram_mem[128595] = 16'b0000000000000000;
	sram_mem[128596] = 16'b0000000000000000;
	sram_mem[128597] = 16'b0000000000000000;
	sram_mem[128598] = 16'b0000000000000000;
	sram_mem[128599] = 16'b0000000000000000;
	sram_mem[128600] = 16'b0000000000000000;
	sram_mem[128601] = 16'b0000000000000000;
	sram_mem[128602] = 16'b0000000000000000;
	sram_mem[128603] = 16'b0000000000000000;
	sram_mem[128604] = 16'b0000000000000000;
	sram_mem[128605] = 16'b0000000000000000;
	sram_mem[128606] = 16'b0000000000000000;
	sram_mem[128607] = 16'b0000000000000000;
	sram_mem[128608] = 16'b0000000000000000;
	sram_mem[128609] = 16'b0000000000000000;
	sram_mem[128610] = 16'b0000000000000000;
	sram_mem[128611] = 16'b0000000000000000;
	sram_mem[128612] = 16'b0000000000000000;
	sram_mem[128613] = 16'b0000000000000000;
	sram_mem[128614] = 16'b0000000000000000;
	sram_mem[128615] = 16'b0000000000000000;
	sram_mem[128616] = 16'b0000000000000000;
	sram_mem[128617] = 16'b0000000000000000;
	sram_mem[128618] = 16'b0000000000000000;
	sram_mem[128619] = 16'b0000000000000000;
	sram_mem[128620] = 16'b0000000000000000;
	sram_mem[128621] = 16'b0000000000000000;
	sram_mem[128622] = 16'b0000000000000000;
	sram_mem[128623] = 16'b0000000000000000;
	sram_mem[128624] = 16'b0000000000000000;
	sram_mem[128625] = 16'b0000000000000000;
	sram_mem[128626] = 16'b0000000000000000;
	sram_mem[128627] = 16'b0000000000000000;
	sram_mem[128628] = 16'b0000000000000000;
	sram_mem[128629] = 16'b0000000000000000;
	sram_mem[128630] = 16'b0000000000000000;
	sram_mem[128631] = 16'b0000000000000000;
	sram_mem[128632] = 16'b0000000000000000;
	sram_mem[128633] = 16'b0000000000000000;
	sram_mem[128634] = 16'b0000000000000000;
	sram_mem[128635] = 16'b0000000000000000;
	sram_mem[128636] = 16'b0000000000000000;
	sram_mem[128637] = 16'b0000000000000000;
	sram_mem[128638] = 16'b0000000000000000;
	sram_mem[128639] = 16'b0000000000000000;
	sram_mem[128640] = 16'b0000000000000000;
	sram_mem[128641] = 16'b0000000000000000;
	sram_mem[128642] = 16'b0000000000000000;
	sram_mem[128643] = 16'b0000000000000000;
	sram_mem[128644] = 16'b0000000000000000;
	sram_mem[128645] = 16'b0000000000000000;
	sram_mem[128646] = 16'b0000000000000000;
	sram_mem[128647] = 16'b0000000000000000;
	sram_mem[128648] = 16'b0000000000000000;
	sram_mem[128649] = 16'b0000000000000000;
	sram_mem[128650] = 16'b0000000000000000;
	sram_mem[128651] = 16'b0000000000000000;
	sram_mem[128652] = 16'b0000000000000000;
	sram_mem[128653] = 16'b0000000000000000;
	sram_mem[128654] = 16'b0000000000000000;
	sram_mem[128655] = 16'b0000000000000000;
	sram_mem[128656] = 16'b0000000000000000;
	sram_mem[128657] = 16'b0000000000000000;
	sram_mem[128658] = 16'b0000000000000000;
	sram_mem[128659] = 16'b0000000000000000;
	sram_mem[128660] = 16'b0000000000000000;
	sram_mem[128661] = 16'b0000000000000000;
	sram_mem[128662] = 16'b0000000000000000;
	sram_mem[128663] = 16'b0000000000000000;
	sram_mem[128664] = 16'b0000000000000000;
	sram_mem[128665] = 16'b0000000000000000;
	sram_mem[128666] = 16'b0000000000000000;
	sram_mem[128667] = 16'b0000000000000000;
	sram_mem[128668] = 16'b0000000000000000;
	sram_mem[128669] = 16'b0000000000000000;
	sram_mem[128670] = 16'b0000000000000000;
	sram_mem[128671] = 16'b0000000000000000;
	sram_mem[128672] = 16'b0000000000000000;
	sram_mem[128673] = 16'b0000000000000000;
	sram_mem[128674] = 16'b0000000000000000;
	sram_mem[128675] = 16'b0000000000000000;
	sram_mem[128676] = 16'b0000000000000000;
	sram_mem[128677] = 16'b0000000000000000;
	sram_mem[128678] = 16'b0000000000000000;
	sram_mem[128679] = 16'b0000000000000000;
	sram_mem[128680] = 16'b0000000000000000;
	sram_mem[128681] = 16'b0000000000000000;
	sram_mem[128682] = 16'b0000000000000000;
	sram_mem[128683] = 16'b0000000000000000;
	sram_mem[128684] = 16'b0000000000000000;
	sram_mem[128685] = 16'b0000000000000000;
	sram_mem[128686] = 16'b0000000000000000;
	sram_mem[128687] = 16'b0000000000000000;
	sram_mem[128688] = 16'b0000000000000000;
	sram_mem[128689] = 16'b0000000000000000;
	sram_mem[128690] = 16'b0000000000000000;
	sram_mem[128691] = 16'b0000000000000000;
	sram_mem[128692] = 16'b0000000000000000;
	sram_mem[128693] = 16'b0000000000000000;
	sram_mem[128694] = 16'b0000000000000000;
	sram_mem[128695] = 16'b0000000000000000;
	sram_mem[128696] = 16'b0000000000000000;
	sram_mem[128697] = 16'b0000000000000000;
	sram_mem[128698] = 16'b0000000000000000;
	sram_mem[128699] = 16'b0000000000000000;
	sram_mem[128700] = 16'b0000000000000000;
	sram_mem[128701] = 16'b0000000000000000;
	sram_mem[128702] = 16'b0000000000000000;
	sram_mem[128703] = 16'b0000000000000000;
	sram_mem[128704] = 16'b0000000000000000;
	sram_mem[128705] = 16'b0000000000000000;
	sram_mem[128706] = 16'b0000000000000000;
	sram_mem[128707] = 16'b0000000000000000;
	sram_mem[128708] = 16'b0000000000000000;
	sram_mem[128709] = 16'b0000000000000000;
	sram_mem[128710] = 16'b0000000000000000;
	sram_mem[128711] = 16'b0000000000000000;
	sram_mem[128712] = 16'b0000000000000000;
	sram_mem[128713] = 16'b0000000000000000;
	sram_mem[128714] = 16'b0000000000000000;
	sram_mem[128715] = 16'b0000000000000000;
	sram_mem[128716] = 16'b0000000000000000;
	sram_mem[128717] = 16'b0000000000000000;
	sram_mem[128718] = 16'b0000000000000000;
	sram_mem[128719] = 16'b0000000000000000;
	sram_mem[128720] = 16'b0000000000000000;
	sram_mem[128721] = 16'b0000000000000000;
	sram_mem[128722] = 16'b0000000000000000;
	sram_mem[128723] = 16'b0000000000000000;
	sram_mem[128724] = 16'b0000000000000000;
	sram_mem[128725] = 16'b0000000000000000;
	sram_mem[128726] = 16'b0000000000000000;
	sram_mem[128727] = 16'b0000000000000000;
	sram_mem[128728] = 16'b0000000000000000;
	sram_mem[128729] = 16'b0000000000000000;
	sram_mem[128730] = 16'b0000000000000000;
	sram_mem[128731] = 16'b0000000000000000;
	sram_mem[128732] = 16'b0000000000000000;
	sram_mem[128733] = 16'b0000000000000000;
	sram_mem[128734] = 16'b0000000000000000;
	sram_mem[128735] = 16'b0000000000000000;
	sram_mem[128736] = 16'b0000000000000000;
	sram_mem[128737] = 16'b0000000000000000;
	sram_mem[128738] = 16'b0000000000000000;
	sram_mem[128739] = 16'b0000000000000000;
	sram_mem[128740] = 16'b0000000000000000;
	sram_mem[128741] = 16'b0000000000000000;
	sram_mem[128742] = 16'b0000000000000000;
	sram_mem[128743] = 16'b0000000000000000;
	sram_mem[128744] = 16'b0000000000000000;
	sram_mem[128745] = 16'b0000000000000000;
	sram_mem[128746] = 16'b0000000000000000;
	sram_mem[128747] = 16'b0000000000000000;
	sram_mem[128748] = 16'b0000000000000000;
	sram_mem[128749] = 16'b0000000000000000;
	sram_mem[128750] = 16'b0000000000000000;
	sram_mem[128751] = 16'b0000000000000000;
	sram_mem[128752] = 16'b0000000000000000;
	sram_mem[128753] = 16'b0000000000000000;
	sram_mem[128754] = 16'b0000000000000000;
	sram_mem[128755] = 16'b0000000000000000;
	sram_mem[128756] = 16'b0000000000000000;
	sram_mem[128757] = 16'b0000000000000000;
	sram_mem[128758] = 16'b0000000000000000;
	sram_mem[128759] = 16'b0000000000000000;
	sram_mem[128760] = 16'b0000000000000000;
	sram_mem[128761] = 16'b0000000000000000;
	sram_mem[128762] = 16'b0000000000000000;
	sram_mem[128763] = 16'b0000000000000000;
	sram_mem[128764] = 16'b0000000000000000;
	sram_mem[128765] = 16'b0000000000000000;
	sram_mem[128766] = 16'b0000000000000000;
	sram_mem[128767] = 16'b0000000000000000;
	sram_mem[128768] = 16'b0000000000000000;
	sram_mem[128769] = 16'b0000000000000000;
	sram_mem[128770] = 16'b0000000000000000;
	sram_mem[128771] = 16'b0000000000000000;
	sram_mem[128772] = 16'b0000000000000000;
	sram_mem[128773] = 16'b0000000000000000;
	sram_mem[128774] = 16'b0000000000000000;
	sram_mem[128775] = 16'b0000000000000000;
	sram_mem[128776] = 16'b0000000000000000;
	sram_mem[128777] = 16'b0000000000000000;
	sram_mem[128778] = 16'b0000000000000000;
	sram_mem[128779] = 16'b0000000000000000;
	sram_mem[128780] = 16'b0000000000000000;
	sram_mem[128781] = 16'b0000000000000000;
	sram_mem[128782] = 16'b0000000000000000;
	sram_mem[128783] = 16'b0000000000000000;
	sram_mem[128784] = 16'b0000000000000000;
	sram_mem[128785] = 16'b0000000000000000;
	sram_mem[128786] = 16'b0000000000000000;
	sram_mem[128787] = 16'b0000000000000000;
	sram_mem[128788] = 16'b0000000000000000;
	sram_mem[128789] = 16'b0000000000000000;
	sram_mem[128790] = 16'b0000000000000000;
	sram_mem[128791] = 16'b0000000000000000;
	sram_mem[128792] = 16'b0000000000000000;
	sram_mem[128793] = 16'b0000000000000000;
	sram_mem[128794] = 16'b0000000000000000;
	sram_mem[128795] = 16'b0000000000000000;
	sram_mem[128796] = 16'b0000000000000000;
	sram_mem[128797] = 16'b0000000000000000;
	sram_mem[128798] = 16'b0000000000000000;
	sram_mem[128799] = 16'b0000000000000000;
	sram_mem[128800] = 16'b0000000000000000;
	sram_mem[128801] = 16'b0000000000000000;
	sram_mem[128802] = 16'b0000000000000000;
	sram_mem[128803] = 16'b0000000000000000;
	sram_mem[128804] = 16'b0000000000000000;
	sram_mem[128805] = 16'b0000000000000000;
	sram_mem[128806] = 16'b0000000000000000;
	sram_mem[128807] = 16'b0000000000000000;
	sram_mem[128808] = 16'b0000000000000000;
	sram_mem[128809] = 16'b0000000000000000;
	sram_mem[128810] = 16'b0000000000000000;
	sram_mem[128811] = 16'b0000000000000000;
	sram_mem[128812] = 16'b0000000000000000;
	sram_mem[128813] = 16'b0000000000000000;
	sram_mem[128814] = 16'b0000000000000000;
	sram_mem[128815] = 16'b0000000000000000;
	sram_mem[128816] = 16'b0000000000000000;
	sram_mem[128817] = 16'b0000000000000000;
	sram_mem[128818] = 16'b0000000000000000;
	sram_mem[128819] = 16'b0000000000000000;
	sram_mem[128820] = 16'b0000000000000000;
	sram_mem[128821] = 16'b0000000000000000;
	sram_mem[128822] = 16'b0000000000000000;
	sram_mem[128823] = 16'b0000000000000000;
	sram_mem[128824] = 16'b0000000000000000;
	sram_mem[128825] = 16'b0000000000000000;
	sram_mem[128826] = 16'b0000000000000000;
	sram_mem[128827] = 16'b0000000000000000;
	sram_mem[128828] = 16'b0000000000000000;
	sram_mem[128829] = 16'b0000000000000000;
	sram_mem[128830] = 16'b0000000000000000;
	sram_mem[128831] = 16'b0000000000000000;
	sram_mem[128832] = 16'b0000000000000000;
	sram_mem[128833] = 16'b0000000000000000;
	sram_mem[128834] = 16'b0000000000000000;
	sram_mem[128835] = 16'b0000000000000000;
	sram_mem[128836] = 16'b0000000000000000;
	sram_mem[128837] = 16'b0000000000000000;
	sram_mem[128838] = 16'b0000000000000000;
	sram_mem[128839] = 16'b0000000000000000;
	sram_mem[128840] = 16'b0000000000000000;
	sram_mem[128841] = 16'b0000000000000000;
	sram_mem[128842] = 16'b0000000000000000;
	sram_mem[128843] = 16'b0000000000000000;
	sram_mem[128844] = 16'b0000000000000000;
	sram_mem[128845] = 16'b0000000000000000;
	sram_mem[128846] = 16'b0000000000000000;
	sram_mem[128847] = 16'b0000000000000000;
	sram_mem[128848] = 16'b0000000000000000;
	sram_mem[128849] = 16'b0000000000000000;
	sram_mem[128850] = 16'b0000000000000000;
	sram_mem[128851] = 16'b0000000000000000;
	sram_mem[128852] = 16'b0000000000000000;
	sram_mem[128853] = 16'b0000000000000000;
	sram_mem[128854] = 16'b0000000000000000;
	sram_mem[128855] = 16'b0000000000000000;
	sram_mem[128856] = 16'b0000000000000000;
	sram_mem[128857] = 16'b0000000000000000;
	sram_mem[128858] = 16'b0000000000000000;
	sram_mem[128859] = 16'b0000000000000000;
	sram_mem[128860] = 16'b0000000000000000;
	sram_mem[128861] = 16'b0000000000000000;
	sram_mem[128862] = 16'b0000000000000000;
	sram_mem[128863] = 16'b0000000000000000;
	sram_mem[128864] = 16'b0000000000000000;
	sram_mem[128865] = 16'b0000000000000000;
	sram_mem[128866] = 16'b0000000000000000;
	sram_mem[128867] = 16'b0000000000000000;
	sram_mem[128868] = 16'b0000000000000000;
	sram_mem[128869] = 16'b0000000000000000;
	sram_mem[128870] = 16'b0000000000000000;
	sram_mem[128871] = 16'b0000000000000000;
	sram_mem[128872] = 16'b0000000000000000;
	sram_mem[128873] = 16'b0000000000000000;
	sram_mem[128874] = 16'b0000000000000000;
	sram_mem[128875] = 16'b0000000000000000;
	sram_mem[128876] = 16'b0000000000000000;
	sram_mem[128877] = 16'b0000000000000000;
	sram_mem[128878] = 16'b0000000000000000;
	sram_mem[128879] = 16'b0000000000000000;
	sram_mem[128880] = 16'b0000000000000000;
	sram_mem[128881] = 16'b0000000000000000;
	sram_mem[128882] = 16'b0000000000000000;
	sram_mem[128883] = 16'b0000000000000000;
	sram_mem[128884] = 16'b0000000000000000;
	sram_mem[128885] = 16'b0000000000000000;
	sram_mem[128886] = 16'b0000000000000000;
	sram_mem[128887] = 16'b0000000000000000;
	sram_mem[128888] = 16'b0000000000000000;
	sram_mem[128889] = 16'b0000000000000000;
	sram_mem[128890] = 16'b0000000000000000;
	sram_mem[128891] = 16'b0000000000000000;
	sram_mem[128892] = 16'b0000000000000000;
	sram_mem[128893] = 16'b0000000000000000;
	sram_mem[128894] = 16'b0000000000000000;
	sram_mem[128895] = 16'b0000000000000000;
	sram_mem[128896] = 16'b0000000000000000;
	sram_mem[128897] = 16'b0000000000000000;
	sram_mem[128898] = 16'b0000000000000000;
	sram_mem[128899] = 16'b0000000000000000;
	sram_mem[128900] = 16'b0000000000000000;
	sram_mem[128901] = 16'b0000000000000000;
	sram_mem[128902] = 16'b0000000000000000;
	sram_mem[128903] = 16'b0000000000000000;
	sram_mem[128904] = 16'b0000000000000000;
	sram_mem[128905] = 16'b0000000000000000;
	sram_mem[128906] = 16'b0000000000000000;
	sram_mem[128907] = 16'b0000000000000000;
	sram_mem[128908] = 16'b0000000000000000;
	sram_mem[128909] = 16'b0000000000000000;
	sram_mem[128910] = 16'b0000000000000000;
	sram_mem[128911] = 16'b0000000000000000;
	sram_mem[128912] = 16'b0000000000000000;
	sram_mem[128913] = 16'b0000000000000000;
	sram_mem[128914] = 16'b0000000000000000;
	sram_mem[128915] = 16'b0000000000000000;
	sram_mem[128916] = 16'b0000000000000000;
	sram_mem[128917] = 16'b0000000000000000;
	sram_mem[128918] = 16'b0000000000000000;
	sram_mem[128919] = 16'b0000000000000000;
	sram_mem[128920] = 16'b0000000000000000;
	sram_mem[128921] = 16'b0000000000000000;
	sram_mem[128922] = 16'b0000000000000000;
	sram_mem[128923] = 16'b0000000000000000;
	sram_mem[128924] = 16'b0000000000000000;
	sram_mem[128925] = 16'b0000000000000000;
	sram_mem[128926] = 16'b0000000000000000;
	sram_mem[128927] = 16'b0000000000000000;
	sram_mem[128928] = 16'b0000000000000000;
	sram_mem[128929] = 16'b0000000000000000;
	sram_mem[128930] = 16'b0000000000000000;
	sram_mem[128931] = 16'b0000000000000000;
	sram_mem[128932] = 16'b0000000000000000;
	sram_mem[128933] = 16'b0000000000000000;
	sram_mem[128934] = 16'b0000000000000000;
	sram_mem[128935] = 16'b0000000000000000;
	sram_mem[128936] = 16'b0000000000000000;
	sram_mem[128937] = 16'b0000000000000000;
	sram_mem[128938] = 16'b0000000000000000;
	sram_mem[128939] = 16'b0000000000000000;
	sram_mem[128940] = 16'b0000000000000000;
	sram_mem[128941] = 16'b0000000000000000;
	sram_mem[128942] = 16'b0000000000000000;
	sram_mem[128943] = 16'b0000000000000000;
	sram_mem[128944] = 16'b0000000000000000;
	sram_mem[128945] = 16'b0000000000000000;
	sram_mem[128946] = 16'b0000000000000000;
	sram_mem[128947] = 16'b0000000000000000;
	sram_mem[128948] = 16'b0000000000000000;
	sram_mem[128949] = 16'b0000000000000000;
	sram_mem[128950] = 16'b0000000000000000;
	sram_mem[128951] = 16'b0000000000000000;
	sram_mem[128952] = 16'b0000000000000000;
	sram_mem[128953] = 16'b0000000000000000;
	sram_mem[128954] = 16'b0000000000000000;
	sram_mem[128955] = 16'b0000000000000000;
	sram_mem[128956] = 16'b0000000000000000;
	sram_mem[128957] = 16'b0000000000000000;
	sram_mem[128958] = 16'b0000000000000000;
	sram_mem[128959] = 16'b0000000000000000;
	sram_mem[128960] = 16'b0000000000000000;
	sram_mem[128961] = 16'b0000000000000000;
	sram_mem[128962] = 16'b0000000000000000;
	sram_mem[128963] = 16'b0000000000000000;
	sram_mem[128964] = 16'b0000000000000000;
	sram_mem[128965] = 16'b0000000000000000;
	sram_mem[128966] = 16'b0000000000000000;
	sram_mem[128967] = 16'b0000000000000000;
	sram_mem[128968] = 16'b0000000000000000;
	sram_mem[128969] = 16'b0000000000000000;
	sram_mem[128970] = 16'b0000000000000000;
	sram_mem[128971] = 16'b0000000000000000;
	sram_mem[128972] = 16'b0000000000000000;
	sram_mem[128973] = 16'b0000000000000000;
	sram_mem[128974] = 16'b0000000000000000;
	sram_mem[128975] = 16'b0000000000000000;
	sram_mem[128976] = 16'b0000000000000000;
	sram_mem[128977] = 16'b0000000000000000;
	sram_mem[128978] = 16'b0000000000000000;
	sram_mem[128979] = 16'b0000000000000000;
	sram_mem[128980] = 16'b0000000000000000;
	sram_mem[128981] = 16'b0000000000000000;
	sram_mem[128982] = 16'b0000000000000000;
	sram_mem[128983] = 16'b0000000000000000;
	sram_mem[128984] = 16'b0000000000000000;
	sram_mem[128985] = 16'b0000000000000000;
	sram_mem[128986] = 16'b0000000000000000;
	sram_mem[128987] = 16'b0000000000000000;
	sram_mem[128988] = 16'b0000000000000000;
	sram_mem[128989] = 16'b0000000000000000;
	sram_mem[128990] = 16'b0000000000000000;
	sram_mem[128991] = 16'b0000000000000000;
	sram_mem[128992] = 16'b0000000000000000;
	sram_mem[128993] = 16'b0000000000000000;
	sram_mem[128994] = 16'b0000000000000000;
	sram_mem[128995] = 16'b0000000000000000;
	sram_mem[128996] = 16'b0000000000000000;
	sram_mem[128997] = 16'b0000000000000000;
	sram_mem[128998] = 16'b0000000000000000;
	sram_mem[128999] = 16'b0000000000000000;
	sram_mem[129000] = 16'b0000000000000000;
	sram_mem[129001] = 16'b0000000000000000;
	sram_mem[129002] = 16'b0000000000000000;
	sram_mem[129003] = 16'b0000000000000000;
	sram_mem[129004] = 16'b0000000000000000;
	sram_mem[129005] = 16'b0000000000000000;
	sram_mem[129006] = 16'b0000000000000000;
	sram_mem[129007] = 16'b0000000000000000;
	sram_mem[129008] = 16'b0000000000000000;
	sram_mem[129009] = 16'b0000000000000000;
	sram_mem[129010] = 16'b0000000000000000;
	sram_mem[129011] = 16'b0000000000000000;
	sram_mem[129012] = 16'b0000000000000000;
	sram_mem[129013] = 16'b0000000000000000;
	sram_mem[129014] = 16'b0000000000000000;
	sram_mem[129015] = 16'b0000000000000000;
	sram_mem[129016] = 16'b0000000000000000;
	sram_mem[129017] = 16'b0000000000000000;
	sram_mem[129018] = 16'b0000000000000000;
	sram_mem[129019] = 16'b0000000000000000;
	sram_mem[129020] = 16'b0000000000000000;
	sram_mem[129021] = 16'b0000000000000000;
	sram_mem[129022] = 16'b0000000000000000;
	sram_mem[129023] = 16'b0000000000000000;
	sram_mem[129024] = 16'b0000000000000000;
	sram_mem[129025] = 16'b0000000000000000;
	sram_mem[129026] = 16'b0000000000000000;
	sram_mem[129027] = 16'b0000000000000000;
	sram_mem[129028] = 16'b0000000000000000;
	sram_mem[129029] = 16'b0000000000000000;
	sram_mem[129030] = 16'b0000000000000000;
	sram_mem[129031] = 16'b0000000000000000;
	sram_mem[129032] = 16'b0000000000000000;
	sram_mem[129033] = 16'b0000000000000000;
	sram_mem[129034] = 16'b0000000000000000;
	sram_mem[129035] = 16'b0000000000000000;
	sram_mem[129036] = 16'b0000000000000000;
	sram_mem[129037] = 16'b0000000000000000;
	sram_mem[129038] = 16'b0000000000000000;
	sram_mem[129039] = 16'b0000000000000000;
	sram_mem[129040] = 16'b0000000000000000;
	sram_mem[129041] = 16'b0000000000000000;
	sram_mem[129042] = 16'b0000000000000000;
	sram_mem[129043] = 16'b0000000000000000;
	sram_mem[129044] = 16'b0000000000000000;
	sram_mem[129045] = 16'b0000000000000000;
	sram_mem[129046] = 16'b0000000000000000;
	sram_mem[129047] = 16'b0000000000000000;
	sram_mem[129048] = 16'b0000000000000000;
	sram_mem[129049] = 16'b0000000000000000;
	sram_mem[129050] = 16'b0000000000000000;
	sram_mem[129051] = 16'b0000000000000000;
	sram_mem[129052] = 16'b0000000000000000;
	sram_mem[129053] = 16'b0000000000000000;
	sram_mem[129054] = 16'b0000000000000000;
	sram_mem[129055] = 16'b0000000000000000;
	sram_mem[129056] = 16'b0000000000000000;
	sram_mem[129057] = 16'b0000000000000000;
	sram_mem[129058] = 16'b0000000000000000;
	sram_mem[129059] = 16'b0000000000000000;
	sram_mem[129060] = 16'b0000000000000000;
	sram_mem[129061] = 16'b0000000000000000;
	sram_mem[129062] = 16'b0000000000000000;
	sram_mem[129063] = 16'b0000000000000000;
	sram_mem[129064] = 16'b0000000000000000;
	sram_mem[129065] = 16'b0000000000000000;
	sram_mem[129066] = 16'b0000000000000000;
	sram_mem[129067] = 16'b0000000000000000;
	sram_mem[129068] = 16'b0000000000000000;
	sram_mem[129069] = 16'b0000000000000000;
	sram_mem[129070] = 16'b0000000000000000;
	sram_mem[129071] = 16'b0000000000000000;
	sram_mem[129072] = 16'b0000000000000000;
	sram_mem[129073] = 16'b0000000000000000;
	sram_mem[129074] = 16'b0000000000000000;
	sram_mem[129075] = 16'b0000000000000000;
	sram_mem[129076] = 16'b0000000000000000;
	sram_mem[129077] = 16'b0000000000000000;
	sram_mem[129078] = 16'b0000000000000000;
	sram_mem[129079] = 16'b0000000000000000;
	sram_mem[129080] = 16'b0000000000000000;
	sram_mem[129081] = 16'b0000000000000000;
	sram_mem[129082] = 16'b0000000000000000;
	sram_mem[129083] = 16'b0000000000000000;
	sram_mem[129084] = 16'b0000000000000000;
	sram_mem[129085] = 16'b0000000000000000;
	sram_mem[129086] = 16'b0000000000000000;
	sram_mem[129087] = 16'b0000000000000000;
	sram_mem[129088] = 16'b0000000000000000;
	sram_mem[129089] = 16'b0000000000000000;
	sram_mem[129090] = 16'b0000000000000000;
	sram_mem[129091] = 16'b0000000000000000;
	sram_mem[129092] = 16'b0000000000000000;
	sram_mem[129093] = 16'b0000000000000000;
	sram_mem[129094] = 16'b0000000000000000;
	sram_mem[129095] = 16'b0000000000000000;
	sram_mem[129096] = 16'b0000000000000000;
	sram_mem[129097] = 16'b0000000000000000;
	sram_mem[129098] = 16'b0000000000000000;
	sram_mem[129099] = 16'b0000000000000000;
	sram_mem[129100] = 16'b0000000000000000;
	sram_mem[129101] = 16'b0000000000000000;
	sram_mem[129102] = 16'b0000000000000000;
	sram_mem[129103] = 16'b0000000000000000;
	sram_mem[129104] = 16'b0000000000000000;
	sram_mem[129105] = 16'b0000000000000000;
	sram_mem[129106] = 16'b0000000000000000;
	sram_mem[129107] = 16'b0000000000000000;
	sram_mem[129108] = 16'b0000000000000000;
	sram_mem[129109] = 16'b0000000000000000;
	sram_mem[129110] = 16'b0000000000000000;
	sram_mem[129111] = 16'b0000000000000000;
	sram_mem[129112] = 16'b0000000000000000;
	sram_mem[129113] = 16'b0000000000000000;
	sram_mem[129114] = 16'b0000000000000000;
	sram_mem[129115] = 16'b0000000000000000;
	sram_mem[129116] = 16'b0000000000000000;
	sram_mem[129117] = 16'b0000000000000000;
	sram_mem[129118] = 16'b0000000000000000;
	sram_mem[129119] = 16'b0000000000000000;
	sram_mem[129120] = 16'b0000000000000000;
	sram_mem[129121] = 16'b0000000000000000;
	sram_mem[129122] = 16'b0000000000000000;
	sram_mem[129123] = 16'b0000000000000000;
	sram_mem[129124] = 16'b0000000000000000;
	sram_mem[129125] = 16'b0000000000000000;
	sram_mem[129126] = 16'b0000000000000000;
	sram_mem[129127] = 16'b0000000000000000;
	sram_mem[129128] = 16'b0000000000000000;
	sram_mem[129129] = 16'b0000000000000000;
	sram_mem[129130] = 16'b0000000000000000;
	sram_mem[129131] = 16'b0000000000000000;
	sram_mem[129132] = 16'b0000000000000000;
	sram_mem[129133] = 16'b0000000000000000;
	sram_mem[129134] = 16'b0000000000000000;
	sram_mem[129135] = 16'b0000000000000000;
	sram_mem[129136] = 16'b0000000000000000;
	sram_mem[129137] = 16'b0000000000000000;
	sram_mem[129138] = 16'b0000000000000000;
	sram_mem[129139] = 16'b0000000000000000;
	sram_mem[129140] = 16'b0000000000000000;
	sram_mem[129141] = 16'b0000000000000000;
	sram_mem[129142] = 16'b0000000000000000;
	sram_mem[129143] = 16'b0000000000000000;
	sram_mem[129144] = 16'b0000000000000000;
	sram_mem[129145] = 16'b0000000000000000;
	sram_mem[129146] = 16'b0000000000000000;
	sram_mem[129147] = 16'b0000000000000000;
	sram_mem[129148] = 16'b0000000000000000;
	sram_mem[129149] = 16'b0000000000000000;
	sram_mem[129150] = 16'b0000000000000000;
	sram_mem[129151] = 16'b0000000000000000;
	sram_mem[129152] = 16'b0000000000000000;
	sram_mem[129153] = 16'b0000000000000000;
	sram_mem[129154] = 16'b0000000000000000;
	sram_mem[129155] = 16'b0000000000000000;
	sram_mem[129156] = 16'b0000000000000000;
	sram_mem[129157] = 16'b0000000000000000;
	sram_mem[129158] = 16'b0000000000000000;
	sram_mem[129159] = 16'b0000000000000000;
	sram_mem[129160] = 16'b0000000000000000;
	sram_mem[129161] = 16'b0000000000000000;
	sram_mem[129162] = 16'b0000000000000000;
	sram_mem[129163] = 16'b0000000000000000;
	sram_mem[129164] = 16'b0000000000000000;
	sram_mem[129165] = 16'b0000000000000000;
	sram_mem[129166] = 16'b0000000000000000;
	sram_mem[129167] = 16'b0000000000000000;
	sram_mem[129168] = 16'b0000000000000000;
	sram_mem[129169] = 16'b0000000000000000;
	sram_mem[129170] = 16'b0000000000000000;
	sram_mem[129171] = 16'b0000000000000000;
	sram_mem[129172] = 16'b0000000000000000;
	sram_mem[129173] = 16'b0000000000000000;
	sram_mem[129174] = 16'b0000000000000000;
	sram_mem[129175] = 16'b0000000000000000;
	sram_mem[129176] = 16'b0000000000000000;
	sram_mem[129177] = 16'b0000000000000000;
	sram_mem[129178] = 16'b0000000000000000;
	sram_mem[129179] = 16'b0000000000000000;
	sram_mem[129180] = 16'b0000000000000000;
	sram_mem[129181] = 16'b0000000000000000;
	sram_mem[129182] = 16'b0000000000000000;
	sram_mem[129183] = 16'b0000000000000000;
	sram_mem[129184] = 16'b0000000000000000;
	sram_mem[129185] = 16'b0000000000000000;
	sram_mem[129186] = 16'b0000000000000000;
	sram_mem[129187] = 16'b0000000000000000;
	sram_mem[129188] = 16'b0000000000000000;
	sram_mem[129189] = 16'b0000000000000000;
	sram_mem[129190] = 16'b0000000000000000;
	sram_mem[129191] = 16'b0000000000000000;
	sram_mem[129192] = 16'b0000000000000000;
	sram_mem[129193] = 16'b0000000000000000;
	sram_mem[129194] = 16'b0000000000000000;
	sram_mem[129195] = 16'b0000000000000000;
	sram_mem[129196] = 16'b0000000000000000;
	sram_mem[129197] = 16'b0000000000000000;
	sram_mem[129198] = 16'b0000000000000000;
	sram_mem[129199] = 16'b0000000000000000;
	sram_mem[129200] = 16'b0000000000000000;
	sram_mem[129201] = 16'b0000000000000000;
	sram_mem[129202] = 16'b0000000000000000;
	sram_mem[129203] = 16'b0000000000000000;
	sram_mem[129204] = 16'b0000000000000000;
	sram_mem[129205] = 16'b0000000000000000;
	sram_mem[129206] = 16'b0000000000000000;
	sram_mem[129207] = 16'b0000000000000000;
	sram_mem[129208] = 16'b0000000000000000;
	sram_mem[129209] = 16'b0000000000000000;
	sram_mem[129210] = 16'b0000000000000000;
	sram_mem[129211] = 16'b0000000000000000;
	sram_mem[129212] = 16'b0000000000000000;
	sram_mem[129213] = 16'b0000000000000000;
	sram_mem[129214] = 16'b0000000000000000;
	sram_mem[129215] = 16'b0000000000000000;
	sram_mem[129216] = 16'b0000000000000000;
	sram_mem[129217] = 16'b0000000000000000;
	sram_mem[129218] = 16'b0000000000000000;
	sram_mem[129219] = 16'b0000000000000000;
	sram_mem[129220] = 16'b0000000000000000;
	sram_mem[129221] = 16'b0000000000000000;
	sram_mem[129222] = 16'b0000000000000000;
	sram_mem[129223] = 16'b0000000000000000;
	sram_mem[129224] = 16'b0000000000000000;
	sram_mem[129225] = 16'b0000000000000000;
	sram_mem[129226] = 16'b0000000000000000;
	sram_mem[129227] = 16'b0000000000000000;
	sram_mem[129228] = 16'b0000000000000000;
	sram_mem[129229] = 16'b0000000000000000;
	sram_mem[129230] = 16'b0000000000000000;
	sram_mem[129231] = 16'b0000000000000000;
	sram_mem[129232] = 16'b0000000000000000;
	sram_mem[129233] = 16'b0000000000000000;
	sram_mem[129234] = 16'b0000000000000000;
	sram_mem[129235] = 16'b0000000000000000;
	sram_mem[129236] = 16'b0000000000000000;
	sram_mem[129237] = 16'b0000000000000000;
	sram_mem[129238] = 16'b0000000000000000;
	sram_mem[129239] = 16'b0000000000000000;
	sram_mem[129240] = 16'b0000000000000000;
	sram_mem[129241] = 16'b0000000000000000;
	sram_mem[129242] = 16'b0000000000000000;
	sram_mem[129243] = 16'b0000000000000000;
	sram_mem[129244] = 16'b0000000000000000;
	sram_mem[129245] = 16'b0000000000000000;
	sram_mem[129246] = 16'b0000000000000000;
	sram_mem[129247] = 16'b0000000000000000;
	sram_mem[129248] = 16'b0000000000000000;
	sram_mem[129249] = 16'b0000000000000000;
	sram_mem[129250] = 16'b0000000000000000;
	sram_mem[129251] = 16'b0000000000000000;
	sram_mem[129252] = 16'b0000000000000000;
	sram_mem[129253] = 16'b0000000000000000;
	sram_mem[129254] = 16'b0000000000000000;
	sram_mem[129255] = 16'b0000000000000000;
	sram_mem[129256] = 16'b0000000000000000;
	sram_mem[129257] = 16'b0000000000000000;
	sram_mem[129258] = 16'b0000000000000000;
	sram_mem[129259] = 16'b0000000000000000;
	sram_mem[129260] = 16'b0000000000000000;
	sram_mem[129261] = 16'b0000000000000000;
	sram_mem[129262] = 16'b0000000000000000;
	sram_mem[129263] = 16'b0000000000000000;
	sram_mem[129264] = 16'b0000000000000000;
	sram_mem[129265] = 16'b0000000000000000;
	sram_mem[129266] = 16'b0000000000000000;
	sram_mem[129267] = 16'b0000000000000000;
	sram_mem[129268] = 16'b0000000000000000;
	sram_mem[129269] = 16'b0000000000000000;
	sram_mem[129270] = 16'b0000000000000000;
	sram_mem[129271] = 16'b0000000000000000;
	sram_mem[129272] = 16'b0000000000000000;
	sram_mem[129273] = 16'b0000000000000000;
	sram_mem[129274] = 16'b0000000000000000;
	sram_mem[129275] = 16'b0000000000000000;
	sram_mem[129276] = 16'b0000000000000000;
	sram_mem[129277] = 16'b0000000000000000;
	sram_mem[129278] = 16'b0000000000000000;
	sram_mem[129279] = 16'b0000000000000000;
	sram_mem[129280] = 16'b0000000000000000;
	sram_mem[129281] = 16'b0000000000000000;
	sram_mem[129282] = 16'b0000000000000000;
	sram_mem[129283] = 16'b0000000000000000;
	sram_mem[129284] = 16'b0000000000000000;
	sram_mem[129285] = 16'b0000000000000000;
	sram_mem[129286] = 16'b0000000000000000;
	sram_mem[129287] = 16'b0000000000000000;
	sram_mem[129288] = 16'b0000000000000000;
	sram_mem[129289] = 16'b0000000000000000;
	sram_mem[129290] = 16'b0000000000000000;
	sram_mem[129291] = 16'b0000000000000000;
	sram_mem[129292] = 16'b0000000000000000;
	sram_mem[129293] = 16'b0000000000000000;
	sram_mem[129294] = 16'b0000000000000000;
	sram_mem[129295] = 16'b0000000000000000;
	sram_mem[129296] = 16'b0000000000000000;
	sram_mem[129297] = 16'b0000000000000000;
	sram_mem[129298] = 16'b0000000000000000;
	sram_mem[129299] = 16'b0000000000000000;
	sram_mem[129300] = 16'b0000000000000000;
	sram_mem[129301] = 16'b0000000000000000;
	sram_mem[129302] = 16'b0000000000000000;
	sram_mem[129303] = 16'b0000000000000000;
	sram_mem[129304] = 16'b0000000000000000;
	sram_mem[129305] = 16'b0000000000000000;
	sram_mem[129306] = 16'b0000000000000000;
	sram_mem[129307] = 16'b0000000000000000;
	sram_mem[129308] = 16'b0000000000000000;
	sram_mem[129309] = 16'b0000000000000000;
	sram_mem[129310] = 16'b0000000000000000;
	sram_mem[129311] = 16'b0000000000000000;
	sram_mem[129312] = 16'b0000000000000000;
	sram_mem[129313] = 16'b0000000000000000;
	sram_mem[129314] = 16'b0000000000000000;
	sram_mem[129315] = 16'b0000000000000000;
	sram_mem[129316] = 16'b0000000000000000;
	sram_mem[129317] = 16'b0000000000000000;
	sram_mem[129318] = 16'b0000000000000000;
	sram_mem[129319] = 16'b0000000000000000;
	sram_mem[129320] = 16'b0000000000000000;
	sram_mem[129321] = 16'b0000000000000000;
	sram_mem[129322] = 16'b0000000000000000;
	sram_mem[129323] = 16'b0000000000000000;
	sram_mem[129324] = 16'b0000000000000000;
	sram_mem[129325] = 16'b0000000000000000;
	sram_mem[129326] = 16'b0000000000000000;
	sram_mem[129327] = 16'b0000000000000000;
	sram_mem[129328] = 16'b0000000000000000;
	sram_mem[129329] = 16'b0000000000000000;
	sram_mem[129330] = 16'b0000000000000000;
	sram_mem[129331] = 16'b0000000000000000;
	sram_mem[129332] = 16'b0000000000000000;
	sram_mem[129333] = 16'b0000000000000000;
	sram_mem[129334] = 16'b0000000000000000;
	sram_mem[129335] = 16'b0000000000000000;
	sram_mem[129336] = 16'b0000000000000000;
	sram_mem[129337] = 16'b0000000000000000;
	sram_mem[129338] = 16'b0000000000000000;
	sram_mem[129339] = 16'b0000000000000000;
	sram_mem[129340] = 16'b0000000000000000;
	sram_mem[129341] = 16'b0000000000000000;
	sram_mem[129342] = 16'b0000000000000000;
	sram_mem[129343] = 16'b0000000000000000;
	sram_mem[129344] = 16'b0000000000000000;
	sram_mem[129345] = 16'b0000000000000000;
	sram_mem[129346] = 16'b0000000000000000;
	sram_mem[129347] = 16'b0000000000000000;
	sram_mem[129348] = 16'b0000000000000000;
	sram_mem[129349] = 16'b0000000000000000;
	sram_mem[129350] = 16'b0000000000000000;
	sram_mem[129351] = 16'b0000000000000000;
	sram_mem[129352] = 16'b0000000000000000;
	sram_mem[129353] = 16'b0000000000000000;
	sram_mem[129354] = 16'b0000000000000000;
	sram_mem[129355] = 16'b0000000000000000;
	sram_mem[129356] = 16'b0000000000000000;
	sram_mem[129357] = 16'b0000000000000000;
	sram_mem[129358] = 16'b0000000000000000;
	sram_mem[129359] = 16'b0000000000000000;
	sram_mem[129360] = 16'b0000000000000000;
	sram_mem[129361] = 16'b0000000000000000;
	sram_mem[129362] = 16'b0000000000000000;
	sram_mem[129363] = 16'b0000000000000000;
	sram_mem[129364] = 16'b0000000000000000;
	sram_mem[129365] = 16'b0000000000000000;
	sram_mem[129366] = 16'b0000000000000000;
	sram_mem[129367] = 16'b0000000000000000;
	sram_mem[129368] = 16'b0000000000000000;
	sram_mem[129369] = 16'b0000000000000000;
	sram_mem[129370] = 16'b0000000000000000;
	sram_mem[129371] = 16'b0000000000000000;
	sram_mem[129372] = 16'b0000000000000000;
	sram_mem[129373] = 16'b0000000000000000;
	sram_mem[129374] = 16'b0000000000000000;
	sram_mem[129375] = 16'b0000000000000000;
	sram_mem[129376] = 16'b0000000000000000;
	sram_mem[129377] = 16'b0000000000000000;
	sram_mem[129378] = 16'b0000000000000000;
	sram_mem[129379] = 16'b0000000000000000;
	sram_mem[129380] = 16'b0000000000000000;
	sram_mem[129381] = 16'b0000000000000000;
	sram_mem[129382] = 16'b0000000000000000;
	sram_mem[129383] = 16'b0000000000000000;
	sram_mem[129384] = 16'b0000000000000000;
	sram_mem[129385] = 16'b0000000000000000;
	sram_mem[129386] = 16'b0000000000000000;
	sram_mem[129387] = 16'b0000000000000000;
	sram_mem[129388] = 16'b0000000000000000;
	sram_mem[129389] = 16'b0000000000000000;
	sram_mem[129390] = 16'b0000000000000000;
	sram_mem[129391] = 16'b0000000000000000;
	sram_mem[129392] = 16'b0000000000000000;
	sram_mem[129393] = 16'b0000000000000000;
	sram_mem[129394] = 16'b0000000000000000;
	sram_mem[129395] = 16'b0000000000000000;
	sram_mem[129396] = 16'b0000000000000000;
	sram_mem[129397] = 16'b0000000000000000;
	sram_mem[129398] = 16'b0000000000000000;
	sram_mem[129399] = 16'b0000000000000000;
	sram_mem[129400] = 16'b0000000000000000;
	sram_mem[129401] = 16'b0000000000000000;
	sram_mem[129402] = 16'b0000000000000000;
	sram_mem[129403] = 16'b0000000000000000;
	sram_mem[129404] = 16'b0000000000000000;
	sram_mem[129405] = 16'b0000000000000000;
	sram_mem[129406] = 16'b0000000000000000;
	sram_mem[129407] = 16'b0000000000000000;
	sram_mem[129408] = 16'b0000000000000000;
	sram_mem[129409] = 16'b0000000000000000;
	sram_mem[129410] = 16'b0000000000000000;
	sram_mem[129411] = 16'b0000000000000000;
	sram_mem[129412] = 16'b0000000000000000;
	sram_mem[129413] = 16'b0000000000000000;
	sram_mem[129414] = 16'b0000000000000000;
	sram_mem[129415] = 16'b0000000000000000;
	sram_mem[129416] = 16'b0000000000000000;
	sram_mem[129417] = 16'b0000000000000000;
	sram_mem[129418] = 16'b0000000000000000;
	sram_mem[129419] = 16'b0000000000000000;
	sram_mem[129420] = 16'b0000000000000000;
	sram_mem[129421] = 16'b0000000000000000;
	sram_mem[129422] = 16'b0000000000000000;
	sram_mem[129423] = 16'b0000000000000000;
	sram_mem[129424] = 16'b0000000000000000;
	sram_mem[129425] = 16'b0000000000000000;
	sram_mem[129426] = 16'b0000000000000000;
	sram_mem[129427] = 16'b0000000000000000;
	sram_mem[129428] = 16'b0000000000000000;
	sram_mem[129429] = 16'b0000000000000000;
	sram_mem[129430] = 16'b0000000000000000;
	sram_mem[129431] = 16'b0000000000000000;
	sram_mem[129432] = 16'b0000000000000000;
	sram_mem[129433] = 16'b0000000000000000;
	sram_mem[129434] = 16'b0000000000000000;
	sram_mem[129435] = 16'b0000000000000000;
	sram_mem[129436] = 16'b0000000000000000;
	sram_mem[129437] = 16'b0000000000000000;
	sram_mem[129438] = 16'b0000000000000000;
	sram_mem[129439] = 16'b0000000000000000;
	sram_mem[129440] = 16'b0000000000000000;
	sram_mem[129441] = 16'b0000000000000000;
	sram_mem[129442] = 16'b0000000000000000;
	sram_mem[129443] = 16'b0000000000000000;
	sram_mem[129444] = 16'b0000000000000000;
	sram_mem[129445] = 16'b0000000000000000;
	sram_mem[129446] = 16'b0000000000000000;
	sram_mem[129447] = 16'b0000000000000000;
	sram_mem[129448] = 16'b0000000000000000;
	sram_mem[129449] = 16'b0000000000000000;
	sram_mem[129450] = 16'b0000000000000000;
	sram_mem[129451] = 16'b0000000000000000;
	sram_mem[129452] = 16'b0000000000000000;
	sram_mem[129453] = 16'b0000000000000000;
	sram_mem[129454] = 16'b0000000000000000;
	sram_mem[129455] = 16'b0000000000000000;
	sram_mem[129456] = 16'b0000000000000000;
	sram_mem[129457] = 16'b0000000000000000;
	sram_mem[129458] = 16'b0000000000000000;
	sram_mem[129459] = 16'b0000000000000000;
	sram_mem[129460] = 16'b0000000000000000;
	sram_mem[129461] = 16'b0000000000000000;
	sram_mem[129462] = 16'b0000000000000000;
	sram_mem[129463] = 16'b0000000000000000;
	sram_mem[129464] = 16'b0000000000000000;
	sram_mem[129465] = 16'b0000000000000000;
	sram_mem[129466] = 16'b0000000000000000;
	sram_mem[129467] = 16'b0000000000000000;
	sram_mem[129468] = 16'b0000000000000000;
	sram_mem[129469] = 16'b0000000000000000;
	sram_mem[129470] = 16'b0000000000000000;
	sram_mem[129471] = 16'b0000000000000000;
	sram_mem[129472] = 16'b0000000000000000;
	sram_mem[129473] = 16'b0000000000000000;
	sram_mem[129474] = 16'b0000000000000000;
	sram_mem[129475] = 16'b0000000000000000;
	sram_mem[129476] = 16'b0000000000000000;
	sram_mem[129477] = 16'b0000000000000000;
	sram_mem[129478] = 16'b0000000000000000;
	sram_mem[129479] = 16'b0000000000000000;
	sram_mem[129480] = 16'b0000000000000000;
	sram_mem[129481] = 16'b0000000000000000;
	sram_mem[129482] = 16'b0000000000000000;
	sram_mem[129483] = 16'b0000000000000000;
	sram_mem[129484] = 16'b0000000000000000;
	sram_mem[129485] = 16'b0000000000000000;
	sram_mem[129486] = 16'b0000000000000000;
	sram_mem[129487] = 16'b0000000000000000;
	sram_mem[129488] = 16'b0000000000000000;
	sram_mem[129489] = 16'b0000000000000000;
	sram_mem[129490] = 16'b0000000000000000;
	sram_mem[129491] = 16'b0000000000000000;
	sram_mem[129492] = 16'b0000000000000000;
	sram_mem[129493] = 16'b0000000000000000;
	sram_mem[129494] = 16'b0000000000000000;
	sram_mem[129495] = 16'b0000000000000000;
	sram_mem[129496] = 16'b0000000000000000;
	sram_mem[129497] = 16'b0000000000000000;
	sram_mem[129498] = 16'b0000000000000000;
	sram_mem[129499] = 16'b0000000000000000;
	sram_mem[129500] = 16'b0000000000000000;
	sram_mem[129501] = 16'b0000000000000000;
	sram_mem[129502] = 16'b0000000000000000;
	sram_mem[129503] = 16'b0000000000000000;
	sram_mem[129504] = 16'b0000000000000000;
	sram_mem[129505] = 16'b0000000000000000;
	sram_mem[129506] = 16'b0000000000000000;
	sram_mem[129507] = 16'b0000000000000000;
	sram_mem[129508] = 16'b0000000000000000;
	sram_mem[129509] = 16'b0000000000000000;
	sram_mem[129510] = 16'b0000000000000000;
	sram_mem[129511] = 16'b0000000000000000;
	sram_mem[129512] = 16'b0000000000000000;
	sram_mem[129513] = 16'b0000000000000000;
	sram_mem[129514] = 16'b0000000000000000;
	sram_mem[129515] = 16'b0000000000000000;
	sram_mem[129516] = 16'b0000000000000000;
	sram_mem[129517] = 16'b0000000000000000;
	sram_mem[129518] = 16'b0000000000000000;
	sram_mem[129519] = 16'b0000000000000000;
	sram_mem[129520] = 16'b0000000000000000;
	sram_mem[129521] = 16'b0000000000000000;
	sram_mem[129522] = 16'b0000000000000000;
	sram_mem[129523] = 16'b0000000000000000;
	sram_mem[129524] = 16'b0000000000000000;
	sram_mem[129525] = 16'b0000000000000000;
	sram_mem[129526] = 16'b0000000000000000;
	sram_mem[129527] = 16'b0000000000000000;
	sram_mem[129528] = 16'b0000000000000000;
	sram_mem[129529] = 16'b0000000000000000;
	sram_mem[129530] = 16'b0000000000000000;
	sram_mem[129531] = 16'b0000000000000000;
	sram_mem[129532] = 16'b0000000000000000;
	sram_mem[129533] = 16'b0000000000000000;
	sram_mem[129534] = 16'b0000000000000000;
	sram_mem[129535] = 16'b0000000000000000;
	sram_mem[129536] = 16'b0000000000000000;
	sram_mem[129537] = 16'b0000000000000000;
	sram_mem[129538] = 16'b0000000000000000;
	sram_mem[129539] = 16'b0000000000000000;
	sram_mem[129540] = 16'b0000000000000000;
	sram_mem[129541] = 16'b0000000000000000;
	sram_mem[129542] = 16'b0000000000000000;
	sram_mem[129543] = 16'b0000000000000000;
	sram_mem[129544] = 16'b0000000000000000;
	sram_mem[129545] = 16'b0000000000000000;
	sram_mem[129546] = 16'b0000000000000000;
	sram_mem[129547] = 16'b0000000000000000;
	sram_mem[129548] = 16'b0000000000000000;
	sram_mem[129549] = 16'b0000000000000000;
	sram_mem[129550] = 16'b0000000000000000;
	sram_mem[129551] = 16'b0000000000000000;
	sram_mem[129552] = 16'b0000000000000000;
	sram_mem[129553] = 16'b0000000000000000;
	sram_mem[129554] = 16'b0000000000000000;
	sram_mem[129555] = 16'b0000000000000000;
	sram_mem[129556] = 16'b0000000000000000;
	sram_mem[129557] = 16'b0000000000000000;
	sram_mem[129558] = 16'b0000000000000000;
	sram_mem[129559] = 16'b0000000000000000;
	sram_mem[129560] = 16'b0000000000000000;
	sram_mem[129561] = 16'b0000000000000000;
	sram_mem[129562] = 16'b0000000000000000;
	sram_mem[129563] = 16'b0000000000000000;
	sram_mem[129564] = 16'b0000000000000000;
	sram_mem[129565] = 16'b0000000000000000;
	sram_mem[129566] = 16'b0000000000000000;
	sram_mem[129567] = 16'b0000000000000000;
	sram_mem[129568] = 16'b0000000000000000;
	sram_mem[129569] = 16'b0000000000000000;
	sram_mem[129570] = 16'b0000000000000000;
	sram_mem[129571] = 16'b0000000000000000;
	sram_mem[129572] = 16'b0000000000000000;
	sram_mem[129573] = 16'b0000000000000000;
	sram_mem[129574] = 16'b0000000000000000;
	sram_mem[129575] = 16'b0000000000000000;
	sram_mem[129576] = 16'b0000000000000000;
	sram_mem[129577] = 16'b0000000000000000;
	sram_mem[129578] = 16'b0000000000000000;
	sram_mem[129579] = 16'b0000000000000000;
	sram_mem[129580] = 16'b0000000000000000;
	sram_mem[129581] = 16'b0000000000000000;
	sram_mem[129582] = 16'b0000000000000000;
	sram_mem[129583] = 16'b0000000000000000;
	sram_mem[129584] = 16'b0000000000000000;
	sram_mem[129585] = 16'b0000000000000000;
	sram_mem[129586] = 16'b0000000000000000;
	sram_mem[129587] = 16'b0000000000000000;
	sram_mem[129588] = 16'b0000000000000000;
	sram_mem[129589] = 16'b0000000000000000;
	sram_mem[129590] = 16'b0000000000000000;
	sram_mem[129591] = 16'b0000000000000000;
	sram_mem[129592] = 16'b0000000000000000;
	sram_mem[129593] = 16'b0000000000000000;
	sram_mem[129594] = 16'b0000000000000000;
	sram_mem[129595] = 16'b0000000000000000;
	sram_mem[129596] = 16'b0000000000000000;
	sram_mem[129597] = 16'b0000000000000000;
	sram_mem[129598] = 16'b0000000000000000;
	sram_mem[129599] = 16'b0000000000000000;
	sram_mem[129600] = 16'b0000000000000000;
	sram_mem[129601] = 16'b0000000000000000;
	sram_mem[129602] = 16'b0000000000000000;
	sram_mem[129603] = 16'b0000000000000000;
	sram_mem[129604] = 16'b0000000000000000;
	sram_mem[129605] = 16'b0000000000000000;
	sram_mem[129606] = 16'b0000000000000000;
	sram_mem[129607] = 16'b0000000000000000;
	sram_mem[129608] = 16'b0000000000000000;
	sram_mem[129609] = 16'b0000000000000000;
	sram_mem[129610] = 16'b0000000000000000;
	sram_mem[129611] = 16'b0000000000000000;
	sram_mem[129612] = 16'b0000000000000000;
	sram_mem[129613] = 16'b0000000000000000;
	sram_mem[129614] = 16'b0000000000000000;
	sram_mem[129615] = 16'b0000000000000000;
	sram_mem[129616] = 16'b0000000000000000;
	sram_mem[129617] = 16'b0000000000000000;
	sram_mem[129618] = 16'b0000000000000000;
	sram_mem[129619] = 16'b0000000000000000;
	sram_mem[129620] = 16'b0000000000000000;
	sram_mem[129621] = 16'b0000000000000000;
	sram_mem[129622] = 16'b0000000000000000;
	sram_mem[129623] = 16'b0000000000000000;
	sram_mem[129624] = 16'b0000000000000000;
	sram_mem[129625] = 16'b0000000000000000;
	sram_mem[129626] = 16'b0000000000000000;
	sram_mem[129627] = 16'b0000000000000000;
	sram_mem[129628] = 16'b0000000000000000;
	sram_mem[129629] = 16'b0000000000000000;
	sram_mem[129630] = 16'b0000000000000000;
	sram_mem[129631] = 16'b0000000000000000;
	sram_mem[129632] = 16'b0000000000000000;
	sram_mem[129633] = 16'b0000000000000000;
	sram_mem[129634] = 16'b0000000000000000;
	sram_mem[129635] = 16'b0000000000000000;
	sram_mem[129636] = 16'b0000000000000000;
	sram_mem[129637] = 16'b0000000000000000;
	sram_mem[129638] = 16'b0000000000000000;
	sram_mem[129639] = 16'b0000000000000000;
	sram_mem[129640] = 16'b0000000000000000;
	sram_mem[129641] = 16'b0000000000000000;
	sram_mem[129642] = 16'b0000000000000000;
	sram_mem[129643] = 16'b0000000000000000;
	sram_mem[129644] = 16'b0000000000000000;
	sram_mem[129645] = 16'b0000000000000000;
	sram_mem[129646] = 16'b0000000000000000;
	sram_mem[129647] = 16'b0000000000000000;
	sram_mem[129648] = 16'b0000000000000000;
	sram_mem[129649] = 16'b0000000000000000;
	sram_mem[129650] = 16'b0000000000000000;
	sram_mem[129651] = 16'b0000000000000000;
	sram_mem[129652] = 16'b0000000000000000;
	sram_mem[129653] = 16'b0000000000000000;
	sram_mem[129654] = 16'b0000000000000000;
	sram_mem[129655] = 16'b0000000000000000;
	sram_mem[129656] = 16'b0000000000000000;
	sram_mem[129657] = 16'b0000000000000000;
	sram_mem[129658] = 16'b0000000000000000;
	sram_mem[129659] = 16'b0000000000000000;
	sram_mem[129660] = 16'b0000000000000000;
	sram_mem[129661] = 16'b0000000000000000;
	sram_mem[129662] = 16'b0000000000000000;
	sram_mem[129663] = 16'b0000000000000000;
	sram_mem[129664] = 16'b0000000000000000;
	sram_mem[129665] = 16'b0000000000000000;
	sram_mem[129666] = 16'b0000000000000000;
	sram_mem[129667] = 16'b0000000000000000;
	sram_mem[129668] = 16'b0000000000000000;
	sram_mem[129669] = 16'b0000000000000000;
	sram_mem[129670] = 16'b0000000000000000;
	sram_mem[129671] = 16'b0000000000000000;
	sram_mem[129672] = 16'b0000000000000000;
	sram_mem[129673] = 16'b0000000000000000;
	sram_mem[129674] = 16'b0000000000000000;
	sram_mem[129675] = 16'b0000000000000000;
	sram_mem[129676] = 16'b0000000000000000;
	sram_mem[129677] = 16'b0000000000000000;
	sram_mem[129678] = 16'b0000000000000000;
	sram_mem[129679] = 16'b0000000000000000;
	sram_mem[129680] = 16'b0000000000000000;
	sram_mem[129681] = 16'b0000000000000000;
	sram_mem[129682] = 16'b0000000000000000;
	sram_mem[129683] = 16'b0000000000000000;
	sram_mem[129684] = 16'b0000000000000000;
	sram_mem[129685] = 16'b0000000000000000;
	sram_mem[129686] = 16'b0000000000000000;
	sram_mem[129687] = 16'b0000000000000000;
	sram_mem[129688] = 16'b0000000000000000;
	sram_mem[129689] = 16'b0000000000000000;
	sram_mem[129690] = 16'b0000000000000000;
	sram_mem[129691] = 16'b0000000000000000;
	sram_mem[129692] = 16'b0000000000000000;
	sram_mem[129693] = 16'b0000000000000000;
	sram_mem[129694] = 16'b0000000000000000;
	sram_mem[129695] = 16'b0000000000000000;
	sram_mem[129696] = 16'b0000000000000000;
	sram_mem[129697] = 16'b0000000000000000;
	sram_mem[129698] = 16'b0000000000000000;
	sram_mem[129699] = 16'b0000000000000000;
	sram_mem[129700] = 16'b0000000000000000;
	sram_mem[129701] = 16'b0000000000000000;
	sram_mem[129702] = 16'b0000000000000000;
	sram_mem[129703] = 16'b0000000000000000;
	sram_mem[129704] = 16'b0000000000000000;
	sram_mem[129705] = 16'b0000000000000000;
	sram_mem[129706] = 16'b0000000000000000;
	sram_mem[129707] = 16'b0000000000000000;
	sram_mem[129708] = 16'b0000000000000000;
	sram_mem[129709] = 16'b0000000000000000;
	sram_mem[129710] = 16'b0000000000000000;
	sram_mem[129711] = 16'b0000000000000000;
	sram_mem[129712] = 16'b0000000000000000;
	sram_mem[129713] = 16'b0000000000000000;
	sram_mem[129714] = 16'b0000000000000000;
	sram_mem[129715] = 16'b0000000000000000;
	sram_mem[129716] = 16'b0000000000000000;
	sram_mem[129717] = 16'b0000000000000000;
	sram_mem[129718] = 16'b0000000000000000;
	sram_mem[129719] = 16'b0000000000000000;
	sram_mem[129720] = 16'b0000000000000000;
	sram_mem[129721] = 16'b0000000000000000;
	sram_mem[129722] = 16'b0000000000000000;
	sram_mem[129723] = 16'b0000000000000000;
	sram_mem[129724] = 16'b0000000000000000;
	sram_mem[129725] = 16'b0000000000000000;
	sram_mem[129726] = 16'b0000000000000000;
	sram_mem[129727] = 16'b0000000000000000;
	sram_mem[129728] = 16'b0000000000000000;
	sram_mem[129729] = 16'b0000000000000000;
	sram_mem[129730] = 16'b0000000000000000;
	sram_mem[129731] = 16'b0000000000000000;
	sram_mem[129732] = 16'b0000000000000000;
	sram_mem[129733] = 16'b0000000000000000;
	sram_mem[129734] = 16'b0000000000000000;
	sram_mem[129735] = 16'b0000000000000000;
	sram_mem[129736] = 16'b0000000000000000;
	sram_mem[129737] = 16'b0000000000000000;
	sram_mem[129738] = 16'b0000000000000000;
	sram_mem[129739] = 16'b0000000000000000;
	sram_mem[129740] = 16'b0000000000000000;
	sram_mem[129741] = 16'b0000000000000000;
	sram_mem[129742] = 16'b0000000000000000;
	sram_mem[129743] = 16'b0000000000000000;
	sram_mem[129744] = 16'b0000000000000000;
	sram_mem[129745] = 16'b0000000000000000;
	sram_mem[129746] = 16'b0000000000000000;
	sram_mem[129747] = 16'b0000000000000000;
	sram_mem[129748] = 16'b0000000000000000;
	sram_mem[129749] = 16'b0000000000000000;
	sram_mem[129750] = 16'b0000000000000000;
	sram_mem[129751] = 16'b0000000000000000;
	sram_mem[129752] = 16'b0000000000000000;
	sram_mem[129753] = 16'b0000000000000000;
	sram_mem[129754] = 16'b0000000000000000;
	sram_mem[129755] = 16'b0000000000000000;
	sram_mem[129756] = 16'b0000000000000000;
	sram_mem[129757] = 16'b0000000000000000;
	sram_mem[129758] = 16'b0000000000000000;
	sram_mem[129759] = 16'b0000000000000000;
	sram_mem[129760] = 16'b0000000000000000;
	sram_mem[129761] = 16'b0000000000000000;
	sram_mem[129762] = 16'b0000000000000000;
	sram_mem[129763] = 16'b0000000000000000;
	sram_mem[129764] = 16'b0000000000000000;
	sram_mem[129765] = 16'b0000000000000000;
	sram_mem[129766] = 16'b0000000000000000;
	sram_mem[129767] = 16'b0000000000000000;
	sram_mem[129768] = 16'b0000000000000000;
	sram_mem[129769] = 16'b0000000000000000;
	sram_mem[129770] = 16'b0000000000000000;
	sram_mem[129771] = 16'b0000000000000000;
	sram_mem[129772] = 16'b0000000000000000;
	sram_mem[129773] = 16'b0000000000000000;
	sram_mem[129774] = 16'b0000000000000000;
	sram_mem[129775] = 16'b0000000000000000;
	sram_mem[129776] = 16'b0000000000000000;
	sram_mem[129777] = 16'b0000000000000000;
	sram_mem[129778] = 16'b0000000000000000;
	sram_mem[129779] = 16'b0000000000000000;
	sram_mem[129780] = 16'b0000000000000000;
	sram_mem[129781] = 16'b0000000000000000;
	sram_mem[129782] = 16'b0000000000000000;
	sram_mem[129783] = 16'b0000000000000000;
	sram_mem[129784] = 16'b0000000000000000;
	sram_mem[129785] = 16'b0000000000000000;
	sram_mem[129786] = 16'b0000000000000000;
	sram_mem[129787] = 16'b0000000000000000;
	sram_mem[129788] = 16'b0000000000000000;
	sram_mem[129789] = 16'b0000000000000000;
	sram_mem[129790] = 16'b0000000000000000;
	sram_mem[129791] = 16'b0000000000000000;
	sram_mem[129792] = 16'b0000000000000000;
	sram_mem[129793] = 16'b0000000000000000;
	sram_mem[129794] = 16'b0000000000000000;
	sram_mem[129795] = 16'b0000000000000000;
	sram_mem[129796] = 16'b0000000000000000;
	sram_mem[129797] = 16'b0000000000000000;
	sram_mem[129798] = 16'b0000000000000000;
	sram_mem[129799] = 16'b0000000000000000;
	sram_mem[129800] = 16'b0000000000000000;
	sram_mem[129801] = 16'b0000000000000000;
	sram_mem[129802] = 16'b0000000000000000;
	sram_mem[129803] = 16'b0000000000000000;
	sram_mem[129804] = 16'b0000000000000000;
	sram_mem[129805] = 16'b0000000000000000;
	sram_mem[129806] = 16'b0000000000000000;
	sram_mem[129807] = 16'b0000000000000000;
	sram_mem[129808] = 16'b0000000000000000;
	sram_mem[129809] = 16'b0000000000000000;
	sram_mem[129810] = 16'b0000000000000000;
	sram_mem[129811] = 16'b0000000000000000;
	sram_mem[129812] = 16'b0000000000000000;
	sram_mem[129813] = 16'b0000000000000000;
	sram_mem[129814] = 16'b0000000000000000;
	sram_mem[129815] = 16'b0000000000000000;
	sram_mem[129816] = 16'b0000000000000000;
	sram_mem[129817] = 16'b0000000000000000;
	sram_mem[129818] = 16'b0000000000000000;
	sram_mem[129819] = 16'b0000000000000000;
	sram_mem[129820] = 16'b0000000000000000;
	sram_mem[129821] = 16'b0000000000000000;
	sram_mem[129822] = 16'b0000000000000000;
	sram_mem[129823] = 16'b0000000000000000;
	sram_mem[129824] = 16'b0000000000000000;
	sram_mem[129825] = 16'b0000000000000000;
	sram_mem[129826] = 16'b0000000000000000;
	sram_mem[129827] = 16'b0000000000000000;
	sram_mem[129828] = 16'b0000000000000000;
	sram_mem[129829] = 16'b0000000000000000;
	sram_mem[129830] = 16'b0000000000000000;
	sram_mem[129831] = 16'b0000000000000000;
	sram_mem[129832] = 16'b0000000000000000;
	sram_mem[129833] = 16'b0000000000000000;
	sram_mem[129834] = 16'b0000000000000000;
	sram_mem[129835] = 16'b0000000000000000;
	sram_mem[129836] = 16'b0000000000000000;
	sram_mem[129837] = 16'b0000000000000000;
	sram_mem[129838] = 16'b0000000000000000;
	sram_mem[129839] = 16'b0000000000000000;
	sram_mem[129840] = 16'b0000000000000000;
	sram_mem[129841] = 16'b0000000000000000;
	sram_mem[129842] = 16'b0000000000000000;
	sram_mem[129843] = 16'b0000000000000000;
	sram_mem[129844] = 16'b0000000000000000;
	sram_mem[129845] = 16'b0000000000000000;
	sram_mem[129846] = 16'b0000000000000000;
	sram_mem[129847] = 16'b0000000000000000;
	sram_mem[129848] = 16'b0000000000000000;
	sram_mem[129849] = 16'b0000000000000000;
	sram_mem[129850] = 16'b0000000000000000;
	sram_mem[129851] = 16'b0000000000000000;
	sram_mem[129852] = 16'b0000000000000000;
	sram_mem[129853] = 16'b0000000000000000;
	sram_mem[129854] = 16'b0000000000000000;
	sram_mem[129855] = 16'b0000000000000000;
	sram_mem[129856] = 16'b0000000000000000;
	sram_mem[129857] = 16'b0000000000000000;
	sram_mem[129858] = 16'b0000000000000000;
	sram_mem[129859] = 16'b0000000000000000;
	sram_mem[129860] = 16'b0000000000000000;
	sram_mem[129861] = 16'b0000000000000000;
	sram_mem[129862] = 16'b0000000000000000;
	sram_mem[129863] = 16'b0000000000000000;
	sram_mem[129864] = 16'b0000000000000000;
	sram_mem[129865] = 16'b0000000000000000;
	sram_mem[129866] = 16'b0000000000000000;
	sram_mem[129867] = 16'b0000000000000000;
	sram_mem[129868] = 16'b0000000000000000;
	sram_mem[129869] = 16'b0000000000000000;
	sram_mem[129870] = 16'b0000000000000000;
	sram_mem[129871] = 16'b0000000000000000;
	sram_mem[129872] = 16'b0000000000000000;
	sram_mem[129873] = 16'b0000000000000000;
	sram_mem[129874] = 16'b0000000000000000;
	sram_mem[129875] = 16'b0000000000000000;
	sram_mem[129876] = 16'b0000000000000000;
	sram_mem[129877] = 16'b0000000000000000;
	sram_mem[129878] = 16'b0000000000000000;
	sram_mem[129879] = 16'b0000000000000000;
	sram_mem[129880] = 16'b0000000000000000;
	sram_mem[129881] = 16'b0000000000000000;
	sram_mem[129882] = 16'b0000000000000000;
	sram_mem[129883] = 16'b0000000000000000;
	sram_mem[129884] = 16'b0000000000000000;
	sram_mem[129885] = 16'b0000000000000000;
	sram_mem[129886] = 16'b0000000000000000;
	sram_mem[129887] = 16'b0000000000000000;
	sram_mem[129888] = 16'b0000000000000000;
	sram_mem[129889] = 16'b0000000000000000;
	sram_mem[129890] = 16'b0000000000000000;
	sram_mem[129891] = 16'b0000000000000000;
	sram_mem[129892] = 16'b0000000000000000;
	sram_mem[129893] = 16'b0000000000000000;
	sram_mem[129894] = 16'b0000000000000000;
	sram_mem[129895] = 16'b0000000000000000;
	sram_mem[129896] = 16'b0000000000000000;
	sram_mem[129897] = 16'b0000000000000000;
	sram_mem[129898] = 16'b0000000000000000;
	sram_mem[129899] = 16'b0000000000000000;
	sram_mem[129900] = 16'b0000000000000000;
	sram_mem[129901] = 16'b0000000000000000;
	sram_mem[129902] = 16'b0000000000000000;
	sram_mem[129903] = 16'b0000000000000000;
	sram_mem[129904] = 16'b0000000000000000;
	sram_mem[129905] = 16'b0000000000000000;
	sram_mem[129906] = 16'b0000000000000000;
	sram_mem[129907] = 16'b0000000000000000;
	sram_mem[129908] = 16'b0000000000000000;
	sram_mem[129909] = 16'b0000000000000000;
	sram_mem[129910] = 16'b0000000000000000;
	sram_mem[129911] = 16'b0000000000000000;
	sram_mem[129912] = 16'b0000000000000000;
	sram_mem[129913] = 16'b0000000000000000;
	sram_mem[129914] = 16'b0000000000000000;
	sram_mem[129915] = 16'b0000000000000000;
	sram_mem[129916] = 16'b0000000000000000;
	sram_mem[129917] = 16'b0000000000000000;
	sram_mem[129918] = 16'b0000000000000000;
	sram_mem[129919] = 16'b0000000000000000;
	sram_mem[129920] = 16'b0000000000000000;
	sram_mem[129921] = 16'b0000000000000000;
	sram_mem[129922] = 16'b0000000000000000;
	sram_mem[129923] = 16'b0000000000000000;
	sram_mem[129924] = 16'b0000000000000000;
	sram_mem[129925] = 16'b0000000000000000;
	sram_mem[129926] = 16'b0000000000000000;
	sram_mem[129927] = 16'b0000000000000000;
	sram_mem[129928] = 16'b0000000000000000;
	sram_mem[129929] = 16'b0000000000000000;
	sram_mem[129930] = 16'b0000000000000000;
	sram_mem[129931] = 16'b0000000000000000;
	sram_mem[129932] = 16'b0000000000000000;
	sram_mem[129933] = 16'b0000000000000000;
	sram_mem[129934] = 16'b0000000000000000;
	sram_mem[129935] = 16'b0000000000000000;
	sram_mem[129936] = 16'b0000000000000000;
	sram_mem[129937] = 16'b0000000000000000;
	sram_mem[129938] = 16'b0000000000000000;
	sram_mem[129939] = 16'b0000000000000000;
	sram_mem[129940] = 16'b0000000000000000;
	sram_mem[129941] = 16'b0000000000000000;
	sram_mem[129942] = 16'b0000000000000000;
	sram_mem[129943] = 16'b0000000000000000;
	sram_mem[129944] = 16'b0000000000000000;
	sram_mem[129945] = 16'b0000000000000000;
	sram_mem[129946] = 16'b0000000000000000;
	sram_mem[129947] = 16'b0000000000000000;
	sram_mem[129948] = 16'b0000000000000000;
	sram_mem[129949] = 16'b0000000000000000;
	sram_mem[129950] = 16'b0000000000000000;
	sram_mem[129951] = 16'b0000000000000000;
	sram_mem[129952] = 16'b0000000000000000;
	sram_mem[129953] = 16'b0000000000000000;
	sram_mem[129954] = 16'b0000000000000000;
	sram_mem[129955] = 16'b0000000000000000;
	sram_mem[129956] = 16'b0000000000000000;
	sram_mem[129957] = 16'b0000000000000000;
	sram_mem[129958] = 16'b0000000000000000;
	sram_mem[129959] = 16'b0000000000000000;
	sram_mem[129960] = 16'b0000000000000000;
	sram_mem[129961] = 16'b0000000000000000;
	sram_mem[129962] = 16'b0000000000000000;
	sram_mem[129963] = 16'b0000000000000000;
	sram_mem[129964] = 16'b0000000000000000;
	sram_mem[129965] = 16'b0000000000000000;
	sram_mem[129966] = 16'b0000000000000000;
	sram_mem[129967] = 16'b0000000000000000;
	sram_mem[129968] = 16'b0000000000000000;
	sram_mem[129969] = 16'b0000000000000000;
	sram_mem[129970] = 16'b0000000000000000;
	sram_mem[129971] = 16'b0000000000000000;
	sram_mem[129972] = 16'b0000000000000000;
	sram_mem[129973] = 16'b0000000000000000;
	sram_mem[129974] = 16'b0000000000000000;
	sram_mem[129975] = 16'b0000000000000000;
	sram_mem[129976] = 16'b0000000000000000;
	sram_mem[129977] = 16'b0000000000000000;
	sram_mem[129978] = 16'b0000000000000000;
	sram_mem[129979] = 16'b0000000000000000;
	sram_mem[129980] = 16'b0000000000000000;
	sram_mem[129981] = 16'b0000000000000000;
	sram_mem[129982] = 16'b0000000000000000;
	sram_mem[129983] = 16'b0000000000000000;
	sram_mem[129984] = 16'b0000000000000000;
	sram_mem[129985] = 16'b0000000000000000;
	sram_mem[129986] = 16'b0000000000000000;
	sram_mem[129987] = 16'b0000000000000000;
	sram_mem[129988] = 16'b0000000000000000;
	sram_mem[129989] = 16'b0000000000000000;
	sram_mem[129990] = 16'b0000000000000000;
	sram_mem[129991] = 16'b0000000000000000;
	sram_mem[129992] = 16'b0000000000000000;
	sram_mem[129993] = 16'b0000000000000000;
	sram_mem[129994] = 16'b0000000000000000;
	sram_mem[129995] = 16'b0000000000000000;
	sram_mem[129996] = 16'b0000000000000000;
	sram_mem[129997] = 16'b0000000000000000;
	sram_mem[129998] = 16'b0000000000000000;
	sram_mem[129999] = 16'b0000000000000000;
	sram_mem[130000] = 16'b0000000000000000;
	sram_mem[130001] = 16'b0000000000000000;
	sram_mem[130002] = 16'b0000000000000000;
	sram_mem[130003] = 16'b0000000000000000;
	sram_mem[130004] = 16'b0000000000000000;
	sram_mem[130005] = 16'b0000000000000000;
	sram_mem[130006] = 16'b0000000000000000;
	sram_mem[130007] = 16'b0000000000000000;
	sram_mem[130008] = 16'b0000000000000000;
	sram_mem[130009] = 16'b0000000000000000;
	sram_mem[130010] = 16'b0000000000000000;
	sram_mem[130011] = 16'b0000000000000000;
	sram_mem[130012] = 16'b0000000000000000;
	sram_mem[130013] = 16'b0000000000000000;
	sram_mem[130014] = 16'b0000000000000000;
	sram_mem[130015] = 16'b0000000000000000;
	sram_mem[130016] = 16'b0000000000000000;
	sram_mem[130017] = 16'b0000000000000000;
	sram_mem[130018] = 16'b0000000000000000;
	sram_mem[130019] = 16'b0000000000000000;
	sram_mem[130020] = 16'b0000000000000000;
	sram_mem[130021] = 16'b0000000000000000;
	sram_mem[130022] = 16'b0000000000000000;
	sram_mem[130023] = 16'b0000000000000000;
	sram_mem[130024] = 16'b0000000000000000;
	sram_mem[130025] = 16'b0000000000000000;
	sram_mem[130026] = 16'b0000000000000000;
	sram_mem[130027] = 16'b0000000000000000;
	sram_mem[130028] = 16'b0000000000000000;
	sram_mem[130029] = 16'b0000000000000000;
	sram_mem[130030] = 16'b0000000000000000;
	sram_mem[130031] = 16'b0000000000000000;
	sram_mem[130032] = 16'b0000000000000000;
	sram_mem[130033] = 16'b0000000000000000;
	sram_mem[130034] = 16'b0000000000000000;
	sram_mem[130035] = 16'b0000000000000000;
	sram_mem[130036] = 16'b0000000000000000;
	sram_mem[130037] = 16'b0000000000000000;
	sram_mem[130038] = 16'b0000000000000000;
	sram_mem[130039] = 16'b0000000000000000;
	sram_mem[130040] = 16'b0000000000000000;
	sram_mem[130041] = 16'b0000000000000000;
	sram_mem[130042] = 16'b0000000000000000;
	sram_mem[130043] = 16'b0000000000000000;
	sram_mem[130044] = 16'b0000000000000000;
	sram_mem[130045] = 16'b0000000000000000;
	sram_mem[130046] = 16'b0000000000000000;
	sram_mem[130047] = 16'b0000000000000000;
	sram_mem[130048] = 16'b0000000000000000;
	sram_mem[130049] = 16'b0000000000000000;
	sram_mem[130050] = 16'b0000000000000000;
	sram_mem[130051] = 16'b0000000000000000;
	sram_mem[130052] = 16'b0000000000000000;
	sram_mem[130053] = 16'b0000000000000000;
	sram_mem[130054] = 16'b0000000000000000;
	sram_mem[130055] = 16'b0000000000000000;
	sram_mem[130056] = 16'b0000000000000000;
	sram_mem[130057] = 16'b0000000000000000;
	sram_mem[130058] = 16'b0000000000000000;
	sram_mem[130059] = 16'b0000000000000000;
	sram_mem[130060] = 16'b0000000000000000;
	sram_mem[130061] = 16'b0000000000000000;
	sram_mem[130062] = 16'b0000000000000000;
	sram_mem[130063] = 16'b0000000000000000;
	sram_mem[130064] = 16'b0000000000000000;
	sram_mem[130065] = 16'b0000000000000000;
	sram_mem[130066] = 16'b0000000000000000;
	sram_mem[130067] = 16'b0000000000000000;
	sram_mem[130068] = 16'b0000000000000000;
	sram_mem[130069] = 16'b0000000000000000;
	sram_mem[130070] = 16'b0000000000000000;
	sram_mem[130071] = 16'b0000000000000000;
	sram_mem[130072] = 16'b0000000000000000;
	sram_mem[130073] = 16'b0000000000000000;
	sram_mem[130074] = 16'b0000000000000000;
	sram_mem[130075] = 16'b0000000000000000;
	sram_mem[130076] = 16'b0000000000000000;
	sram_mem[130077] = 16'b0000000000000000;
	sram_mem[130078] = 16'b0000000000000000;
	sram_mem[130079] = 16'b0000000000000000;
	sram_mem[130080] = 16'b0000000000000000;
	sram_mem[130081] = 16'b0000000000000000;
	sram_mem[130082] = 16'b0000000000000000;
	sram_mem[130083] = 16'b0000000000000000;
	sram_mem[130084] = 16'b0000000000000000;
	sram_mem[130085] = 16'b0000000000000000;
	sram_mem[130086] = 16'b0000000000000000;
	sram_mem[130087] = 16'b0000000000000000;
	sram_mem[130088] = 16'b0000000000000000;
	sram_mem[130089] = 16'b0000000000000000;
	sram_mem[130090] = 16'b0000000000000000;
	sram_mem[130091] = 16'b0000000000000000;
	sram_mem[130092] = 16'b0000000000000000;
	sram_mem[130093] = 16'b0000000000000000;
	sram_mem[130094] = 16'b0000000000000000;
	sram_mem[130095] = 16'b0000000000000000;
	sram_mem[130096] = 16'b0000000000000000;
	sram_mem[130097] = 16'b0000000000000000;
	sram_mem[130098] = 16'b0000000000000000;
	sram_mem[130099] = 16'b0000000000000000;
	sram_mem[130100] = 16'b0000000000000000;
	sram_mem[130101] = 16'b0000000000000000;
	sram_mem[130102] = 16'b0000000000000000;
	sram_mem[130103] = 16'b0000000000000000;
	sram_mem[130104] = 16'b0000000000000000;
	sram_mem[130105] = 16'b0000000000000000;
	sram_mem[130106] = 16'b0000000000000000;
	sram_mem[130107] = 16'b0000000000000000;
	sram_mem[130108] = 16'b0000000000000000;
	sram_mem[130109] = 16'b0000000000000000;
	sram_mem[130110] = 16'b0000000000000000;
	sram_mem[130111] = 16'b0000000000000000;
	sram_mem[130112] = 16'b0000000000000000;
	sram_mem[130113] = 16'b0000000000000000;
	sram_mem[130114] = 16'b0000000000000000;
	sram_mem[130115] = 16'b0000000000000000;
	sram_mem[130116] = 16'b0000000000000000;
	sram_mem[130117] = 16'b0000000000000000;
	sram_mem[130118] = 16'b0000000000000000;
	sram_mem[130119] = 16'b0000000000000000;
	sram_mem[130120] = 16'b0000000000000000;
	sram_mem[130121] = 16'b0000000000000000;
	sram_mem[130122] = 16'b0000000000000000;
	sram_mem[130123] = 16'b0000000000000000;
	sram_mem[130124] = 16'b0000000000000000;
	sram_mem[130125] = 16'b0000000000000000;
	sram_mem[130126] = 16'b0000000000000000;
	sram_mem[130127] = 16'b0000000000000000;
	sram_mem[130128] = 16'b0000000000000000;
	sram_mem[130129] = 16'b0000000000000000;
	sram_mem[130130] = 16'b0000000000000000;
	sram_mem[130131] = 16'b0000000000000000;
	sram_mem[130132] = 16'b0000000000000000;
	sram_mem[130133] = 16'b0000000000000000;
	sram_mem[130134] = 16'b0000000000000000;
	sram_mem[130135] = 16'b0000000000000000;
	sram_mem[130136] = 16'b0000000000000000;
	sram_mem[130137] = 16'b0000000000000000;
	sram_mem[130138] = 16'b0000000000000000;
	sram_mem[130139] = 16'b0000000000000000;
	sram_mem[130140] = 16'b0000000000000000;
	sram_mem[130141] = 16'b0000000000000000;
	sram_mem[130142] = 16'b0000000000000000;
	sram_mem[130143] = 16'b0000000000000000;
	sram_mem[130144] = 16'b0000000000000000;
	sram_mem[130145] = 16'b0000000000000000;
	sram_mem[130146] = 16'b0000000000000000;
	sram_mem[130147] = 16'b0000000000000000;
	sram_mem[130148] = 16'b0000000000000000;
	sram_mem[130149] = 16'b0000000000000000;
	sram_mem[130150] = 16'b0000000000000000;
	sram_mem[130151] = 16'b0000000000000000;
	sram_mem[130152] = 16'b0000000000000000;
	sram_mem[130153] = 16'b0000000000000000;
	sram_mem[130154] = 16'b0000000000000000;
	sram_mem[130155] = 16'b0000000000000000;
	sram_mem[130156] = 16'b0000000000000000;
	sram_mem[130157] = 16'b0000000000000000;
	sram_mem[130158] = 16'b0000000000000000;
	sram_mem[130159] = 16'b0000000000000000;
	sram_mem[130160] = 16'b0000000000000000;
	sram_mem[130161] = 16'b0000000000000000;
	sram_mem[130162] = 16'b0000000000000000;
	sram_mem[130163] = 16'b0000000000000000;
	sram_mem[130164] = 16'b0000000000000000;
	sram_mem[130165] = 16'b0000000000000000;
	sram_mem[130166] = 16'b0000000000000000;
	sram_mem[130167] = 16'b0000000000000000;
	sram_mem[130168] = 16'b0000000000000000;
	sram_mem[130169] = 16'b0000000000000000;
	sram_mem[130170] = 16'b0000000000000000;
	sram_mem[130171] = 16'b0000000000000000;
	sram_mem[130172] = 16'b0000000000000000;
	sram_mem[130173] = 16'b0000000000000000;
	sram_mem[130174] = 16'b0000000000000000;
	sram_mem[130175] = 16'b0000000000000000;
	sram_mem[130176] = 16'b0000000000000000;
	sram_mem[130177] = 16'b0000000000000000;
	sram_mem[130178] = 16'b0000000000000000;
	sram_mem[130179] = 16'b0000000000000000;
	sram_mem[130180] = 16'b0000000000000000;
	sram_mem[130181] = 16'b0000000000000000;
	sram_mem[130182] = 16'b0000000000000000;
	sram_mem[130183] = 16'b0000000000000000;
	sram_mem[130184] = 16'b0000000000000000;
	sram_mem[130185] = 16'b0000000000000000;
	sram_mem[130186] = 16'b0000000000000000;
	sram_mem[130187] = 16'b0000000000000000;
	sram_mem[130188] = 16'b0000000000000000;
	sram_mem[130189] = 16'b0000000000000000;
	sram_mem[130190] = 16'b0000000000000000;
	sram_mem[130191] = 16'b0000000000000000;
	sram_mem[130192] = 16'b0000000000000000;
	sram_mem[130193] = 16'b0000000000000000;
	sram_mem[130194] = 16'b0000000000000000;
	sram_mem[130195] = 16'b0000000000000000;
	sram_mem[130196] = 16'b0000000000000000;
	sram_mem[130197] = 16'b0000000000000000;
	sram_mem[130198] = 16'b0000000000000000;
	sram_mem[130199] = 16'b0000000000000000;
	sram_mem[130200] = 16'b0000000000000000;
	sram_mem[130201] = 16'b0000000000000000;
	sram_mem[130202] = 16'b0000000000000000;
	sram_mem[130203] = 16'b0000000000000000;
	sram_mem[130204] = 16'b0000000000000000;
	sram_mem[130205] = 16'b0000000000000000;
	sram_mem[130206] = 16'b0000000000000000;
	sram_mem[130207] = 16'b0000000000000000;
	sram_mem[130208] = 16'b0000000000000000;
	sram_mem[130209] = 16'b0000000000000000;
	sram_mem[130210] = 16'b0000000000000000;
	sram_mem[130211] = 16'b0000000000000000;
	sram_mem[130212] = 16'b0000000000000000;
	sram_mem[130213] = 16'b0000000000000000;
	sram_mem[130214] = 16'b0000000000000000;
	sram_mem[130215] = 16'b0000000000000000;
	sram_mem[130216] = 16'b0000000000000000;
	sram_mem[130217] = 16'b0000000000000000;
	sram_mem[130218] = 16'b0000000000000000;
	sram_mem[130219] = 16'b0000000000000000;
	sram_mem[130220] = 16'b0000000000000000;
	sram_mem[130221] = 16'b0000000000000000;
	sram_mem[130222] = 16'b0000000000000000;
	sram_mem[130223] = 16'b0000000000000000;
	sram_mem[130224] = 16'b0000000000000000;
	sram_mem[130225] = 16'b0000000000000000;
	sram_mem[130226] = 16'b0000000000000000;
	sram_mem[130227] = 16'b0000000000000000;
	sram_mem[130228] = 16'b0000000000000000;
	sram_mem[130229] = 16'b0000000000000000;
	sram_mem[130230] = 16'b0000000000000000;
	sram_mem[130231] = 16'b0000000000000000;
	sram_mem[130232] = 16'b0000000000000000;
	sram_mem[130233] = 16'b0000000000000000;
	sram_mem[130234] = 16'b0000000000000000;
	sram_mem[130235] = 16'b0000000000000000;
	sram_mem[130236] = 16'b0000000000000000;
	sram_mem[130237] = 16'b0000000000000000;
	sram_mem[130238] = 16'b0000000000000000;
	sram_mem[130239] = 16'b0000000000000000;
	sram_mem[130240] = 16'b0000000000000000;
	sram_mem[130241] = 16'b0000000000000000;
	sram_mem[130242] = 16'b0000000000000000;
	sram_mem[130243] = 16'b0000000000000000;
	sram_mem[130244] = 16'b0000000000000000;
	sram_mem[130245] = 16'b0000000000000000;
	sram_mem[130246] = 16'b0000000000000000;
	sram_mem[130247] = 16'b0000000000000000;
	sram_mem[130248] = 16'b0000000000000000;
	sram_mem[130249] = 16'b0000000000000000;
	sram_mem[130250] = 16'b0000000000000000;
	sram_mem[130251] = 16'b0000000000000000;
	sram_mem[130252] = 16'b0000000000000000;
	sram_mem[130253] = 16'b0000000000000000;
	sram_mem[130254] = 16'b0000000000000000;
	sram_mem[130255] = 16'b0000000000000000;
	sram_mem[130256] = 16'b0000000000000000;
	sram_mem[130257] = 16'b0000000000000000;
	sram_mem[130258] = 16'b0000000000000000;
	sram_mem[130259] = 16'b0000000000000000;
	sram_mem[130260] = 16'b0000000000000000;
	sram_mem[130261] = 16'b0000000000000000;
	sram_mem[130262] = 16'b0000000000000000;
	sram_mem[130263] = 16'b0000000000000000;
	sram_mem[130264] = 16'b0000000000000000;
	sram_mem[130265] = 16'b0000000000000000;
	sram_mem[130266] = 16'b0000000000000000;
	sram_mem[130267] = 16'b0000000000000000;
	sram_mem[130268] = 16'b0000000000000000;
	sram_mem[130269] = 16'b0000000000000000;
	sram_mem[130270] = 16'b0000000000000000;
	sram_mem[130271] = 16'b0000000000000000;
	sram_mem[130272] = 16'b0000000000000000;
	sram_mem[130273] = 16'b0000000000000000;
	sram_mem[130274] = 16'b0000000000000000;
	sram_mem[130275] = 16'b0000000000000000;
	sram_mem[130276] = 16'b0000000000000000;
	sram_mem[130277] = 16'b0000000000000000;
	sram_mem[130278] = 16'b0000000000000000;
	sram_mem[130279] = 16'b0000000000000000;
	sram_mem[130280] = 16'b0000000000000000;
	sram_mem[130281] = 16'b0000000000000000;
	sram_mem[130282] = 16'b0000000000000000;
	sram_mem[130283] = 16'b0000000000000000;
	sram_mem[130284] = 16'b0000000000000000;
	sram_mem[130285] = 16'b0000000000000000;
	sram_mem[130286] = 16'b0000000000000000;
	sram_mem[130287] = 16'b0000000000000000;
	sram_mem[130288] = 16'b0000000000000000;
	sram_mem[130289] = 16'b0000000000000000;
	sram_mem[130290] = 16'b0000000000000000;
	sram_mem[130291] = 16'b0000000000000000;
	sram_mem[130292] = 16'b0000000000000000;
	sram_mem[130293] = 16'b0000000000000000;
	sram_mem[130294] = 16'b0000000000000000;
	sram_mem[130295] = 16'b0000000000000000;
	sram_mem[130296] = 16'b0000000000000000;
	sram_mem[130297] = 16'b0000000000000000;
	sram_mem[130298] = 16'b0000000000000000;
	sram_mem[130299] = 16'b0000000000000000;
	sram_mem[130300] = 16'b0000000000000000;
	sram_mem[130301] = 16'b0000000000000000;
	sram_mem[130302] = 16'b0000000000000000;
	sram_mem[130303] = 16'b0000000000000000;
	sram_mem[130304] = 16'b0000000000000000;
	sram_mem[130305] = 16'b0000000000000000;
	sram_mem[130306] = 16'b0000000000000000;
	sram_mem[130307] = 16'b0000000000000000;
	sram_mem[130308] = 16'b0000000000000000;
	sram_mem[130309] = 16'b0000000000000000;
	sram_mem[130310] = 16'b0000000000000000;
	sram_mem[130311] = 16'b0000000000000000;
	sram_mem[130312] = 16'b0000000000000000;
	sram_mem[130313] = 16'b0000000000000000;
	sram_mem[130314] = 16'b0000000000000000;
	sram_mem[130315] = 16'b0000000000000000;
	sram_mem[130316] = 16'b0000000000000000;
	sram_mem[130317] = 16'b0000000000000000;
	sram_mem[130318] = 16'b0000000000000000;
	sram_mem[130319] = 16'b0000000000000000;
	sram_mem[130320] = 16'b0000000000000000;
	sram_mem[130321] = 16'b0000000000000000;
	sram_mem[130322] = 16'b0000000000000000;
	sram_mem[130323] = 16'b0000000000000000;
	sram_mem[130324] = 16'b0000000000000000;
	sram_mem[130325] = 16'b0000000000000000;
	sram_mem[130326] = 16'b0000000000000000;
	sram_mem[130327] = 16'b0000000000000000;
	sram_mem[130328] = 16'b0000000000000000;
	sram_mem[130329] = 16'b0000000000000000;
	sram_mem[130330] = 16'b0000000000000000;
	sram_mem[130331] = 16'b0000000000000000;
	sram_mem[130332] = 16'b0000000000000000;
	sram_mem[130333] = 16'b0000000000000000;
	sram_mem[130334] = 16'b0000000000000000;
	sram_mem[130335] = 16'b0000000000000000;
	sram_mem[130336] = 16'b0000000000000000;
	sram_mem[130337] = 16'b0000000000000000;
	sram_mem[130338] = 16'b0000000000000000;
	sram_mem[130339] = 16'b0000000000000000;
	sram_mem[130340] = 16'b0000000000000000;
	sram_mem[130341] = 16'b0000000000000000;
	sram_mem[130342] = 16'b0000000000000000;
	sram_mem[130343] = 16'b0000000000000000;
	sram_mem[130344] = 16'b0000000000000000;
	sram_mem[130345] = 16'b0000000000000000;
	sram_mem[130346] = 16'b0000000000000000;
	sram_mem[130347] = 16'b0000000000000000;
	sram_mem[130348] = 16'b0000000000000000;
	sram_mem[130349] = 16'b0000000000000000;
	sram_mem[130350] = 16'b0000000000000000;
	sram_mem[130351] = 16'b0000000000000000;
	sram_mem[130352] = 16'b0000000000000000;
	sram_mem[130353] = 16'b0000000000000000;
	sram_mem[130354] = 16'b0000000000000000;
	sram_mem[130355] = 16'b0000000000000000;
	sram_mem[130356] = 16'b0000000000000000;
	sram_mem[130357] = 16'b0000000000000000;
	sram_mem[130358] = 16'b0000000000000000;
	sram_mem[130359] = 16'b0000000000000000;
	sram_mem[130360] = 16'b0000000000000000;
	sram_mem[130361] = 16'b0000000000000000;
	sram_mem[130362] = 16'b0000000000000000;
	sram_mem[130363] = 16'b0000000000000000;
	sram_mem[130364] = 16'b0000000000000000;
	sram_mem[130365] = 16'b0000000000000000;
	sram_mem[130366] = 16'b0000000000000000;
	sram_mem[130367] = 16'b0000000000000000;
	sram_mem[130368] = 16'b0000000000000000;
	sram_mem[130369] = 16'b0000000000000000;
	sram_mem[130370] = 16'b0000000000000000;
	sram_mem[130371] = 16'b0000000000000000;
	sram_mem[130372] = 16'b0000000000000000;
	sram_mem[130373] = 16'b0000000000000000;
	sram_mem[130374] = 16'b0000000000000000;
	sram_mem[130375] = 16'b0000000000000000;
	sram_mem[130376] = 16'b0000000000000000;
	sram_mem[130377] = 16'b0000000000000000;
	sram_mem[130378] = 16'b0000000000000000;
	sram_mem[130379] = 16'b0000000000000000;
	sram_mem[130380] = 16'b0000000000000000;
	sram_mem[130381] = 16'b0000000000000000;
	sram_mem[130382] = 16'b0000000000000000;
	sram_mem[130383] = 16'b0000000000000000;
	sram_mem[130384] = 16'b0000000000000000;
	sram_mem[130385] = 16'b0000000000000000;
	sram_mem[130386] = 16'b0000000000000000;
	sram_mem[130387] = 16'b0000000000000000;
	sram_mem[130388] = 16'b0000000000000000;
	sram_mem[130389] = 16'b0000000000000000;
	sram_mem[130390] = 16'b0000000000000000;
	sram_mem[130391] = 16'b0000000000000000;
	sram_mem[130392] = 16'b0000000000000000;
	sram_mem[130393] = 16'b0000000000000000;
	sram_mem[130394] = 16'b0000000000000000;
	sram_mem[130395] = 16'b0000000000000000;
	sram_mem[130396] = 16'b0000000000000000;
	sram_mem[130397] = 16'b0000000000000000;
	sram_mem[130398] = 16'b0000000000000000;
	sram_mem[130399] = 16'b0000000000000000;
	sram_mem[130400] = 16'b0000000000000000;
	sram_mem[130401] = 16'b0000000000000000;
	sram_mem[130402] = 16'b0000000000000000;
	sram_mem[130403] = 16'b0000000000000000;
	sram_mem[130404] = 16'b0000000000000000;
	sram_mem[130405] = 16'b0000000000000000;
	sram_mem[130406] = 16'b0000000000000000;
	sram_mem[130407] = 16'b0000000000000000;
	sram_mem[130408] = 16'b0000000000000000;
	sram_mem[130409] = 16'b0000000000000000;
	sram_mem[130410] = 16'b0000000000000000;
	sram_mem[130411] = 16'b0000000000000000;
	sram_mem[130412] = 16'b0000000000000000;
	sram_mem[130413] = 16'b0000000000000000;
	sram_mem[130414] = 16'b0000000000000000;
	sram_mem[130415] = 16'b0000000000000000;
	sram_mem[130416] = 16'b0000000000000000;
	sram_mem[130417] = 16'b0000000000000000;
	sram_mem[130418] = 16'b0000000000000000;
	sram_mem[130419] = 16'b0000000000000000;
	sram_mem[130420] = 16'b0000000000000000;
	sram_mem[130421] = 16'b0000000000000000;
	sram_mem[130422] = 16'b0000000000000000;
	sram_mem[130423] = 16'b0000000000000000;
	sram_mem[130424] = 16'b0000000000000000;
	sram_mem[130425] = 16'b0000000000000000;
	sram_mem[130426] = 16'b0000000000000000;
	sram_mem[130427] = 16'b0000000000000000;
	sram_mem[130428] = 16'b0000000000000000;
	sram_mem[130429] = 16'b0000000000000000;
	sram_mem[130430] = 16'b0000000000000000;
	sram_mem[130431] = 16'b0000000000000000;
	sram_mem[130432] = 16'b0000000000000000;
	sram_mem[130433] = 16'b0000000000000000;
	sram_mem[130434] = 16'b0000000000000000;
	sram_mem[130435] = 16'b0000000000000000;
	sram_mem[130436] = 16'b0000000000000000;
	sram_mem[130437] = 16'b0000000000000000;
	sram_mem[130438] = 16'b0000000000000000;
	sram_mem[130439] = 16'b0000000000000000;
	sram_mem[130440] = 16'b0000000000000000;
	sram_mem[130441] = 16'b0000000000000000;
	sram_mem[130442] = 16'b0000000000000000;
	sram_mem[130443] = 16'b0000000000000000;
	sram_mem[130444] = 16'b0000000000000000;
	sram_mem[130445] = 16'b0000000000000000;
	sram_mem[130446] = 16'b0000000000000000;
	sram_mem[130447] = 16'b0000000000000000;
	sram_mem[130448] = 16'b0000000000000000;
	sram_mem[130449] = 16'b0000000000000000;
	sram_mem[130450] = 16'b0000000000000000;
	sram_mem[130451] = 16'b0000000000000000;
	sram_mem[130452] = 16'b0000000000000000;
	sram_mem[130453] = 16'b0000000000000000;
	sram_mem[130454] = 16'b0000000000000000;
	sram_mem[130455] = 16'b0000000000000000;
	sram_mem[130456] = 16'b0000000000000000;
	sram_mem[130457] = 16'b0000000000000000;
	sram_mem[130458] = 16'b0000000000000000;
	sram_mem[130459] = 16'b0000000000000000;
	sram_mem[130460] = 16'b0000000000000000;
	sram_mem[130461] = 16'b0000000000000000;
	sram_mem[130462] = 16'b0000000000000000;
	sram_mem[130463] = 16'b0000000000000000;
	sram_mem[130464] = 16'b0000000000000000;
	sram_mem[130465] = 16'b0000000000000000;
	sram_mem[130466] = 16'b0000000000000000;
	sram_mem[130467] = 16'b0000000000000000;
	sram_mem[130468] = 16'b0000000000000000;
	sram_mem[130469] = 16'b0000000000000000;
	sram_mem[130470] = 16'b0000000000000000;
	sram_mem[130471] = 16'b0000000000000000;
	sram_mem[130472] = 16'b0000000000000000;
	sram_mem[130473] = 16'b0000000000000000;
	sram_mem[130474] = 16'b0000000000000000;
	sram_mem[130475] = 16'b0000000000000000;
	sram_mem[130476] = 16'b0000000000000000;
	sram_mem[130477] = 16'b0000000000000000;
	sram_mem[130478] = 16'b0000000000000000;
	sram_mem[130479] = 16'b0000000000000000;
	sram_mem[130480] = 16'b0000000000000000;
	sram_mem[130481] = 16'b0000000000000000;
	sram_mem[130482] = 16'b0000000000000000;
	sram_mem[130483] = 16'b0000000000000000;
	sram_mem[130484] = 16'b0000000000000000;
	sram_mem[130485] = 16'b0000000000000000;
	sram_mem[130486] = 16'b0000000000000000;
	sram_mem[130487] = 16'b0000000000000000;
	sram_mem[130488] = 16'b0000000000000000;
	sram_mem[130489] = 16'b0000000000000000;
	sram_mem[130490] = 16'b0000000000000000;
	sram_mem[130491] = 16'b0000000000000000;
	sram_mem[130492] = 16'b0000000000000000;
	sram_mem[130493] = 16'b0000000000000000;
	sram_mem[130494] = 16'b0000000000000000;
	sram_mem[130495] = 16'b0000000000000000;
	sram_mem[130496] = 16'b0000000000000000;
	sram_mem[130497] = 16'b0000000000000000;
	sram_mem[130498] = 16'b0000000000000000;
	sram_mem[130499] = 16'b0000000000000000;
	sram_mem[130500] = 16'b0000000000000000;
	sram_mem[130501] = 16'b0000000000000000;
	sram_mem[130502] = 16'b0000000000000000;
	sram_mem[130503] = 16'b0000000000000000;
	sram_mem[130504] = 16'b0000000000000000;
	sram_mem[130505] = 16'b0000000000000000;
	sram_mem[130506] = 16'b0000000000000000;
	sram_mem[130507] = 16'b0000000000000000;
	sram_mem[130508] = 16'b0000000000000000;
	sram_mem[130509] = 16'b0000000000000000;
	sram_mem[130510] = 16'b0000000000000000;
	sram_mem[130511] = 16'b0000000000000000;
	sram_mem[130512] = 16'b0000000000000000;
	sram_mem[130513] = 16'b0000000000000000;
	sram_mem[130514] = 16'b0000000000000000;
	sram_mem[130515] = 16'b0000000000000000;
	sram_mem[130516] = 16'b0000000000000000;
	sram_mem[130517] = 16'b0000000000000000;
	sram_mem[130518] = 16'b0000000000000000;
	sram_mem[130519] = 16'b0000000000000000;
	sram_mem[130520] = 16'b0000000000000000;
	sram_mem[130521] = 16'b0000000000000000;
	sram_mem[130522] = 16'b0000000000000000;
	sram_mem[130523] = 16'b0000000000000000;
	sram_mem[130524] = 16'b0000000000000000;
	sram_mem[130525] = 16'b0000000000000000;
	sram_mem[130526] = 16'b0000000000000000;
	sram_mem[130527] = 16'b0000000000000000;
	sram_mem[130528] = 16'b0000000000000000;
	sram_mem[130529] = 16'b0000000000000000;
	sram_mem[130530] = 16'b0000000000000000;
	sram_mem[130531] = 16'b0000000000000000;
	sram_mem[130532] = 16'b0000000000000000;
	sram_mem[130533] = 16'b0000000000000000;
	sram_mem[130534] = 16'b0000000000000000;
	sram_mem[130535] = 16'b0000000000000000;
	sram_mem[130536] = 16'b0000000000000000;
	sram_mem[130537] = 16'b0000000000000000;
	sram_mem[130538] = 16'b0000000000000000;
	sram_mem[130539] = 16'b0000000000000000;
	sram_mem[130540] = 16'b0000000000000000;
	sram_mem[130541] = 16'b0000000000000000;
	sram_mem[130542] = 16'b0000000000000000;
	sram_mem[130543] = 16'b0000000000000000;
	sram_mem[130544] = 16'b0000000000000000;
	sram_mem[130545] = 16'b0000000000000000;
	sram_mem[130546] = 16'b0000000000000000;
	sram_mem[130547] = 16'b0000000000000000;
	sram_mem[130548] = 16'b0000000000000000;
	sram_mem[130549] = 16'b0000000000000000;
	sram_mem[130550] = 16'b0000000000000000;
	sram_mem[130551] = 16'b0000000000000000;
	sram_mem[130552] = 16'b0000000000000000;
	sram_mem[130553] = 16'b0000000000000000;
	sram_mem[130554] = 16'b0000000000000000;
	sram_mem[130555] = 16'b0000000000000000;
	sram_mem[130556] = 16'b0000000000000000;
	sram_mem[130557] = 16'b0000000000000000;
	sram_mem[130558] = 16'b0000000000000000;
	sram_mem[130559] = 16'b0000000000000000;
	sram_mem[130560] = 16'b0000000000000000;
	sram_mem[130561] = 16'b0000000000000000;
	sram_mem[130562] = 16'b0000000000000000;
	sram_mem[130563] = 16'b0000000000000000;
	sram_mem[130564] = 16'b0000000000000000;
	sram_mem[130565] = 16'b0000000000000000;
	sram_mem[130566] = 16'b0000000000000000;
	sram_mem[130567] = 16'b0000000000000000;
	sram_mem[130568] = 16'b0000000000000000;
	sram_mem[130569] = 16'b0000000000000000;
	sram_mem[130570] = 16'b0000000000000000;
	sram_mem[130571] = 16'b0000000000000000;
	sram_mem[130572] = 16'b0000000000000000;
	sram_mem[130573] = 16'b0000000000000000;
	sram_mem[130574] = 16'b0000000000000000;
	sram_mem[130575] = 16'b0000000000000000;
	sram_mem[130576] = 16'b0000000000000000;
	sram_mem[130577] = 16'b0000000000000000;
	sram_mem[130578] = 16'b0000000000000000;
	sram_mem[130579] = 16'b0000000000000000;
	sram_mem[130580] = 16'b0000000000000000;
	sram_mem[130581] = 16'b0000000000000000;
	sram_mem[130582] = 16'b0000000000000000;
	sram_mem[130583] = 16'b0000000000000000;
	sram_mem[130584] = 16'b0000000000000000;
	sram_mem[130585] = 16'b0000000000000000;
	sram_mem[130586] = 16'b0000000000000000;
	sram_mem[130587] = 16'b0000000000000000;
	sram_mem[130588] = 16'b0000000000000000;
	sram_mem[130589] = 16'b0000000000000000;
	sram_mem[130590] = 16'b0000000000000000;
	sram_mem[130591] = 16'b0000000000000000;
	sram_mem[130592] = 16'b0000000000000000;
	sram_mem[130593] = 16'b0000000000000000;
	sram_mem[130594] = 16'b0000000000000000;
	sram_mem[130595] = 16'b0000000000000000;
	sram_mem[130596] = 16'b0000000000000000;
	sram_mem[130597] = 16'b0000000000000000;
	sram_mem[130598] = 16'b0000000000000000;
	sram_mem[130599] = 16'b0000000000000000;
	sram_mem[130600] = 16'b0000000000000000;
	sram_mem[130601] = 16'b0000000000000000;
	sram_mem[130602] = 16'b0000000000000000;
	sram_mem[130603] = 16'b0000000000000000;
	sram_mem[130604] = 16'b0000000000000000;
	sram_mem[130605] = 16'b0000000000000000;
	sram_mem[130606] = 16'b0000000000000000;
	sram_mem[130607] = 16'b0000000000000000;
	sram_mem[130608] = 16'b0000000000000000;
	sram_mem[130609] = 16'b0000000000000000;
	sram_mem[130610] = 16'b0000000000000000;
	sram_mem[130611] = 16'b0000000000000000;
	sram_mem[130612] = 16'b0000000000000000;
	sram_mem[130613] = 16'b0000000000000000;
	sram_mem[130614] = 16'b0000000000000000;
	sram_mem[130615] = 16'b0000000000000000;
	sram_mem[130616] = 16'b0000000000000000;
	sram_mem[130617] = 16'b0000000000000000;
	sram_mem[130618] = 16'b0000000000000000;
	sram_mem[130619] = 16'b0000000000000000;
	sram_mem[130620] = 16'b0000000000000000;
	sram_mem[130621] = 16'b0000000000000000;
	sram_mem[130622] = 16'b0000000000000000;
	sram_mem[130623] = 16'b0000000000000000;
	sram_mem[130624] = 16'b0000000000000000;
	sram_mem[130625] = 16'b0000000000000000;
	sram_mem[130626] = 16'b0000000000000000;
	sram_mem[130627] = 16'b0000000000000000;
	sram_mem[130628] = 16'b0000000000000000;
	sram_mem[130629] = 16'b0000000000000000;
	sram_mem[130630] = 16'b0000000000000000;
	sram_mem[130631] = 16'b0000000000000000;
	sram_mem[130632] = 16'b0000000000000000;
	sram_mem[130633] = 16'b0000000000000000;
	sram_mem[130634] = 16'b0000000000000000;
	sram_mem[130635] = 16'b0000000000000000;
	sram_mem[130636] = 16'b0000000000000000;
	sram_mem[130637] = 16'b0000000000000000;
	sram_mem[130638] = 16'b0000000000000000;
	sram_mem[130639] = 16'b0000000000000000;
	sram_mem[130640] = 16'b0000000000000000;
	sram_mem[130641] = 16'b0000000000000000;
	sram_mem[130642] = 16'b0000000000000000;
	sram_mem[130643] = 16'b0000000000000000;
	sram_mem[130644] = 16'b0000000000000000;
	sram_mem[130645] = 16'b0000000000000000;
	sram_mem[130646] = 16'b0000000000000000;
	sram_mem[130647] = 16'b0000000000000000;
	sram_mem[130648] = 16'b0000000000000000;
	sram_mem[130649] = 16'b0000000000000000;
	sram_mem[130650] = 16'b0000000000000000;
	sram_mem[130651] = 16'b0000000000000000;
	sram_mem[130652] = 16'b0000000000000000;
	sram_mem[130653] = 16'b0000000000000000;
	sram_mem[130654] = 16'b0000000000000000;
	sram_mem[130655] = 16'b0000000000000000;
	sram_mem[130656] = 16'b0000000000000000;
	sram_mem[130657] = 16'b0000000000000000;
	sram_mem[130658] = 16'b0000000000000000;
	sram_mem[130659] = 16'b0000000000000000;
	sram_mem[130660] = 16'b0000000000000000;
	sram_mem[130661] = 16'b0000000000000000;
	sram_mem[130662] = 16'b0000000000000000;
	sram_mem[130663] = 16'b0000000000000000;
	sram_mem[130664] = 16'b0000000000000000;
	sram_mem[130665] = 16'b0000000000000000;
	sram_mem[130666] = 16'b0000000000000000;
	sram_mem[130667] = 16'b0000000000000000;
	sram_mem[130668] = 16'b0000000000000000;
	sram_mem[130669] = 16'b0000000000000000;
	sram_mem[130670] = 16'b0000000000000000;
	sram_mem[130671] = 16'b0000000000000000;
	sram_mem[130672] = 16'b0000000000000000;
	sram_mem[130673] = 16'b0000000000000000;
	sram_mem[130674] = 16'b0000000000000000;
	sram_mem[130675] = 16'b0000000000000000;
	sram_mem[130676] = 16'b0000000000000000;
	sram_mem[130677] = 16'b0000000000000000;
	sram_mem[130678] = 16'b0000000000000000;
	sram_mem[130679] = 16'b0000000000000000;
	sram_mem[130680] = 16'b0000000000000000;
	sram_mem[130681] = 16'b0000000000000000;
	sram_mem[130682] = 16'b0000000000000000;
	sram_mem[130683] = 16'b0000000000000000;
	sram_mem[130684] = 16'b0000000000000000;
	sram_mem[130685] = 16'b0000000000000000;
	sram_mem[130686] = 16'b0000000000000000;
	sram_mem[130687] = 16'b0000000000000000;
	sram_mem[130688] = 16'b0000000000000000;
	sram_mem[130689] = 16'b0000000000000000;
	sram_mem[130690] = 16'b0000000000000000;
	sram_mem[130691] = 16'b0000000000000000;
	sram_mem[130692] = 16'b0000000000000000;
	sram_mem[130693] = 16'b0000000000000000;
	sram_mem[130694] = 16'b0000000000000000;
	sram_mem[130695] = 16'b0000000000000000;
	sram_mem[130696] = 16'b0000000000000000;
	sram_mem[130697] = 16'b0000000000000000;
	sram_mem[130698] = 16'b0000000000000000;
	sram_mem[130699] = 16'b0000000000000000;
	sram_mem[130700] = 16'b0000000000000000;
	sram_mem[130701] = 16'b0000000000000000;
	sram_mem[130702] = 16'b0000000000000000;
	sram_mem[130703] = 16'b0000000000000000;
	sram_mem[130704] = 16'b0000000000000000;
	sram_mem[130705] = 16'b0000000000000000;
	sram_mem[130706] = 16'b0000000000000000;
	sram_mem[130707] = 16'b0000000000000000;
	sram_mem[130708] = 16'b0000000000000000;
	sram_mem[130709] = 16'b0000000000000000;
	sram_mem[130710] = 16'b0000000000000000;
	sram_mem[130711] = 16'b0000000000000000;
	sram_mem[130712] = 16'b0000000000000000;
	sram_mem[130713] = 16'b0000000000000000;
	sram_mem[130714] = 16'b0000000000000000;
	sram_mem[130715] = 16'b0000000000000000;
	sram_mem[130716] = 16'b0000000000000000;
	sram_mem[130717] = 16'b0000000000000000;
	sram_mem[130718] = 16'b0000000000000000;
	sram_mem[130719] = 16'b0000000000000000;
	sram_mem[130720] = 16'b0000000000000000;
	sram_mem[130721] = 16'b0000000000000000;
	sram_mem[130722] = 16'b0000000000000000;
	sram_mem[130723] = 16'b0000000000000000;
	sram_mem[130724] = 16'b0000000000000000;
	sram_mem[130725] = 16'b0000000000000000;
	sram_mem[130726] = 16'b0000000000000000;
	sram_mem[130727] = 16'b0000000000000000;
	sram_mem[130728] = 16'b0000000000000000;
	sram_mem[130729] = 16'b0000000000000000;
	sram_mem[130730] = 16'b0000000000000000;
	sram_mem[130731] = 16'b0000000000000000;
	sram_mem[130732] = 16'b0000000000000000;
	sram_mem[130733] = 16'b0000000000000000;
	sram_mem[130734] = 16'b0000000000000000;
	sram_mem[130735] = 16'b0000000000000000;
	sram_mem[130736] = 16'b0000000000000000;
	sram_mem[130737] = 16'b0000000000000000;
	sram_mem[130738] = 16'b0000000000000000;
	sram_mem[130739] = 16'b0000000000000000;
	sram_mem[130740] = 16'b0000000000000000;
	sram_mem[130741] = 16'b0000000000000000;
	sram_mem[130742] = 16'b0000000000000000;
	sram_mem[130743] = 16'b0000000000000000;
	sram_mem[130744] = 16'b0000000000000000;
	sram_mem[130745] = 16'b0000000000000000;
	sram_mem[130746] = 16'b0000000000000000;
	sram_mem[130747] = 16'b0000000000000000;
	sram_mem[130748] = 16'b0000000000000000;
	sram_mem[130749] = 16'b0000000000000000;
	sram_mem[130750] = 16'b0000000000000000;
	sram_mem[130751] = 16'b0000000000000000;
	sram_mem[130752] = 16'b0000000000000000;
	sram_mem[130753] = 16'b0000000000000000;
	sram_mem[130754] = 16'b0000000000000000;
	sram_mem[130755] = 16'b0000000000000000;
	sram_mem[130756] = 16'b0000000000000000;
	sram_mem[130757] = 16'b0000000000000000;
	sram_mem[130758] = 16'b0000000000000000;
	sram_mem[130759] = 16'b0000000000000000;
	sram_mem[130760] = 16'b0000000000000000;
	sram_mem[130761] = 16'b0000000000000000;
	sram_mem[130762] = 16'b0000000000000000;
	sram_mem[130763] = 16'b0000000000000000;
	sram_mem[130764] = 16'b0000000000000000;
	sram_mem[130765] = 16'b0000000000000000;
	sram_mem[130766] = 16'b0000000000000000;
	sram_mem[130767] = 16'b0000000000000000;
	sram_mem[130768] = 16'b0000000000000000;
	sram_mem[130769] = 16'b0000000000000000;
	sram_mem[130770] = 16'b0000000000000000;
	sram_mem[130771] = 16'b0000000000000000;
	sram_mem[130772] = 16'b0000000000000000;
	sram_mem[130773] = 16'b0000000000000000;
	sram_mem[130774] = 16'b0000000000000000;
	sram_mem[130775] = 16'b0000000000000000;
	sram_mem[130776] = 16'b0000000000000000;
	sram_mem[130777] = 16'b0000000000000000;
	sram_mem[130778] = 16'b0000000000000000;
	sram_mem[130779] = 16'b0000000000000000;
	sram_mem[130780] = 16'b0000000000000000;
	sram_mem[130781] = 16'b0000000000000000;
	sram_mem[130782] = 16'b0000000000000000;
	sram_mem[130783] = 16'b0000000000000000;
	sram_mem[130784] = 16'b0000000000000000;
	sram_mem[130785] = 16'b0000000000000000;
	sram_mem[130786] = 16'b0000000000000000;
	sram_mem[130787] = 16'b0000000000000000;
	sram_mem[130788] = 16'b0000000000000000;
	sram_mem[130789] = 16'b0000000000000000;
	sram_mem[130790] = 16'b0000000000000000;
	sram_mem[130791] = 16'b0000000000000000;
	sram_mem[130792] = 16'b0000000000000000;
	sram_mem[130793] = 16'b0000000000000000;
	sram_mem[130794] = 16'b0000000000000000;
	sram_mem[130795] = 16'b0000000000000000;
	sram_mem[130796] = 16'b0000000000000000;
	sram_mem[130797] = 16'b0000000000000000;
	sram_mem[130798] = 16'b0000000000000000;
	sram_mem[130799] = 16'b0000000000000000;
	sram_mem[130800] = 16'b0000000000000000;
	sram_mem[130801] = 16'b0000000000000000;
	sram_mem[130802] = 16'b0000000000000000;
	sram_mem[130803] = 16'b0000000000000000;
	sram_mem[130804] = 16'b0000000000000000;
	sram_mem[130805] = 16'b0000000000000000;
	sram_mem[130806] = 16'b0000000000000000;
	sram_mem[130807] = 16'b0000000000000000;
	sram_mem[130808] = 16'b0000000000000000;
	sram_mem[130809] = 16'b0000000000000000;
	sram_mem[130810] = 16'b0000000000000000;
	sram_mem[130811] = 16'b0000000000000000;
	sram_mem[130812] = 16'b0000000000000000;
	sram_mem[130813] = 16'b0000000000000000;
	sram_mem[130814] = 16'b0000000000000000;
	sram_mem[130815] = 16'b0000000000000000;
	sram_mem[130816] = 16'b0000000000000000;
	sram_mem[130817] = 16'b0000000000000000;
	sram_mem[130818] = 16'b0000000000000000;
	sram_mem[130819] = 16'b0000000000000000;
	sram_mem[130820] = 16'b0000000000000000;
	sram_mem[130821] = 16'b0000000000000000;
	sram_mem[130822] = 16'b0000000000000000;
	sram_mem[130823] = 16'b0000000000000000;
	sram_mem[130824] = 16'b0000000000000000;
	sram_mem[130825] = 16'b0000000000000000;
	sram_mem[130826] = 16'b0000000000000000;
	sram_mem[130827] = 16'b0000000000000000;
	sram_mem[130828] = 16'b0000000000000000;
	sram_mem[130829] = 16'b0000000000000000;
	sram_mem[130830] = 16'b0000000000000000;
	sram_mem[130831] = 16'b0000000000000000;
	sram_mem[130832] = 16'b0000000000000000;
	sram_mem[130833] = 16'b0000000000000000;
	sram_mem[130834] = 16'b0000000000000000;
	sram_mem[130835] = 16'b0000000000000000;
	sram_mem[130836] = 16'b0000000000000000;
	sram_mem[130837] = 16'b0000000000000000;
	sram_mem[130838] = 16'b0000000000000000;
	sram_mem[130839] = 16'b0000000000000000;
	sram_mem[130840] = 16'b0000000000000000;
	sram_mem[130841] = 16'b0000000000000000;
	sram_mem[130842] = 16'b0000000000000000;
	sram_mem[130843] = 16'b0000000000000000;
	sram_mem[130844] = 16'b0000000000000000;
	sram_mem[130845] = 16'b0000000000000000;
	sram_mem[130846] = 16'b0000000000000000;
	sram_mem[130847] = 16'b0000000000000000;
	sram_mem[130848] = 16'b0000000000000000;
	sram_mem[130849] = 16'b0000000000000000;
	sram_mem[130850] = 16'b0000000000000000;
	sram_mem[130851] = 16'b0000000000000000;
	sram_mem[130852] = 16'b0000000000000000;
	sram_mem[130853] = 16'b0000000000000000;
	sram_mem[130854] = 16'b0000000000000000;
	sram_mem[130855] = 16'b0000000000000000;
	sram_mem[130856] = 16'b0000000000000000;
	sram_mem[130857] = 16'b0000000000000000;
	sram_mem[130858] = 16'b0000000000000000;
	sram_mem[130859] = 16'b0000000000000000;
	sram_mem[130860] = 16'b0000000000000000;
	sram_mem[130861] = 16'b0000000000000000;
	sram_mem[130862] = 16'b0000000000000000;
	sram_mem[130863] = 16'b0000000000000000;
	sram_mem[130864] = 16'b0000000000000000;
	sram_mem[130865] = 16'b0000000000000000;
	sram_mem[130866] = 16'b0000000000000000;
	sram_mem[130867] = 16'b0000000000000000;
	sram_mem[130868] = 16'b0000000000000000;
	sram_mem[130869] = 16'b0000000000000000;
	sram_mem[130870] = 16'b0000000000000000;
	sram_mem[130871] = 16'b0000000000000000;
	sram_mem[130872] = 16'b0000000000000000;
	sram_mem[130873] = 16'b0000000000000000;
	sram_mem[130874] = 16'b0000000000000000;
	sram_mem[130875] = 16'b0000000000000000;
	sram_mem[130876] = 16'b0000000000000000;
	sram_mem[130877] = 16'b0000000000000000;
	sram_mem[130878] = 16'b0000000000000000;
	sram_mem[130879] = 16'b0000000000000000;
	sram_mem[130880] = 16'b0000000000000000;
	sram_mem[130881] = 16'b0000000000000000;
	sram_mem[130882] = 16'b0000000000000000;
	sram_mem[130883] = 16'b0000000000000000;
	sram_mem[130884] = 16'b0000000000000000;
	sram_mem[130885] = 16'b0000000000000000;
	sram_mem[130886] = 16'b0000000000000000;
	sram_mem[130887] = 16'b0000000000000000;
	sram_mem[130888] = 16'b0000000000000000;
	sram_mem[130889] = 16'b0000000000000000;
	sram_mem[130890] = 16'b0000000000000000;
	sram_mem[130891] = 16'b0000000000000000;
	sram_mem[130892] = 16'b0000000000000000;
	sram_mem[130893] = 16'b0000000000000000;
	sram_mem[130894] = 16'b0000000000000000;
	sram_mem[130895] = 16'b0000000000000000;
	sram_mem[130896] = 16'b0000000000000000;
	sram_mem[130897] = 16'b0000000000000000;
	sram_mem[130898] = 16'b0000000000000000;
	sram_mem[130899] = 16'b0000000000000000;
	sram_mem[130900] = 16'b0000000000000000;
	sram_mem[130901] = 16'b0000000000000000;
	sram_mem[130902] = 16'b0000000000000000;
	sram_mem[130903] = 16'b0000000000000000;
	sram_mem[130904] = 16'b0000000000000000;
	sram_mem[130905] = 16'b0000000000000000;
	sram_mem[130906] = 16'b0000000000000000;
	sram_mem[130907] = 16'b0000000000000000;
	sram_mem[130908] = 16'b0000000000000000;
	sram_mem[130909] = 16'b0000000000000000;
	sram_mem[130910] = 16'b0000000000000000;
	sram_mem[130911] = 16'b0000000000000000;
	sram_mem[130912] = 16'b0000000000000000;
	sram_mem[130913] = 16'b0000000000000000;
	sram_mem[130914] = 16'b0000000000000000;
	sram_mem[130915] = 16'b0000000000000000;
	sram_mem[130916] = 16'b0000000000000000;
	sram_mem[130917] = 16'b0000000000000000;
	sram_mem[130918] = 16'b0000000000000000;
	sram_mem[130919] = 16'b0000000000000000;
	sram_mem[130920] = 16'b0000000000000000;
	sram_mem[130921] = 16'b0000000000000000;
	sram_mem[130922] = 16'b0000000000000000;
	sram_mem[130923] = 16'b0000000000000000;
	sram_mem[130924] = 16'b0000000000000000;
	sram_mem[130925] = 16'b0000000000000000;
	sram_mem[130926] = 16'b0000000000000000;
	sram_mem[130927] = 16'b0000000000000000;
	sram_mem[130928] = 16'b0000000000000000;
	sram_mem[130929] = 16'b0000000000000000;
	sram_mem[130930] = 16'b0000000000000000;
	sram_mem[130931] = 16'b0000000000000000;
	sram_mem[130932] = 16'b0000000000000000;
	sram_mem[130933] = 16'b0000000000000000;
	sram_mem[130934] = 16'b0000000000000000;
	sram_mem[130935] = 16'b0000000000000000;
	sram_mem[130936] = 16'b0000000000000000;
	sram_mem[130937] = 16'b0000000000000000;
	sram_mem[130938] = 16'b0000000000000000;
	sram_mem[130939] = 16'b0000000000000000;
	sram_mem[130940] = 16'b0000000000000000;
	sram_mem[130941] = 16'b0000000000000000;
	sram_mem[130942] = 16'b0000000000000000;
	sram_mem[130943] = 16'b0000000000000000;
	sram_mem[130944] = 16'b0000000000000000;
	sram_mem[130945] = 16'b0000000000000000;
	sram_mem[130946] = 16'b0000000000000000;
	sram_mem[130947] = 16'b0000000000000000;
	sram_mem[130948] = 16'b0000000000000000;
	sram_mem[130949] = 16'b0000000000000000;
	sram_mem[130950] = 16'b0000000000000000;
	sram_mem[130951] = 16'b0000000000000000;
	sram_mem[130952] = 16'b0000000000000000;
	sram_mem[130953] = 16'b0000000000000000;
	sram_mem[130954] = 16'b0000000000000000;
	sram_mem[130955] = 16'b0000000000000000;
	sram_mem[130956] = 16'b0000000000000000;
	sram_mem[130957] = 16'b0000000000000000;
	sram_mem[130958] = 16'b0000000000000000;
	sram_mem[130959] = 16'b0000000000000000;
	sram_mem[130960] = 16'b0000000000000000;
	sram_mem[130961] = 16'b0000000000000000;
	sram_mem[130962] = 16'b0000000000000000;
	sram_mem[130963] = 16'b0000000000000000;
	sram_mem[130964] = 16'b0000000000000000;
	sram_mem[130965] = 16'b0000000000000000;
	sram_mem[130966] = 16'b0000000000000000;
	sram_mem[130967] = 16'b0000000000000000;
	sram_mem[130968] = 16'b0000000000000000;
	sram_mem[130969] = 16'b0000000000000000;
	sram_mem[130970] = 16'b0000000000000000;
	sram_mem[130971] = 16'b0000000000000000;
	sram_mem[130972] = 16'b0000000000000000;
	sram_mem[130973] = 16'b0000000000000000;
	sram_mem[130974] = 16'b0000000000000000;
	sram_mem[130975] = 16'b0000000000000000;
	sram_mem[130976] = 16'b0000000000000000;
	sram_mem[130977] = 16'b0000000000000000;
	sram_mem[130978] = 16'b0000000000000000;
	sram_mem[130979] = 16'b0000000000000000;
	sram_mem[130980] = 16'b0000000000000000;
	sram_mem[130981] = 16'b0000000000000000;
	sram_mem[130982] = 16'b0000000000000000;
	sram_mem[130983] = 16'b0000000000000000;
	sram_mem[130984] = 16'b0000000000000000;
	sram_mem[130985] = 16'b0000000000000000;
	sram_mem[130986] = 16'b0000000000000000;
	sram_mem[130987] = 16'b0000000000000000;
	sram_mem[130988] = 16'b0000000000000000;
	sram_mem[130989] = 16'b0000000000000000;
	sram_mem[130990] = 16'b0000000000000000;
	sram_mem[130991] = 16'b0000000000000000;
	sram_mem[130992] = 16'b0000000000000000;
	sram_mem[130993] = 16'b0000000000000000;
	sram_mem[130994] = 16'b0000000000000000;
	sram_mem[130995] = 16'b0000000000000000;
	sram_mem[130996] = 16'b0000000000000000;
	sram_mem[130997] = 16'b0000000000000000;
	sram_mem[130998] = 16'b0000000000000000;
	sram_mem[130999] = 16'b0000000000000000;
	sram_mem[131000] = 16'b0000000000000000;
	sram_mem[131001] = 16'b0000000000000000;
	sram_mem[131002] = 16'b0000000000000000;
	sram_mem[131003] = 16'b0000000000000000;
	sram_mem[131004] = 16'b0000000000000000;
	sram_mem[131005] = 16'b0000000000000000;
	sram_mem[131006] = 16'b0000000000000000;
	sram_mem[131007] = 16'b0000000000000000;
	sram_mem[131008] = 16'b0000000000000000;
	sram_mem[131009] = 16'b0000000000000000;
	sram_mem[131010] = 16'b0000000000000000;
	sram_mem[131011] = 16'b0000000000000000;
	sram_mem[131012] = 16'b0000000000000000;
	sram_mem[131013] = 16'b0000000000000000;
	sram_mem[131014] = 16'b0000000000000000;
	sram_mem[131015] = 16'b0000000000000000;
	sram_mem[131016] = 16'b0000000000000000;
	sram_mem[131017] = 16'b0000000000000000;
	sram_mem[131018] = 16'b0000000000000000;
	sram_mem[131019] = 16'b0000000000000000;
	sram_mem[131020] = 16'b0000000000000000;
	sram_mem[131021] = 16'b0000000000000000;
	sram_mem[131022] = 16'b0000000000000000;
	sram_mem[131023] = 16'b0000000000000000;
	sram_mem[131024] = 16'b0000000000000000;
	sram_mem[131025] = 16'b0000000000000000;
	sram_mem[131026] = 16'b0000000000000000;
	sram_mem[131027] = 16'b0000000000000000;
	sram_mem[131028] = 16'b0000000000000000;
	sram_mem[131029] = 16'b0000000000000000;
	sram_mem[131030] = 16'b0000000000000000;
	sram_mem[131031] = 16'b0000000000000000;
	sram_mem[131032] = 16'b0000000000000000;
	sram_mem[131033] = 16'b0000000000000000;
	sram_mem[131034] = 16'b0000000000000000;
	sram_mem[131035] = 16'b0000000000000000;
	sram_mem[131036] = 16'b0000000000000000;
	sram_mem[131037] = 16'b0000000000000000;
	sram_mem[131038] = 16'b0000000000000000;
	sram_mem[131039] = 16'b0000000000000000;
	sram_mem[131040] = 16'b0000000000000000;
	sram_mem[131041] = 16'b0000000000000000;
	sram_mem[131042] = 16'b0000000000000000;
	sram_mem[131043] = 16'b0000000000000000;
	sram_mem[131044] = 16'b0000000000000000;
	sram_mem[131045] = 16'b0000000000000000;
	sram_mem[131046] = 16'b0000000000000000;
	sram_mem[131047] = 16'b0000000000000000;
	sram_mem[131048] = 16'b0000000000000000;
	sram_mem[131049] = 16'b0000000000000000;
	sram_mem[131050] = 16'b0000000000000000;
	sram_mem[131051] = 16'b0000000000000000;
	sram_mem[131052] = 16'b0000000000000000;
	sram_mem[131053] = 16'b0000000000000000;
	sram_mem[131054] = 16'b0000000000000000;
	sram_mem[131055] = 16'b0000000000000000;
	sram_mem[131056] = 16'b0000000000000000;
	sram_mem[131057] = 16'b0000000000000000;
	sram_mem[131058] = 16'b0000000000000000;
	sram_mem[131059] = 16'b0000000000000000;
	sram_mem[131060] = 16'b0000000000000000;
	sram_mem[131061] = 16'b0000000000000000;
	sram_mem[131062] = 16'b0000000000000000;
	sram_mem[131063] = 16'b0000000000000000;
	sram_mem[131064] = 16'b0000000000000000;
	sram_mem[131065] = 16'b0000000000000000;
	sram_mem[131066] = 16'b0000000000000000;
	sram_mem[131067] = 16'b0000000000000000;
	sram_mem[131068] = 16'b0000000000000000;
	sram_mem[131069] = 16'b0000000000000000;
	sram_mem[131070] = 16'b0000000000000000;
	sram_mem[131071] = 16'b0000000000000000;
end
endmodule